module alu_fsm_tb();

reg     in_clka,
        in_clkb,
        reset_in,
        n_dec_in,
        z_dec_in,
        p_dec_in,
        n_alu_in,
        z_alu_in,
        p_alu_in,
        we_reg_in,
        br_in;

wire [2:0] state_out;
wire pc_ctl_0_out;

//create an FSM instance.
ALU_FSM fsm (
        .clka (in_clka),
        .clkb (in_clkb),
        .reset_in (reset_in),
        .n_dec_in (n_dec_in),
        .z_dec_in (z_dec_in),
        .p_dec_in (p_dec_in),
        .n_alu_in (n_alu_in),
        .z_alu_in (z_alu_in),
        .p_alu_in (p_alu_in),
        .we_reg_in (we_reg_in),
        .br_in (br_in),
        .pc_ctl_0_out (pc_ctl_0_out),
        .state_out (state_out)
);

initial begin

reset_in = 0;
n_dec_in = 0;
z_dec_in = 0;
p_dec_in = 0;
n_alu_in = 0;
z_alu_in = 0;
p_alu_in = 0;
we_reg_in = 0;
br_in = 0;
in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

reset_in = 1; //reset fsm

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

reset_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

/**
The following blocks test that the state is not updated when the we signal is 
not asserted 
**/ 

n_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

n_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

/**
The following tests verify that the FSM moves between states properly
**/
we_reg_in = 1;
n_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

n_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

/**
The following test check that the ALU Properly asserts the 
branch out bit when it should
**/

n_alu_in = 1; //set state to n

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

n_alu_in = 0;
n_dec_in = 1;
br_in = 1; //should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 1;
n_dec_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_alu_in = 0;
z_dec_in = 1;
br_in = 1; // should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 1;
z_dec_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 0;
p_dec_in = 1;
br_in = 1; //should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


/**
The following tests verify that the branch is asserted soon enough
**/

n_alu_in = 1;
n_dec_in = 1;
p_dec_in = 0;
br_in = 1; //should assert branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 1;
p_dec_in = 1; //should cause branch
n_alu_in = 0;
n_dec_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


p_alu_in = 0;
p_dec_in = 0;
z_dec_in = 1;
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


z_dec_in = 0;
z_alu_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


/**
The following tests verify that the FSM does not assert branch at the wrong time
**/

//cases when br is not asserted
n_dec_in = 1;
n_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


p_dec_in = 1;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

z_dec_in = 1;
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

//cases when wrong dec asserted
br_in = 1;
n_alu_in = 1;
p_dec_in = 1;
z_dec_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


n_alu_in = 0;
p_dec_in = 0;
n_dec_in = 1;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

p_alu_in = 0;
p_dec_in = 1;
z_alu_in = 1;
z_dec_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

//clear all signals
reset_in = 0;
n_dec_in = 0;
z_dec_in = 0;
p_dec_in = 0;
n_alu_in = 0;
z_alu_in = 0;
p_alu_in = 0;
we_reg_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

//assert reset

reset_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

reset_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

//verify no branches taken in idle

br_in = 1;
n_dec_in = 1;
p_dec_in = 1;
z_dec_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;


















end

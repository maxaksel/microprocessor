magic
tech scmos
timestamp 1682896469
<< polysilicon >>
rect -1464 3339 -1221 3340
rect -1464 2931 3239 3339
rect -1464 2928 3243 2931
rect -1464 -1358 -1221 2928
rect 2996 -1351 3243 2928
<< metal1 >>
rect -1368 4094 -1336 4124
rect -1064 4091 -1026 4122
rect -768 4093 -734 4123
rect -468 4097 -431 4123
rect -173 4089 -116 4133
rect 128 4093 180 4132
rect 422 4091 473 4124
rect 731 4090 780 4127
rect 1034 4095 1080 4129
rect 1329 4097 1378 4128
rect 1638 4094 1679 4129
rect 1925 4098 1982 4132
rect 1931 4096 1972 4098
rect 2227 4097 2273 4132
rect 2525 4095 2583 4127
rect 2838 4101 2869 4125
rect 3130 4093 3181 4131
rect -1493 3385 -1394 3395
rect -1389 3388 -1380 3392
rect -1376 3385 -1248 3394
rect -1493 3372 -1248 3385
rect -1489 3357 -1398 3366
rect -2223 3227 -2201 3273
rect -1495 3221 -1418 3352
rect -1492 3211 -1488 3215
rect -1485 3119 -1418 3221
rect -1414 3135 -1398 3357
rect -1395 3138 -1248 3372
rect -1243 3151 -1234 3389
rect -1230 3383 -1099 3393
rect -1089 3388 -1085 3392
rect -1077 3383 -947 3394
rect -1230 3155 -947 3383
rect -943 3168 -934 3390
rect -931 3384 -794 3393
rect -789 3388 -785 3392
rect -779 3384 -647 3392
rect -931 3172 -647 3384
rect -643 3184 -634 3390
rect -630 3383 -495 3393
rect -489 3388 -485 3392
rect -478 3383 -348 3395
rect -630 3379 -348 3383
rect -629 3189 -348 3379
rect -343 3199 -334 3390
rect -330 3384 -197 3393
rect -189 3388 -185 3393
rect -177 3384 -47 3395
rect -330 3203 -47 3384
rect -43 3214 -34 3390
rect -29 3383 102 3394
rect 111 3388 115 3392
rect 121 3383 253 3394
rect -29 3217 253 3383
rect 257 3229 266 3390
rect 270 3273 395 3391
rect 402 3277 498 3391
rect 506 3379 702 3393
rect 711 3388 715 3392
rect 721 3379 853 3395
rect 506 3375 853 3379
rect 506 3273 742 3375
rect 857 3372 866 3389
rect 873 3385 1007 3393
rect 1011 3388 1015 3392
rect 1020 3385 1153 3394
rect 873 3383 1153 3385
rect 873 3382 1152 3383
rect 270 3232 742 3273
rect 747 3362 866 3372
rect 257 3218 730 3229
rect -43 3203 714 3214
rect -343 3188 698 3199
rect -643 3173 682 3184
rect -943 3157 658 3168
rect -1243 3140 642 3151
rect -1414 3124 626 3135
rect -1485 2997 614 3119
rect -1485 2919 -625 2997
rect -1485 2851 -1212 2919
rect -621 2895 -372 2993
rect -365 2918 614 2997
rect 621 2921 626 3124
rect 637 2921 642 3140
rect 653 2921 658 3157
rect 677 2921 682 3173
rect 693 2921 698 3188
rect 709 2921 714 3203
rect 725 2921 730 3218
rect 747 2920 756 3362
rect 874 3361 1152 3382
rect 1157 3358 1166 3389
rect 1169 3384 1307 3394
rect 1311 3388 1315 3392
rect 1320 3384 1453 3393
rect 1169 3375 1453 3384
rect 763 3347 1166 3358
rect 763 2920 772 3347
rect 1170 3341 1453 3375
rect 1457 3337 1466 3390
rect 1611 3388 1615 3392
rect 779 3329 1466 3337
rect 779 2920 788 3329
rect 1472 3321 1754 3385
rect 1757 3317 1766 3386
rect 795 3309 1766 3317
rect 1772 3384 1906 3394
rect 1911 3388 1915 3392
rect 1919 3384 2053 3394
rect 795 2920 804 3309
rect 1772 3306 2053 3384
rect 2057 3301 2066 3386
rect 2073 3384 2203 3393
rect 2211 3388 2215 3392
rect 2223 3384 2353 3394
rect 2073 3380 2353 3384
rect 811 3293 2068 3301
rect 811 2920 820 3293
rect 2074 3291 2353 3380
rect 2357 3286 2366 3385
rect 827 3275 2366 3286
rect 2371 3275 2496 3392
rect 2502 3276 2598 3392
rect 2811 3388 2815 3392
rect 3111 3388 3115 3392
rect 827 2920 836 3275
rect 2606 3274 2951 3385
rect 2957 3268 2966 3385
rect 843 3259 2966 3268
rect 2970 3259 3175 3384
rect 3257 3375 3266 3384
rect 3178 3367 3266 3375
rect 843 2920 852 3259
rect 3178 3254 3187 3367
rect 3281 3357 3290 3366
rect 859 3246 3187 3254
rect 3204 3349 3290 3357
rect 859 2920 868 3246
rect 3204 3241 3213 3349
rect 875 3233 3213 3241
rect 875 2920 884 3233
rect 3217 3231 3295 3345
rect 3993 3231 4023 3271
rect 891 3218 3262 3226
rect 3267 3218 3295 3231
rect 891 2920 900 3218
rect 904 2918 1456 3215
rect 1461 3206 3228 3213
rect 1461 2924 1466 3206
rect 1469 2919 1514 3203
rect 1517 3194 3207 3201
rect 1517 2924 1522 3194
rect 1525 2919 1530 3190
rect 1533 3182 3191 3189
rect 1533 2924 1538 3182
rect 1541 2920 1592 3179
rect 1597 3172 3158 3179
rect 1597 2924 1602 3172
rect 1605 2920 1720 3168
rect 1725 3162 3146 3169
rect 1725 2924 1730 3162
rect 1735 2919 1886 3157
rect 1893 3151 3134 3158
rect 1893 2924 1898 3151
rect 1901 2919 2081 3147
rect 2085 3140 3122 3147
rect 2085 2924 2090 3140
rect 2095 2989 3111 3136
rect 2095 2988 2637 2989
rect 2095 2919 2609 2988
rect 2619 2895 2889 2982
rect 2895 2921 3111 2989
rect 2995 2852 3111 2921
rect -1485 2765 -1162 2851
rect 2942 2765 3111 2852
rect -1485 2750 -1212 2765
rect 2995 2752 3111 2765
rect -1485 2664 -1162 2750
rect 2943 2665 3111 2752
rect -1485 2651 -1212 2664
rect 2995 2652 3111 2665
rect -1485 2565 -1162 2651
rect 2944 2565 3111 2652
rect -1485 2550 -1212 2565
rect 2995 2552 3111 2565
rect -1485 2464 -1162 2550
rect 2944 2465 3111 2552
rect -1485 2450 -1212 2464
rect 2995 2452 3111 2465
rect -1485 2365 -1162 2450
rect 2944 2365 3111 2452
rect -1485 2349 -1212 2365
rect 2995 2351 3111 2365
rect -1485 2264 -1162 2349
rect 2944 2264 3111 2351
rect -1485 2251 -1212 2264
rect 2995 2252 3111 2264
rect -1485 2166 -1162 2251
rect -1485 2149 -1212 2166
rect 2944 2165 3111 2252
rect 2995 2161 3111 2165
rect 3007 2149 3110 2156
rect -1485 2104 -1162 2149
rect 3007 2119 3098 2126
rect -2224 2022 -2190 2076
rect -1489 2002 -1478 2098
rect -1469 2064 -1162 2104
rect 3007 2099 3087 2106
rect -1469 2049 -1212 2064
rect 2996 2051 3076 2094
rect -1469 2017 -1162 2049
rect -1471 1997 -1162 2017
rect -1484 1964 -1162 1997
rect 2944 1964 3076 2051
rect -1484 1950 -1212 1964
rect 2996 1951 3076 1964
rect -1484 1865 -1162 1950
rect -1484 1851 -1212 1865
rect 2944 1864 3076 1951
rect 2996 1851 3076 1864
rect -1484 1766 -1162 1851
rect -1484 1750 -1212 1766
rect 2943 1764 3076 1851
rect 2996 1751 3076 1764
rect -1484 1665 -1162 1750
rect -1484 1651 -1212 1665
rect 2944 1664 3076 1751
rect 2996 1651 3076 1664
rect -1484 1566 -1162 1651
rect -1484 1550 -1185 1566
rect 2944 1564 3076 1651
rect 2996 1552 3076 1564
rect -1484 1465 -1162 1550
rect 2944 1465 3076 1552
rect -1484 1450 -1212 1465
rect -1484 1365 -1162 1450
rect 2996 1398 3076 1465
rect 3012 1385 3076 1398
rect 2996 1379 3076 1385
rect -1484 1347 -1187 1365
rect 2996 1351 3073 1379
rect -1484 1269 -1162 1347
rect -1489 1257 -1228 1266
rect 2944 1264 3073 1351
rect -2225 1132 -2200 1171
rect -1492 1111 -1488 1115
rect -1485 1105 -1240 1254
rect -1235 1116 -1228 1257
rect 2996 1252 3073 1264
rect -1224 1164 -1162 1251
rect 2944 1165 3073 1252
rect -1224 1151 -1186 1164
rect 2996 1151 3073 1165
rect -1224 1121 -1162 1151
rect -1235 1109 -1221 1116
rect -1210 1105 -1162 1121
rect -1485 1065 -1162 1105
rect 2945 1066 3073 1151
rect -1485 1050 -1210 1065
rect 2996 1051 3073 1066
rect -1485 964 -1162 1050
rect 2945 966 3073 1051
rect -1485 950 -1210 964
rect 2996 950 3073 966
rect -1485 864 -1162 950
rect 2944 865 3073 950
rect -1485 852 -1210 864
rect -1485 764 -1162 852
rect 2996 850 3073 865
rect 2944 765 3073 850
rect -1485 751 -1210 764
rect -1485 665 -1162 751
rect 2996 750 3073 765
rect 2943 665 3073 750
rect -1485 652 -1210 665
rect 2996 652 3073 665
rect -1485 566 -1162 652
rect 2944 567 3073 652
rect -1485 551 -1210 566
rect -1485 465 -1162 551
rect 2996 550 3073 567
rect 2944 465 3073 550
rect -1485 451 -1210 465
rect 2996 452 3073 465
rect -1485 364 -1162 451
rect 2944 367 3073 452
rect -1485 352 -1210 364
rect -1485 312 -1162 352
rect 2996 350 3073 367
rect -2218 233 -2192 265
rect -1489 202 -1480 298
rect -1469 265 -1162 312
rect 2943 265 3073 350
rect -1469 252 -1209 265
rect -1469 195 -1162 252
rect 2996 251 3073 265
rect -1484 165 -1162 195
rect 2944 166 3073 251
rect -1484 152 -1209 165
rect -1484 65 -1162 152
rect 2996 149 3073 166
rect -1484 51 -1209 65
rect 2944 64 3073 149
rect 2996 51 3073 64
rect -1484 -36 -1162 51
rect 2944 -34 3073 51
rect -1484 -48 -1209 -36
rect -1484 -135 -1162 -48
rect 2996 -51 3073 -34
rect -1484 -148 -1209 -135
rect 2944 -136 3073 -51
rect -1484 -235 -1162 -148
rect 2996 -150 3073 -136
rect 2945 -235 3073 -150
rect -1484 -249 -1209 -235
rect -1484 -336 -1162 -249
rect 2996 -250 3073 -235
rect 2944 -335 3073 -250
rect -1484 -349 -1209 -336
rect -1484 -436 -1162 -349
rect 2996 -350 3073 -335
rect 2943 -435 3073 -350
rect -1484 -448 -1209 -436
rect -1484 -535 -1162 -448
rect 2996 -451 3073 -435
rect -1484 -552 -1209 -535
rect 2944 -536 3073 -451
rect 2996 -548 3073 -536
rect -1484 -636 -1162 -552
rect 2944 -633 3073 -548
rect -1484 -649 -1209 -636
rect 2996 -649 3073 -633
rect -1484 -735 -1162 -649
rect 2944 -734 3073 -649
rect -1484 -748 -1209 -735
rect -1484 -834 -1162 -748
rect 2996 -750 3073 -734
rect 2945 -761 3073 -750
rect 3080 -747 3087 2099
rect 3091 -447 3098 2119
rect 3103 153 3110 2149
rect 3115 453 3122 3140
rect 3127 753 3134 3151
rect 3139 1053 3146 3162
rect 3151 1353 3158 3172
rect 3184 2166 3191 3182
rect 3200 2466 3207 3194
rect 3221 2553 3228 3206
rect 3233 3054 3251 3215
rect 3254 3066 3262 3218
rect 3288 3211 3292 3215
rect 3268 3072 3293 3204
rect 3254 3057 3290 3066
rect 3233 3052 3285 3054
rect 3234 2558 3285 3052
rect 3990 2929 4022 2979
rect 3288 2911 3292 2915
rect 3992 2631 4025 2673
rect 3288 2611 3292 2615
rect 3221 2544 3284 2553
rect 3211 2470 3293 2541
rect 3200 2457 3285 2466
rect 3196 2320 3293 2453
rect 3196 2170 3285 2320
rect 3995 2316 4024 2367
rect 3288 2311 3292 2315
rect 3184 2157 3282 2166
rect 3162 1694 3268 2152
rect 4001 2020 4024 2076
rect 3288 2011 3292 2015
rect 3276 1702 3289 1798
rect 3989 1784 4021 1785
rect 3989 1724 4022 1784
rect 3993 1722 4022 1724
rect 3162 1424 3294 1694
rect 3995 1428 4028 1476
rect 3162 1358 3283 1424
rect 3288 1411 3292 1415
rect 3151 1344 3282 1353
rect 3149 1056 3283 1339
rect 3995 1123 4028 1180
rect 3288 1111 3292 1115
rect 3139 1044 3283 1053
rect 3137 758 3284 1041
rect 3992 820 4022 876
rect 3288 811 3292 815
rect 3127 744 3282 753
rect 3126 737 3283 741
rect 3126 457 3284 737
rect 3995 521 4026 576
rect 3288 511 3292 515
rect 3115 444 3282 453
rect 3115 158 3283 438
rect 3985 233 4026 272
rect 3288 211 3292 215
rect 3103 144 3282 153
rect 3102 8 3293 136
rect 3102 -103 3277 8
rect 3283 -98 3289 -2
rect 3987 -70 4024 -20
rect 3102 -381 3294 -103
rect 3995 -376 4026 -319
rect 3102 -443 3277 -381
rect 3288 -389 3292 -385
rect 3091 -456 3283 -447
rect 3091 -743 3280 -462
rect 3995 -676 4029 -614
rect 3288 -689 3292 -685
rect 3080 -756 3282 -747
rect -1484 -855 -1209 -834
rect 2945 -835 3282 -761
rect 2996 -850 3282 -835
rect -1484 -934 -1162 -855
rect -1484 -951 -1209 -934
rect 2944 -935 3282 -850
rect 2996 -950 3282 -935
rect -1484 -1032 -1162 -951
rect -1484 -1053 -1209 -1032
rect 2945 -1035 3282 -950
rect 2996 -1050 3282 -1035
rect -1484 -1134 -1162 -1053
rect -1484 -1204 -1209 -1134
rect 2944 -1135 3282 -1050
rect 2996 -1203 3282 -1135
rect -95 -1204 3284 -1203
rect -1484 -1363 3284 -1204
rect -1484 -1382 -206 -1363
rect -1339 -1383 -206 -1382
rect -198 -1390 -102 -1367
rect -95 -1369 3284 -1363
rect -95 -1384 1588 -1369
rect 1602 -1390 1698 -1374
rect 1703 -1384 3284 -1369
<< metal2 >>
rect -1405 3388 -1401 3392
rect -1477 3378 -1471 3384
rect -1489 3357 -1481 3366
rect -1389 3344 -1380 3392
rect -1243 3381 -1234 3389
rect -1105 3388 -1101 3392
rect -1177 3378 -1171 3383
rect -1089 3379 -1085 3392
rect -943 3381 -934 3390
rect -805 3388 -801 3392
rect -1092 3344 -1082 3379
rect -877 3377 -871 3383
rect -789 3379 -785 3392
rect -643 3381 -634 3390
rect -505 3387 -501 3392
rect -792 3344 -783 3379
rect -577 3378 -571 3384
rect -489 3379 -485 3392
rect -343 3381 -334 3390
rect -205 3388 -201 3392
rect -491 3344 -483 3379
rect -277 3377 -271 3383
rect -189 3379 -185 3393
rect -43 3381 -34 3390
rect 95 3388 99 3392
rect -191 3344 -183 3379
rect 23 3378 29 3383
rect 111 3379 115 3393
rect 257 3381 266 3390
rect 695 3388 699 3393
rect 109 3344 117 3379
rect 402 3344 498 3379
rect 623 3378 629 3383
rect 711 3344 715 3392
rect 857 3381 866 3389
rect 995 3388 999 3392
rect 923 3377 929 3383
rect 1011 3344 1015 3392
rect 1157 3381 1166 3389
rect 1295 3388 1299 3392
rect 1223 3378 1229 3384
rect 1311 3344 1315 3392
rect 1457 3381 1466 3390
rect 1523 3377 1529 3383
rect 1595 3377 1599 3388
rect 1611 3344 1615 3392
rect 1757 3377 1766 3386
rect 1895 3384 1899 3388
rect 1823 3378 1829 3384
rect 1911 3344 1915 3392
rect 2195 3388 2199 3392
rect 2057 3376 2066 3386
rect 2123 3377 2129 3383
rect 2211 3344 2215 3392
rect 2795 3386 2799 3390
rect 2357 3375 2366 3385
rect 2502 3344 2598 3379
rect 2723 3378 2729 3383
rect 2811 3344 2815 3392
rect 3095 3386 3099 3390
rect 2957 3376 2966 3385
rect 3023 3378 3029 3383
rect 3111 3344 3115 3392
rect 3257 3376 3266 3384
rect 3281 3357 3297 3366
rect 3281 3344 3297 3353
rect -1460 3277 3250 3344
rect -1460 3215 -1399 3277
rect -1492 3211 -1399 3215
rect -1492 3195 -1488 3199
rect -1483 3123 -1478 3129
rect -1482 2823 -1476 2829
rect -1482 2523 -1476 2529
rect -1482 2223 -1476 2229
rect -1489 2002 -1467 2098
rect -1489 1257 -1481 1266
rect -1460 1115 -1399 3211
rect -620 2993 -373 3277
rect 2502 3276 2598 3277
rect -621 2895 -372 2993
rect 621 2921 626 3135
rect 637 2921 642 3128
rect 653 2921 658 3128
rect 677 2921 682 3128
rect 693 2921 698 3128
rect 709 2921 714 3128
rect 725 2921 730 3128
rect 2619 2982 2888 3277
rect 3180 3215 3250 3277
rect 3180 3211 3292 3215
rect 747 2920 756 2932
rect 763 2920 772 2932
rect 779 2920 788 2932
rect 795 2920 804 2932
rect 811 2920 820 2932
rect 827 2920 836 2932
rect 843 2920 852 2932
rect 859 2920 868 2932
rect 875 2920 884 2932
rect 891 2920 900 2931
rect 1461 2924 1466 2928
rect 1517 2924 1522 2928
rect 1533 2924 1538 2928
rect 1597 2924 1602 2928
rect 1725 2924 1730 2928
rect 1893 2924 1898 2928
rect 2085 2924 2090 2928
rect 2619 2895 2889 2982
rect 3180 2915 3250 3211
rect 3288 3195 3292 3199
rect 3277 3123 3283 3129
rect 3281 3057 3290 3066
rect 3180 2911 3292 2915
rect 3180 2615 3250 2911
rect 3288 2895 3292 2899
rect 3276 2823 3282 2829
rect 3180 2611 3292 2615
rect 3180 2529 3250 2611
rect 3288 2595 3292 2599
rect 3265 2544 3284 2553
rect 3180 2523 3283 2529
rect 3180 2315 3250 2523
rect 3261 2457 3285 2466
rect 3180 2311 3292 2315
rect 3000 2149 3014 2156
rect 3000 2119 3014 2126
rect 3000 2099 3014 2106
rect 3180 2015 3250 2311
rect 3288 2295 3292 2299
rect 3276 2223 3282 2229
rect 3264 2157 3282 2166
rect 3180 2011 3292 2015
rect 2949 1666 2965 1751
rect 3180 1415 3250 2011
rect 3288 1995 3292 1999
rect 3276 1923 3282 1929
rect 3256 1702 3289 1798
rect 3180 1411 3292 1415
rect 3180 1329 3250 1411
rect 3288 1395 3292 1399
rect 3265 1344 3282 1353
rect 3180 1323 3283 1329
rect -1492 1111 -1399 1115
rect -1492 1095 -1488 1099
rect -1483 1023 -1478 1029
rect -1483 723 -1478 729
rect -1483 423 -1478 429
rect -1489 202 -1471 298
rect -1482 71 -1476 77
rect -1482 -477 -1476 -471
rect -1483 -777 -1477 -771
rect -1483 -1077 -1477 -1071
rect -1460 -1305 -1399 1111
rect -1228 1109 -1214 1116
rect 3180 1115 3250 1323
rect 3180 1111 3292 1115
rect 3180 1029 3250 1111
rect 3288 1095 3292 1099
rect 3265 1044 3283 1053
rect 3180 1023 3283 1029
rect 3180 815 3250 1023
rect 3180 811 3292 815
rect 3180 729 3250 811
rect 3288 795 3292 799
rect 3265 744 3282 753
rect 3180 723 3283 729
rect 3180 515 3250 723
rect 3180 511 3292 515
rect 3180 429 3250 511
rect 3288 495 3292 499
rect 3264 444 3282 453
rect 3180 423 3284 429
rect 3180 215 3250 423
rect 3180 211 3292 215
rect 3180 129 3250 211
rect 3288 195 3292 199
rect 3265 144 3282 153
rect 3180 123 3286 129
rect 2948 -136 2966 -50
rect 3180 -385 3250 123
rect 3277 -98 3289 -2
rect 3180 -389 3292 -385
rect 3180 -471 3250 -389
rect 3288 -405 3292 -401
rect 3265 -456 3283 -447
rect 3180 -477 3286 -471
rect 3180 -685 3250 -477
rect 3180 -689 3292 -685
rect 3180 -771 3250 -689
rect 3288 -705 3292 -701
rect 3265 -756 3282 -747
rect 3180 -777 3283 -771
rect 3180 -1271 3250 -777
rect 3276 -1077 3282 -1071
rect 3179 -1305 3250 -1271
rect -1460 -1345 3250 -1305
rect -1461 -1356 3250 -1345
rect -1482 -1382 -1471 -1371
rect -1177 -1382 -1171 -1376
rect -877 -1382 -871 -1376
rect -577 -1382 -571 -1376
rect -198 -1390 -102 -1356
rect 23 -1382 29 -1376
rect 323 -1382 329 -1376
rect 623 -1382 629 -1376
rect 923 -1382 929 -1376
rect 1223 -1382 1229 -1376
rect 1602 -1390 1698 -1356
rect 1823 -1382 1829 -1376
rect 2123 -1382 2129 -1376
rect 2423 -1382 2429 -1376
rect 2723 -1382 2729 -1376
rect 3023 -1382 3029 -1376
rect 3277 -1377 3283 -1371
<< gv1 >>
rect -1388 3389 -1386 3391
rect -1383 3389 -1381 3391
rect -1088 3389 -1086 3391
rect -788 3389 -786 3391
rect -488 3389 -486 3391
rect -188 3389 -186 3391
rect 112 3389 114 3391
rect 712 3389 714 3391
rect 1012 3389 1014 3391
rect 1312 3389 1314 3391
rect 1612 3389 1614 3391
rect 1912 3389 1914 3391
rect 2212 3389 2214 3391
rect 2812 3389 2814 3391
rect 3112 3389 3114 3391
rect -942 3387 -940 3389
rect -937 3387 -935 3389
rect -642 3387 -640 3389
rect -637 3387 -635 3389
rect -342 3387 -340 3389
rect -337 3387 -335 3389
rect -42 3387 -40 3389
rect -37 3387 -35 3389
rect 258 3387 260 3389
rect 263 3387 265 3389
rect 1458 3387 1460 3389
rect 1463 3387 1465 3389
rect -1242 3384 -1240 3386
rect -1237 3384 -1235 3386
rect 858 3384 860 3386
rect 863 3384 865 3386
rect 1158 3384 1160 3386
rect 1163 3384 1165 3386
rect -942 3382 -940 3384
rect -937 3382 -935 3384
rect -642 3382 -640 3384
rect -637 3382 -635 3384
rect -342 3382 -340 3384
rect -337 3382 -335 3384
rect -42 3382 -40 3384
rect -37 3382 -35 3384
rect 258 3382 260 3384
rect 263 3382 265 3384
rect 1458 3382 1460 3384
rect 1463 3382 1465 3384
rect 1758 3383 1760 3385
rect 1763 3383 1765 3385
rect 2058 3382 2060 3384
rect 2063 3382 2065 3384
rect 2358 3381 2360 3383
rect 2363 3381 2365 3383
rect 2958 3382 2960 3384
rect 2963 3382 2965 3384
rect 1758 3378 1760 3380
rect 1763 3378 1765 3380
rect 3258 3379 3260 3381
rect 3263 3379 3265 3381
rect 2058 3377 2060 3379
rect 2063 3377 2065 3379
rect 2358 3376 2360 3378
rect 2363 3376 2365 3378
rect 2958 3377 2960 3379
rect 2963 3377 2965 3379
rect 404 3374 406 3376
rect 409 3374 411 3376
rect 414 3374 416 3376
rect 419 3374 421 3376
rect 424 3374 426 3376
rect 429 3374 431 3376
rect 434 3374 436 3376
rect 439 3374 441 3376
rect 444 3374 446 3376
rect 449 3374 451 3376
rect 454 3374 456 3376
rect 459 3374 461 3376
rect 464 3374 466 3376
rect 469 3374 471 3376
rect 474 3374 476 3376
rect 479 3374 481 3376
rect 484 3374 486 3376
rect 489 3374 491 3376
rect 494 3374 496 3376
rect 2504 3374 2506 3376
rect 2509 3374 2511 3376
rect 2514 3374 2516 3376
rect 2519 3374 2521 3376
rect 2524 3374 2526 3376
rect 2529 3374 2531 3376
rect 2534 3374 2536 3376
rect 2539 3374 2541 3376
rect 2544 3374 2546 3376
rect 2549 3374 2551 3376
rect 2554 3374 2556 3376
rect 2559 3374 2561 3376
rect 2564 3374 2566 3376
rect 2569 3374 2571 3376
rect 2574 3374 2576 3376
rect 2579 3374 2581 3376
rect 2584 3374 2586 3376
rect 2589 3374 2591 3376
rect 2594 3374 2596 3376
rect 404 3369 406 3371
rect 409 3369 411 3371
rect 414 3369 416 3371
rect 419 3369 421 3371
rect 424 3369 426 3371
rect 429 3369 431 3371
rect 434 3369 436 3371
rect 439 3369 441 3371
rect 444 3369 446 3371
rect 449 3369 451 3371
rect 454 3369 456 3371
rect 459 3369 461 3371
rect 464 3369 466 3371
rect 469 3369 471 3371
rect 474 3369 476 3371
rect 479 3369 481 3371
rect 484 3369 486 3371
rect 489 3369 491 3371
rect 494 3369 496 3371
rect 2504 3369 2506 3371
rect 2509 3369 2511 3371
rect 2514 3369 2516 3371
rect 2519 3369 2521 3371
rect 2524 3369 2526 3371
rect 2529 3369 2531 3371
rect 2534 3369 2536 3371
rect 2539 3369 2541 3371
rect 2544 3369 2546 3371
rect 2549 3369 2551 3371
rect 2554 3369 2556 3371
rect 2559 3369 2561 3371
rect 2564 3369 2566 3371
rect 2569 3369 2571 3371
rect 2574 3369 2576 3371
rect 2579 3369 2581 3371
rect 2584 3369 2586 3371
rect 2589 3369 2591 3371
rect 2594 3369 2596 3371
rect -1486 3363 -1484 3365
rect 404 3364 406 3366
rect 409 3364 411 3366
rect 414 3364 416 3366
rect 419 3364 421 3366
rect 424 3364 426 3366
rect 429 3364 431 3366
rect 434 3364 436 3366
rect 439 3364 441 3366
rect 444 3364 446 3366
rect 449 3364 451 3366
rect 454 3364 456 3366
rect 459 3364 461 3366
rect 464 3364 466 3366
rect 469 3364 471 3366
rect 474 3364 476 3366
rect 479 3364 481 3366
rect 484 3364 486 3366
rect 489 3364 491 3366
rect 494 3364 496 3366
rect 2504 3364 2506 3366
rect 2509 3364 2511 3366
rect 2514 3364 2516 3366
rect 2519 3364 2521 3366
rect 2524 3364 2526 3366
rect 2529 3364 2531 3366
rect 2534 3364 2536 3366
rect 2539 3364 2541 3366
rect 2544 3364 2546 3366
rect 2549 3364 2551 3366
rect 2554 3364 2556 3366
rect 2559 3364 2561 3366
rect 2564 3364 2566 3366
rect 2569 3364 2571 3366
rect 2574 3364 2576 3366
rect 2579 3364 2581 3366
rect 2584 3364 2586 3366
rect 2589 3364 2591 3366
rect 2594 3364 2596 3366
rect 3282 3363 3284 3365
rect 3287 3363 3289 3365
rect -1486 3358 -1484 3360
rect 404 3359 406 3361
rect 409 3359 411 3361
rect 414 3359 416 3361
rect 419 3359 421 3361
rect 424 3359 426 3361
rect 429 3359 431 3361
rect 434 3359 436 3361
rect 439 3359 441 3361
rect 444 3359 446 3361
rect 449 3359 451 3361
rect 454 3359 456 3361
rect 459 3359 461 3361
rect 464 3359 466 3361
rect 469 3359 471 3361
rect 474 3359 476 3361
rect 479 3359 481 3361
rect 484 3359 486 3361
rect 489 3359 491 3361
rect 494 3359 496 3361
rect 2504 3359 2506 3361
rect 2509 3359 2511 3361
rect 2514 3359 2516 3361
rect 2519 3359 2521 3361
rect 2524 3359 2526 3361
rect 2529 3359 2531 3361
rect 2534 3359 2536 3361
rect 2539 3359 2541 3361
rect 2544 3359 2546 3361
rect 2549 3359 2551 3361
rect 2554 3359 2556 3361
rect 2559 3359 2561 3361
rect 2564 3359 2566 3361
rect 2569 3359 2571 3361
rect 2574 3359 2576 3361
rect 2579 3359 2581 3361
rect 2584 3359 2586 3361
rect 2589 3359 2591 3361
rect 2594 3359 2596 3361
rect 3282 3358 3284 3360
rect 3287 3358 3289 3360
rect 404 3354 406 3356
rect 409 3354 411 3356
rect 414 3354 416 3356
rect 419 3354 421 3356
rect 424 3354 426 3356
rect 429 3354 431 3356
rect 434 3354 436 3356
rect 439 3354 441 3356
rect 444 3354 446 3356
rect 449 3354 451 3356
rect 454 3354 456 3356
rect 459 3354 461 3356
rect 464 3354 466 3356
rect 469 3354 471 3356
rect 474 3354 476 3356
rect 479 3354 481 3356
rect 484 3354 486 3356
rect 489 3354 491 3356
rect 494 3354 496 3356
rect 2504 3354 2506 3356
rect 2509 3354 2511 3356
rect 2514 3354 2516 3356
rect 2519 3354 2521 3356
rect 2524 3354 2526 3356
rect 2529 3354 2531 3356
rect 2534 3354 2536 3356
rect 2539 3354 2541 3356
rect 2544 3354 2546 3356
rect 2549 3354 2551 3356
rect 2554 3354 2556 3356
rect 2559 3354 2561 3356
rect 2564 3354 2566 3356
rect 2569 3354 2571 3356
rect 2574 3354 2576 3356
rect 2579 3354 2581 3356
rect 2584 3354 2586 3356
rect 2589 3354 2591 3356
rect 2594 3354 2596 3356
rect 404 3349 406 3351
rect 409 3349 411 3351
rect 414 3349 416 3351
rect 419 3349 421 3351
rect 424 3349 426 3351
rect 429 3349 431 3351
rect 434 3349 436 3351
rect 439 3349 441 3351
rect 444 3349 446 3351
rect 449 3349 451 3351
rect 454 3349 456 3351
rect 459 3349 461 3351
rect 464 3349 466 3351
rect 469 3349 471 3351
rect 474 3349 476 3351
rect 479 3349 481 3351
rect 484 3349 486 3351
rect 489 3349 491 3351
rect 494 3349 496 3351
rect 2504 3349 2506 3351
rect 2509 3349 2511 3351
rect 2514 3349 2516 3351
rect 2519 3349 2521 3351
rect 2524 3349 2526 3351
rect 2529 3349 2531 3351
rect 2534 3349 2536 3351
rect 2539 3349 2541 3351
rect 2544 3349 2546 3351
rect 2549 3349 2551 3351
rect 2554 3349 2556 3351
rect 2559 3349 2561 3351
rect 2564 3349 2566 3351
rect 2569 3349 2571 3351
rect 2574 3349 2576 3351
rect 2579 3349 2581 3351
rect 2584 3349 2586 3351
rect 2589 3349 2591 3351
rect 2594 3349 2596 3351
rect 404 3344 406 3346
rect 409 3344 411 3346
rect 414 3344 416 3346
rect 419 3344 421 3346
rect 424 3344 426 3346
rect 429 3344 431 3346
rect 434 3344 436 3346
rect 439 3344 441 3346
rect 444 3344 446 3346
rect 449 3344 451 3346
rect 454 3344 456 3346
rect 459 3344 461 3346
rect 464 3344 466 3346
rect 469 3344 471 3346
rect 474 3344 476 3346
rect 479 3344 481 3346
rect 484 3344 486 3346
rect 489 3344 491 3346
rect 494 3344 496 3346
rect 2504 3344 2506 3346
rect 2509 3344 2511 3346
rect 2514 3344 2516 3346
rect 2519 3344 2521 3346
rect 2524 3344 2526 3346
rect 2529 3344 2531 3346
rect 2534 3344 2536 3346
rect 2539 3344 2541 3346
rect 2544 3344 2546 3346
rect 2549 3344 2551 3346
rect 2554 3344 2556 3346
rect 2559 3344 2561 3346
rect 2564 3344 2566 3346
rect 2569 3344 2571 3346
rect 2574 3344 2576 3346
rect 2579 3344 2581 3346
rect 2584 3344 2586 3346
rect 2589 3344 2591 3346
rect 2594 3344 2596 3346
rect 404 3339 406 3341
rect 409 3339 411 3341
rect 414 3339 416 3341
rect 419 3339 421 3341
rect 424 3339 426 3341
rect 429 3339 431 3341
rect 434 3339 436 3341
rect 439 3339 441 3341
rect 444 3339 446 3341
rect 449 3339 451 3341
rect 454 3339 456 3341
rect 459 3339 461 3341
rect 464 3339 466 3341
rect 469 3339 471 3341
rect 474 3339 476 3341
rect 479 3339 481 3341
rect 484 3339 486 3341
rect 489 3339 491 3341
rect 494 3339 496 3341
rect 2504 3339 2506 3341
rect 2509 3339 2511 3341
rect 2514 3339 2516 3341
rect 2519 3339 2521 3341
rect 2524 3339 2526 3341
rect 2529 3339 2531 3341
rect 2534 3339 2536 3341
rect 2539 3339 2541 3341
rect 2544 3339 2546 3341
rect 2549 3339 2551 3341
rect 2554 3339 2556 3341
rect 2559 3339 2561 3341
rect 2564 3339 2566 3341
rect 2569 3339 2571 3341
rect 2574 3339 2576 3341
rect 2579 3339 2581 3341
rect 2584 3339 2586 3341
rect 2589 3339 2591 3341
rect 2594 3339 2596 3341
rect 404 3334 406 3336
rect 409 3334 411 3336
rect 414 3334 416 3336
rect 419 3334 421 3336
rect 424 3334 426 3336
rect 429 3334 431 3336
rect 434 3334 436 3336
rect 439 3334 441 3336
rect 444 3334 446 3336
rect 449 3334 451 3336
rect 454 3334 456 3336
rect 459 3334 461 3336
rect 464 3334 466 3336
rect 469 3334 471 3336
rect 474 3334 476 3336
rect 479 3334 481 3336
rect 484 3334 486 3336
rect 489 3334 491 3336
rect 494 3334 496 3336
rect 2504 3334 2506 3336
rect 2509 3334 2511 3336
rect 2514 3334 2516 3336
rect 2519 3334 2521 3336
rect 2524 3334 2526 3336
rect 2529 3334 2531 3336
rect 2534 3334 2536 3336
rect 2539 3334 2541 3336
rect 2544 3334 2546 3336
rect 2549 3334 2551 3336
rect 2554 3334 2556 3336
rect 2559 3334 2561 3336
rect 2564 3334 2566 3336
rect 2569 3334 2571 3336
rect 2574 3334 2576 3336
rect 2579 3334 2581 3336
rect 2584 3334 2586 3336
rect 2589 3334 2591 3336
rect 2594 3334 2596 3336
rect 404 3329 406 3331
rect 409 3329 411 3331
rect 414 3329 416 3331
rect 419 3329 421 3331
rect 424 3329 426 3331
rect 429 3329 431 3331
rect 434 3329 436 3331
rect 439 3329 441 3331
rect 444 3329 446 3331
rect 449 3329 451 3331
rect 454 3329 456 3331
rect 459 3329 461 3331
rect 464 3329 466 3331
rect 469 3329 471 3331
rect 474 3329 476 3331
rect 479 3329 481 3331
rect 484 3329 486 3331
rect 489 3329 491 3331
rect 494 3329 496 3331
rect 2504 3329 2506 3331
rect 2509 3329 2511 3331
rect 2514 3329 2516 3331
rect 2519 3329 2521 3331
rect 2524 3329 2526 3331
rect 2529 3329 2531 3331
rect 2534 3329 2536 3331
rect 2539 3329 2541 3331
rect 2544 3329 2546 3331
rect 2549 3329 2551 3331
rect 2554 3329 2556 3331
rect 2559 3329 2561 3331
rect 2564 3329 2566 3331
rect 2569 3329 2571 3331
rect 2574 3329 2576 3331
rect 2579 3329 2581 3331
rect 2584 3329 2586 3331
rect 2589 3329 2591 3331
rect 2594 3329 2596 3331
rect 404 3324 406 3326
rect 409 3324 411 3326
rect 414 3324 416 3326
rect 419 3324 421 3326
rect 424 3324 426 3326
rect 429 3324 431 3326
rect 434 3324 436 3326
rect 439 3324 441 3326
rect 444 3324 446 3326
rect 449 3324 451 3326
rect 454 3324 456 3326
rect 459 3324 461 3326
rect 464 3324 466 3326
rect 469 3324 471 3326
rect 474 3324 476 3326
rect 479 3324 481 3326
rect 484 3324 486 3326
rect 489 3324 491 3326
rect 494 3324 496 3326
rect 2504 3324 2506 3326
rect 2509 3324 2511 3326
rect 2514 3324 2516 3326
rect 2519 3324 2521 3326
rect 2524 3324 2526 3326
rect 2529 3324 2531 3326
rect 2534 3324 2536 3326
rect 2539 3324 2541 3326
rect 2544 3324 2546 3326
rect 2549 3324 2551 3326
rect 2554 3324 2556 3326
rect 2559 3324 2561 3326
rect 2564 3324 2566 3326
rect 2569 3324 2571 3326
rect 2574 3324 2576 3326
rect 2579 3324 2581 3326
rect 2584 3324 2586 3326
rect 2589 3324 2591 3326
rect 2594 3324 2596 3326
rect 404 3319 406 3321
rect 409 3319 411 3321
rect 414 3319 416 3321
rect 419 3319 421 3321
rect 424 3319 426 3321
rect 429 3319 431 3321
rect 434 3319 436 3321
rect 439 3319 441 3321
rect 444 3319 446 3321
rect 449 3319 451 3321
rect 454 3319 456 3321
rect 459 3319 461 3321
rect 464 3319 466 3321
rect 469 3319 471 3321
rect 474 3319 476 3321
rect 479 3319 481 3321
rect 484 3319 486 3321
rect 489 3319 491 3321
rect 494 3319 496 3321
rect 2504 3319 2506 3321
rect 2509 3319 2511 3321
rect 2514 3319 2516 3321
rect 2519 3319 2521 3321
rect 2524 3319 2526 3321
rect 2529 3319 2531 3321
rect 2534 3319 2536 3321
rect 2539 3319 2541 3321
rect 2544 3319 2546 3321
rect 2549 3319 2551 3321
rect 2554 3319 2556 3321
rect 2559 3319 2561 3321
rect 2564 3319 2566 3321
rect 2569 3319 2571 3321
rect 2574 3319 2576 3321
rect 2579 3319 2581 3321
rect 2584 3319 2586 3321
rect 2589 3319 2591 3321
rect 2594 3319 2596 3321
rect 404 3314 406 3316
rect 409 3314 411 3316
rect 414 3314 416 3316
rect 419 3314 421 3316
rect 424 3314 426 3316
rect 429 3314 431 3316
rect 434 3314 436 3316
rect 439 3314 441 3316
rect 444 3314 446 3316
rect 449 3314 451 3316
rect 454 3314 456 3316
rect 459 3314 461 3316
rect 464 3314 466 3316
rect 469 3314 471 3316
rect 474 3314 476 3316
rect 479 3314 481 3316
rect 484 3314 486 3316
rect 489 3314 491 3316
rect 494 3314 496 3316
rect 2504 3314 2506 3316
rect 2509 3314 2511 3316
rect 2514 3314 2516 3316
rect 2519 3314 2521 3316
rect 2524 3314 2526 3316
rect 2529 3314 2531 3316
rect 2534 3314 2536 3316
rect 2539 3314 2541 3316
rect 2544 3314 2546 3316
rect 2549 3314 2551 3316
rect 2554 3314 2556 3316
rect 2559 3314 2561 3316
rect 2564 3314 2566 3316
rect 2569 3314 2571 3316
rect 2574 3314 2576 3316
rect 2579 3314 2581 3316
rect 2584 3314 2586 3316
rect 2589 3314 2591 3316
rect 2594 3314 2596 3316
rect 404 3309 406 3311
rect 409 3309 411 3311
rect 414 3309 416 3311
rect 419 3309 421 3311
rect 424 3309 426 3311
rect 429 3309 431 3311
rect 434 3309 436 3311
rect 439 3309 441 3311
rect 444 3309 446 3311
rect 449 3309 451 3311
rect 454 3309 456 3311
rect 459 3309 461 3311
rect 464 3309 466 3311
rect 469 3309 471 3311
rect 474 3309 476 3311
rect 479 3309 481 3311
rect 484 3309 486 3311
rect 489 3309 491 3311
rect 494 3309 496 3311
rect 2504 3309 2506 3311
rect 2509 3309 2511 3311
rect 2514 3309 2516 3311
rect 2519 3309 2521 3311
rect 2524 3309 2526 3311
rect 2529 3309 2531 3311
rect 2534 3309 2536 3311
rect 2539 3309 2541 3311
rect 2544 3309 2546 3311
rect 2549 3309 2551 3311
rect 2554 3309 2556 3311
rect 2559 3309 2561 3311
rect 2564 3309 2566 3311
rect 2569 3309 2571 3311
rect 2574 3309 2576 3311
rect 2579 3309 2581 3311
rect 2584 3309 2586 3311
rect 2589 3309 2591 3311
rect 2594 3309 2596 3311
rect 404 3304 406 3306
rect 409 3304 411 3306
rect 414 3304 416 3306
rect 419 3304 421 3306
rect 424 3304 426 3306
rect 429 3304 431 3306
rect 434 3304 436 3306
rect 439 3304 441 3306
rect 444 3304 446 3306
rect 449 3304 451 3306
rect 454 3304 456 3306
rect 459 3304 461 3306
rect 464 3304 466 3306
rect 469 3304 471 3306
rect 474 3304 476 3306
rect 479 3304 481 3306
rect 484 3304 486 3306
rect 489 3304 491 3306
rect 494 3304 496 3306
rect 2504 3304 2506 3306
rect 2509 3304 2511 3306
rect 2514 3304 2516 3306
rect 2519 3304 2521 3306
rect 2524 3304 2526 3306
rect 2529 3304 2531 3306
rect 2534 3304 2536 3306
rect 2539 3304 2541 3306
rect 2544 3304 2546 3306
rect 2549 3304 2551 3306
rect 2554 3304 2556 3306
rect 2559 3304 2561 3306
rect 2564 3304 2566 3306
rect 2569 3304 2571 3306
rect 2574 3304 2576 3306
rect 2579 3304 2581 3306
rect 2584 3304 2586 3306
rect 2589 3304 2591 3306
rect 2594 3304 2596 3306
rect 404 3299 406 3301
rect 409 3299 411 3301
rect 414 3299 416 3301
rect 419 3299 421 3301
rect 424 3299 426 3301
rect 429 3299 431 3301
rect 434 3299 436 3301
rect 439 3299 441 3301
rect 444 3299 446 3301
rect 449 3299 451 3301
rect 454 3299 456 3301
rect 459 3299 461 3301
rect 464 3299 466 3301
rect 469 3299 471 3301
rect 474 3299 476 3301
rect 479 3299 481 3301
rect 484 3299 486 3301
rect 489 3299 491 3301
rect 494 3299 496 3301
rect 2504 3299 2506 3301
rect 2509 3299 2511 3301
rect 2514 3299 2516 3301
rect 2519 3299 2521 3301
rect 2524 3299 2526 3301
rect 2529 3299 2531 3301
rect 2534 3299 2536 3301
rect 2539 3299 2541 3301
rect 2544 3299 2546 3301
rect 2549 3299 2551 3301
rect 2554 3299 2556 3301
rect 2559 3299 2561 3301
rect 2564 3299 2566 3301
rect 2569 3299 2571 3301
rect 2574 3299 2576 3301
rect 2579 3299 2581 3301
rect 2584 3299 2586 3301
rect 2589 3299 2591 3301
rect 2594 3299 2596 3301
rect 404 3294 406 3296
rect 409 3294 411 3296
rect 414 3294 416 3296
rect 419 3294 421 3296
rect 424 3294 426 3296
rect 429 3294 431 3296
rect 434 3294 436 3296
rect 439 3294 441 3296
rect 444 3294 446 3296
rect 449 3294 451 3296
rect 454 3294 456 3296
rect 459 3294 461 3296
rect 464 3294 466 3296
rect 469 3294 471 3296
rect 474 3294 476 3296
rect 479 3294 481 3296
rect 484 3294 486 3296
rect 489 3294 491 3296
rect 494 3294 496 3296
rect 2504 3294 2506 3296
rect 2509 3294 2511 3296
rect 2514 3294 2516 3296
rect 2519 3294 2521 3296
rect 2524 3294 2526 3296
rect 2529 3294 2531 3296
rect 2534 3294 2536 3296
rect 2539 3294 2541 3296
rect 2544 3294 2546 3296
rect 2549 3294 2551 3296
rect 2554 3294 2556 3296
rect 2559 3294 2561 3296
rect 2564 3294 2566 3296
rect 2569 3294 2571 3296
rect 2574 3294 2576 3296
rect 2579 3294 2581 3296
rect 2584 3294 2586 3296
rect 2589 3294 2591 3296
rect 2594 3294 2596 3296
rect 404 3289 406 3291
rect 409 3289 411 3291
rect 414 3289 416 3291
rect 419 3289 421 3291
rect 424 3289 426 3291
rect 429 3289 431 3291
rect 434 3289 436 3291
rect 439 3289 441 3291
rect 444 3289 446 3291
rect 449 3289 451 3291
rect 454 3289 456 3291
rect 459 3289 461 3291
rect 464 3289 466 3291
rect 469 3289 471 3291
rect 474 3289 476 3291
rect 479 3289 481 3291
rect 484 3289 486 3291
rect 489 3289 491 3291
rect 494 3289 496 3291
rect 2504 3289 2506 3291
rect 2509 3289 2511 3291
rect 2514 3289 2516 3291
rect 2519 3289 2521 3291
rect 2524 3289 2526 3291
rect 2529 3289 2531 3291
rect 2534 3289 2536 3291
rect 2539 3289 2541 3291
rect 2544 3289 2546 3291
rect 2549 3289 2551 3291
rect 2554 3289 2556 3291
rect 2559 3289 2561 3291
rect 2564 3289 2566 3291
rect 2569 3289 2571 3291
rect 2574 3289 2576 3291
rect 2579 3289 2581 3291
rect 2584 3289 2586 3291
rect 2589 3289 2591 3291
rect 2594 3289 2596 3291
rect 404 3284 406 3286
rect 409 3284 411 3286
rect 414 3284 416 3286
rect 419 3284 421 3286
rect 424 3284 426 3286
rect 429 3284 431 3286
rect 434 3284 436 3286
rect 439 3284 441 3286
rect 444 3284 446 3286
rect 449 3284 451 3286
rect 454 3284 456 3286
rect 459 3284 461 3286
rect 464 3284 466 3286
rect 469 3284 471 3286
rect 474 3284 476 3286
rect 479 3284 481 3286
rect 484 3284 486 3286
rect 489 3284 491 3286
rect 494 3284 496 3286
rect 2504 3284 2506 3286
rect 2509 3284 2511 3286
rect 2514 3284 2516 3286
rect 2519 3284 2521 3286
rect 2524 3284 2526 3286
rect 2529 3284 2531 3286
rect 2534 3284 2536 3286
rect 2539 3284 2541 3286
rect 2544 3284 2546 3286
rect 2549 3284 2551 3286
rect 2554 3284 2556 3286
rect 2559 3284 2561 3286
rect 2564 3284 2566 3286
rect 2569 3284 2571 3286
rect 2574 3284 2576 3286
rect 2579 3284 2581 3286
rect 2584 3284 2586 3286
rect 2589 3284 2591 3286
rect 2594 3284 2596 3286
rect 404 3279 406 3281
rect 409 3279 411 3281
rect 414 3279 416 3281
rect 419 3279 421 3281
rect 424 3279 426 3281
rect 429 3279 431 3281
rect 434 3279 436 3281
rect 439 3279 441 3281
rect 444 3279 446 3281
rect 449 3279 451 3281
rect 454 3279 456 3281
rect 459 3279 461 3281
rect 464 3279 466 3281
rect 469 3279 471 3281
rect 474 3279 476 3281
rect 479 3279 481 3281
rect 484 3279 486 3281
rect 489 3279 491 3281
rect 494 3279 496 3281
rect 2504 3279 2506 3281
rect 2509 3279 2511 3281
rect 2514 3279 2516 3281
rect 2519 3279 2521 3281
rect 2524 3279 2526 3281
rect 2529 3279 2531 3281
rect 2534 3279 2536 3281
rect 2539 3279 2541 3281
rect 2544 3279 2546 3281
rect 2549 3279 2551 3281
rect 2554 3279 2556 3281
rect 2559 3279 2561 3281
rect 2564 3279 2566 3281
rect 2569 3279 2571 3281
rect 2574 3279 2576 3281
rect 2579 3279 2581 3281
rect 2584 3279 2586 3281
rect 2589 3279 2591 3281
rect 2594 3279 2596 3281
rect -1491 3212 -1489 3214
rect 3289 3212 3291 3214
rect 622 3132 624 3134
rect 622 3127 624 3129
rect 622 3122 624 3124
rect 638 3123 640 3125
rect 654 3123 656 3125
rect 678 3123 680 3125
rect 694 3123 696 3125
rect 710 3123 712 3125
rect 726 3123 728 3125
rect 622 3117 624 3119
rect 638 3118 640 3120
rect 654 3118 656 3120
rect 678 3118 680 3120
rect 694 3118 696 3120
rect 710 3118 712 3120
rect 726 3118 728 3120
rect 622 3112 624 3114
rect 638 3113 640 3115
rect 654 3113 656 3115
rect 678 3113 680 3115
rect 694 3113 696 3115
rect 710 3113 712 3115
rect 726 3113 728 3115
rect 622 3107 624 3109
rect 638 3108 640 3110
rect 654 3108 656 3110
rect 678 3108 680 3110
rect 694 3108 696 3110
rect 710 3108 712 3110
rect 726 3108 728 3110
rect 622 3102 624 3104
rect 638 3103 640 3105
rect 654 3103 656 3105
rect 678 3103 680 3105
rect 694 3103 696 3105
rect 710 3103 712 3105
rect 726 3103 728 3105
rect 622 3097 624 3099
rect 638 3098 640 3100
rect 654 3098 656 3100
rect 678 3098 680 3100
rect 694 3098 696 3100
rect 710 3098 712 3100
rect 726 3098 728 3100
rect 622 3092 624 3094
rect 638 3093 640 3095
rect 654 3093 656 3095
rect 678 3093 680 3095
rect 694 3093 696 3095
rect 710 3093 712 3095
rect 726 3093 728 3095
rect 622 3087 624 3089
rect 638 3088 640 3090
rect 654 3088 656 3090
rect 678 3088 680 3090
rect 694 3088 696 3090
rect 710 3088 712 3090
rect 726 3088 728 3090
rect 622 3082 624 3084
rect 638 3083 640 3085
rect 654 3083 656 3085
rect 678 3083 680 3085
rect 694 3083 696 3085
rect 710 3083 712 3085
rect 726 3083 728 3085
rect 622 3077 624 3079
rect 638 3078 640 3080
rect 654 3078 656 3080
rect 678 3078 680 3080
rect 694 3078 696 3080
rect 710 3078 712 3080
rect 726 3078 728 3080
rect 622 3072 624 3074
rect 638 3073 640 3075
rect 654 3073 656 3075
rect 678 3073 680 3075
rect 694 3073 696 3075
rect 710 3073 712 3075
rect 726 3073 728 3075
rect 622 3067 624 3069
rect 638 3068 640 3070
rect 654 3068 656 3070
rect 678 3068 680 3070
rect 694 3068 696 3070
rect 710 3068 712 3070
rect 726 3068 728 3070
rect 622 3062 624 3064
rect 638 3063 640 3065
rect 654 3063 656 3065
rect 678 3063 680 3065
rect 694 3063 696 3065
rect 710 3063 712 3065
rect 726 3063 728 3065
rect 3282 3063 3284 3065
rect 3287 3063 3289 3065
rect 622 3057 624 3059
rect 638 3058 640 3060
rect 654 3058 656 3060
rect 678 3058 680 3060
rect 694 3058 696 3060
rect 710 3058 712 3060
rect 726 3058 728 3060
rect 3282 3058 3284 3060
rect 3287 3058 3289 3060
rect 622 3052 624 3054
rect 638 3053 640 3055
rect 654 3053 656 3055
rect 678 3053 680 3055
rect 694 3053 696 3055
rect 710 3053 712 3055
rect 726 3053 728 3055
rect 622 3047 624 3049
rect 638 3048 640 3050
rect 654 3048 656 3050
rect 678 3048 680 3050
rect 694 3048 696 3050
rect 710 3048 712 3050
rect 726 3048 728 3050
rect 622 3042 624 3044
rect 638 3043 640 3045
rect 654 3043 656 3045
rect 678 3043 680 3045
rect 694 3043 696 3045
rect 710 3043 712 3045
rect 726 3043 728 3045
rect 622 3037 624 3039
rect 638 3038 640 3040
rect 654 3038 656 3040
rect 678 3038 680 3040
rect 694 3038 696 3040
rect 710 3038 712 3040
rect 726 3038 728 3040
rect 622 3032 624 3034
rect 638 3033 640 3035
rect 654 3033 656 3035
rect 678 3033 680 3035
rect 694 3033 696 3035
rect 710 3033 712 3035
rect 726 3033 728 3035
rect 622 3027 624 3029
rect 638 3028 640 3030
rect 654 3028 656 3030
rect 678 3028 680 3030
rect 694 3028 696 3030
rect 710 3028 712 3030
rect 726 3028 728 3030
rect 622 3022 624 3024
rect 638 3023 640 3025
rect 654 3023 656 3025
rect 678 3023 680 3025
rect 694 3023 696 3025
rect 710 3023 712 3025
rect 726 3023 728 3025
rect 622 3017 624 3019
rect 638 3018 640 3020
rect 654 3018 656 3020
rect 678 3018 680 3020
rect 694 3018 696 3020
rect 710 3018 712 3020
rect 726 3018 728 3020
rect 622 3012 624 3014
rect 638 3013 640 3015
rect 654 3013 656 3015
rect 678 3013 680 3015
rect 694 3013 696 3015
rect 710 3013 712 3015
rect 726 3013 728 3015
rect 622 3007 624 3009
rect 638 3008 640 3010
rect 654 3008 656 3010
rect 678 3008 680 3010
rect 694 3008 696 3010
rect 710 3008 712 3010
rect 726 3008 728 3010
rect 622 3002 624 3004
rect 638 3003 640 3005
rect 654 3003 656 3005
rect 678 3003 680 3005
rect 694 3003 696 3005
rect 710 3003 712 3005
rect 726 3003 728 3005
rect 622 2997 624 2999
rect 638 2998 640 3000
rect 654 2998 656 3000
rect 678 2998 680 3000
rect 694 2998 696 3000
rect 710 2998 712 3000
rect 726 2998 728 3000
rect 622 2992 624 2994
rect 638 2993 640 2995
rect 654 2993 656 2995
rect 678 2993 680 2995
rect 694 2993 696 2995
rect 710 2993 712 2995
rect 726 2993 728 2995
rect -620 2988 -618 2990
rect -615 2988 -613 2990
rect -610 2988 -608 2990
rect -605 2988 -603 2990
rect -600 2988 -598 2990
rect -595 2988 -593 2990
rect -590 2988 -588 2990
rect -585 2988 -583 2990
rect -580 2988 -578 2990
rect -575 2988 -573 2990
rect -570 2988 -568 2990
rect -565 2988 -563 2990
rect -560 2988 -558 2990
rect -555 2988 -553 2990
rect -550 2988 -548 2990
rect -545 2988 -543 2990
rect -540 2988 -538 2990
rect -535 2988 -533 2990
rect -530 2988 -528 2990
rect -525 2988 -523 2990
rect -520 2988 -518 2990
rect -515 2988 -513 2990
rect -510 2988 -508 2990
rect -505 2988 -503 2990
rect -500 2988 -498 2990
rect -495 2988 -493 2990
rect -490 2988 -488 2990
rect -485 2988 -483 2990
rect -480 2988 -478 2990
rect -475 2988 -473 2990
rect -470 2988 -468 2990
rect -465 2988 -463 2990
rect -460 2988 -458 2990
rect -455 2988 -453 2990
rect -450 2988 -448 2990
rect -445 2988 -443 2990
rect -440 2988 -438 2990
rect -435 2988 -433 2990
rect -430 2988 -428 2990
rect -425 2988 -423 2990
rect -420 2988 -418 2990
rect -415 2988 -413 2990
rect -410 2988 -408 2990
rect -405 2988 -403 2990
rect -400 2988 -398 2990
rect -395 2988 -393 2990
rect -390 2988 -388 2990
rect -385 2988 -383 2990
rect -380 2988 -378 2990
rect -375 2988 -373 2990
rect 622 2987 624 2989
rect 638 2988 640 2990
rect 654 2988 656 2990
rect 678 2988 680 2990
rect 694 2988 696 2990
rect 710 2988 712 2990
rect 726 2988 728 2990
rect -620 2983 -618 2985
rect -615 2983 -613 2985
rect -610 2983 -608 2985
rect -605 2983 -603 2985
rect -600 2983 -598 2985
rect -595 2983 -593 2985
rect -590 2983 -588 2985
rect -585 2983 -583 2985
rect -580 2983 -578 2985
rect -575 2983 -573 2985
rect -570 2983 -568 2985
rect -565 2983 -563 2985
rect -560 2983 -558 2985
rect -555 2983 -553 2985
rect -550 2983 -548 2985
rect -545 2983 -543 2985
rect -540 2983 -538 2985
rect -535 2983 -533 2985
rect -530 2983 -528 2985
rect -525 2983 -523 2985
rect -520 2983 -518 2985
rect -515 2983 -513 2985
rect -510 2983 -508 2985
rect -505 2983 -503 2985
rect -500 2983 -498 2985
rect -495 2983 -493 2985
rect -490 2983 -488 2985
rect -485 2983 -483 2985
rect -480 2983 -478 2985
rect -475 2983 -473 2985
rect -470 2983 -468 2985
rect -465 2983 -463 2985
rect -460 2983 -458 2985
rect -455 2983 -453 2985
rect -450 2983 -448 2985
rect -445 2983 -443 2985
rect -440 2983 -438 2985
rect -435 2983 -433 2985
rect -430 2983 -428 2985
rect -425 2983 -423 2985
rect -420 2983 -418 2985
rect -415 2983 -413 2985
rect -410 2983 -408 2985
rect -405 2983 -403 2985
rect -400 2983 -398 2985
rect -395 2983 -393 2985
rect -390 2983 -388 2985
rect -385 2983 -383 2985
rect -380 2983 -378 2985
rect -375 2983 -373 2985
rect 622 2982 624 2984
rect 638 2983 640 2985
rect 654 2983 656 2985
rect 678 2983 680 2985
rect 694 2983 696 2985
rect 710 2983 712 2985
rect 726 2983 728 2985
rect -620 2978 -618 2980
rect -615 2978 -613 2980
rect -610 2978 -608 2980
rect -605 2978 -603 2980
rect -600 2978 -598 2980
rect -595 2978 -593 2980
rect -590 2978 -588 2980
rect -585 2978 -583 2980
rect -580 2978 -578 2980
rect -575 2978 -573 2980
rect -570 2978 -568 2980
rect -565 2978 -563 2980
rect -560 2978 -558 2980
rect -555 2978 -553 2980
rect -550 2978 -548 2980
rect -545 2978 -543 2980
rect -540 2978 -538 2980
rect -535 2978 -533 2980
rect -530 2978 -528 2980
rect -525 2978 -523 2980
rect -520 2978 -518 2980
rect -515 2978 -513 2980
rect -510 2978 -508 2980
rect -505 2978 -503 2980
rect -500 2978 -498 2980
rect -495 2978 -493 2980
rect -490 2978 -488 2980
rect -485 2978 -483 2980
rect -480 2978 -478 2980
rect -475 2978 -473 2980
rect -470 2978 -468 2980
rect -465 2978 -463 2980
rect -460 2978 -458 2980
rect -455 2978 -453 2980
rect -450 2978 -448 2980
rect -445 2978 -443 2980
rect -440 2978 -438 2980
rect -435 2978 -433 2980
rect -430 2978 -428 2980
rect -425 2978 -423 2980
rect -420 2978 -418 2980
rect -415 2978 -413 2980
rect -410 2978 -408 2980
rect -405 2978 -403 2980
rect -400 2978 -398 2980
rect -395 2978 -393 2980
rect -390 2978 -388 2980
rect -385 2978 -383 2980
rect -380 2978 -378 2980
rect -375 2978 -373 2980
rect 622 2977 624 2979
rect 638 2978 640 2980
rect 654 2978 656 2980
rect 678 2978 680 2980
rect 694 2978 696 2980
rect 710 2978 712 2980
rect 726 2978 728 2980
rect 2620 2977 2622 2979
rect 2625 2977 2627 2979
rect 2630 2977 2632 2979
rect 2635 2977 2637 2979
rect 2640 2977 2642 2979
rect 2645 2977 2647 2979
rect 2650 2977 2652 2979
rect 2655 2977 2657 2979
rect 2660 2977 2662 2979
rect 2665 2977 2667 2979
rect 2670 2977 2672 2979
rect 2675 2977 2677 2979
rect 2680 2977 2682 2979
rect 2685 2977 2687 2979
rect 2690 2977 2692 2979
rect 2695 2977 2697 2979
rect 2700 2977 2702 2979
rect 2705 2977 2707 2979
rect 2710 2977 2712 2979
rect 2715 2977 2717 2979
rect 2720 2977 2722 2979
rect 2725 2977 2727 2979
rect 2730 2977 2732 2979
rect 2735 2977 2737 2979
rect 2740 2977 2742 2979
rect 2745 2977 2747 2979
rect 2750 2977 2752 2979
rect 2755 2977 2757 2979
rect 2760 2977 2762 2979
rect 2765 2977 2767 2979
rect 2770 2977 2772 2979
rect 2775 2977 2777 2979
rect 2780 2977 2782 2979
rect 2785 2977 2787 2979
rect 2790 2977 2792 2979
rect 2795 2977 2797 2979
rect 2800 2977 2802 2979
rect 2805 2977 2807 2979
rect 2810 2977 2812 2979
rect 2815 2977 2817 2979
rect 2820 2977 2822 2979
rect 2825 2977 2827 2979
rect 2830 2977 2832 2979
rect 2835 2977 2837 2979
rect 2840 2977 2842 2979
rect 2845 2977 2847 2979
rect 2850 2977 2852 2979
rect 2855 2977 2857 2979
rect 2860 2977 2862 2979
rect 2865 2977 2867 2979
rect 2870 2977 2872 2979
rect 2875 2977 2877 2979
rect 2880 2977 2882 2979
rect 2885 2977 2887 2979
rect -620 2973 -618 2975
rect -615 2973 -613 2975
rect -610 2973 -608 2975
rect -605 2973 -603 2975
rect -600 2973 -598 2975
rect -595 2973 -593 2975
rect -590 2973 -588 2975
rect -585 2973 -583 2975
rect -580 2973 -578 2975
rect -575 2973 -573 2975
rect -570 2973 -568 2975
rect -565 2973 -563 2975
rect -560 2973 -558 2975
rect -555 2973 -553 2975
rect -550 2973 -548 2975
rect -545 2973 -543 2975
rect -540 2973 -538 2975
rect -535 2973 -533 2975
rect -530 2973 -528 2975
rect -525 2973 -523 2975
rect -520 2973 -518 2975
rect -515 2973 -513 2975
rect -510 2973 -508 2975
rect -505 2973 -503 2975
rect -500 2973 -498 2975
rect -495 2973 -493 2975
rect -490 2973 -488 2975
rect -485 2973 -483 2975
rect -480 2973 -478 2975
rect -475 2973 -473 2975
rect -470 2973 -468 2975
rect -465 2973 -463 2975
rect -460 2973 -458 2975
rect -455 2973 -453 2975
rect -450 2973 -448 2975
rect -445 2973 -443 2975
rect -440 2973 -438 2975
rect -435 2973 -433 2975
rect -430 2973 -428 2975
rect -425 2973 -423 2975
rect -420 2973 -418 2975
rect -415 2973 -413 2975
rect -410 2973 -408 2975
rect -405 2973 -403 2975
rect -400 2973 -398 2975
rect -395 2973 -393 2975
rect -390 2973 -388 2975
rect -385 2973 -383 2975
rect -380 2973 -378 2975
rect -375 2973 -373 2975
rect 622 2972 624 2974
rect 638 2973 640 2975
rect 654 2973 656 2975
rect 678 2973 680 2975
rect 694 2973 696 2975
rect 710 2973 712 2975
rect 726 2973 728 2975
rect 2620 2972 2622 2974
rect 2625 2972 2627 2974
rect 2630 2972 2632 2974
rect 2635 2972 2637 2974
rect 2640 2972 2642 2974
rect 2645 2972 2647 2974
rect 2650 2972 2652 2974
rect 2655 2972 2657 2974
rect 2660 2972 2662 2974
rect 2665 2972 2667 2974
rect 2670 2972 2672 2974
rect 2675 2972 2677 2974
rect 2680 2972 2682 2974
rect 2685 2972 2687 2974
rect 2690 2972 2692 2974
rect 2695 2972 2697 2974
rect 2700 2972 2702 2974
rect 2705 2972 2707 2974
rect 2710 2972 2712 2974
rect 2715 2972 2717 2974
rect 2720 2972 2722 2974
rect 2725 2972 2727 2974
rect 2730 2972 2732 2974
rect 2735 2972 2737 2974
rect 2740 2972 2742 2974
rect 2745 2972 2747 2974
rect 2750 2972 2752 2974
rect 2755 2972 2757 2974
rect 2760 2972 2762 2974
rect 2765 2972 2767 2974
rect 2770 2972 2772 2974
rect 2775 2972 2777 2974
rect 2780 2972 2782 2974
rect 2785 2972 2787 2974
rect 2790 2972 2792 2974
rect 2795 2972 2797 2974
rect 2800 2972 2802 2974
rect 2805 2972 2807 2974
rect 2810 2972 2812 2974
rect 2815 2972 2817 2974
rect 2820 2972 2822 2974
rect 2825 2972 2827 2974
rect 2830 2972 2832 2974
rect 2835 2972 2837 2974
rect 2840 2972 2842 2974
rect 2845 2972 2847 2974
rect 2850 2972 2852 2974
rect 2855 2972 2857 2974
rect 2860 2972 2862 2974
rect 2865 2972 2867 2974
rect 2870 2972 2872 2974
rect 2875 2972 2877 2974
rect 2880 2972 2882 2974
rect 2885 2972 2887 2974
rect -620 2968 -618 2970
rect -615 2968 -613 2970
rect -610 2968 -608 2970
rect -605 2968 -603 2970
rect -600 2968 -598 2970
rect -595 2968 -593 2970
rect -590 2968 -588 2970
rect -585 2968 -583 2970
rect -580 2968 -578 2970
rect -575 2968 -573 2970
rect -570 2968 -568 2970
rect -565 2968 -563 2970
rect -560 2968 -558 2970
rect -555 2968 -553 2970
rect -550 2968 -548 2970
rect -545 2968 -543 2970
rect -540 2968 -538 2970
rect -535 2968 -533 2970
rect -530 2968 -528 2970
rect -525 2968 -523 2970
rect -520 2968 -518 2970
rect -515 2968 -513 2970
rect -510 2968 -508 2970
rect -505 2968 -503 2970
rect -500 2968 -498 2970
rect -495 2968 -493 2970
rect -490 2968 -488 2970
rect -485 2968 -483 2970
rect -480 2968 -478 2970
rect -475 2968 -473 2970
rect -470 2968 -468 2970
rect -465 2968 -463 2970
rect -460 2968 -458 2970
rect -455 2968 -453 2970
rect -450 2968 -448 2970
rect -445 2968 -443 2970
rect -440 2968 -438 2970
rect -435 2968 -433 2970
rect -430 2968 -428 2970
rect -425 2968 -423 2970
rect -420 2968 -418 2970
rect -415 2968 -413 2970
rect -410 2968 -408 2970
rect -405 2968 -403 2970
rect -400 2968 -398 2970
rect -395 2968 -393 2970
rect -390 2968 -388 2970
rect -385 2968 -383 2970
rect -380 2968 -378 2970
rect -375 2968 -373 2970
rect 622 2967 624 2969
rect 638 2968 640 2970
rect 654 2968 656 2970
rect 678 2968 680 2970
rect 694 2968 696 2970
rect 710 2968 712 2970
rect 726 2968 728 2970
rect 2620 2967 2622 2969
rect 2625 2967 2627 2969
rect 2630 2967 2632 2969
rect 2635 2967 2637 2969
rect 2640 2967 2642 2969
rect 2645 2967 2647 2969
rect 2650 2967 2652 2969
rect 2655 2967 2657 2969
rect 2660 2967 2662 2969
rect 2665 2967 2667 2969
rect 2670 2967 2672 2969
rect 2675 2967 2677 2969
rect 2680 2967 2682 2969
rect 2685 2967 2687 2969
rect 2690 2967 2692 2969
rect 2695 2967 2697 2969
rect 2700 2967 2702 2969
rect 2705 2967 2707 2969
rect 2710 2967 2712 2969
rect 2715 2967 2717 2969
rect 2720 2967 2722 2969
rect 2725 2967 2727 2969
rect 2730 2967 2732 2969
rect 2735 2967 2737 2969
rect 2740 2967 2742 2969
rect 2745 2967 2747 2969
rect 2750 2967 2752 2969
rect 2755 2967 2757 2969
rect 2760 2967 2762 2969
rect 2765 2967 2767 2969
rect 2770 2967 2772 2969
rect 2775 2967 2777 2969
rect 2780 2967 2782 2969
rect 2785 2967 2787 2969
rect 2790 2967 2792 2969
rect 2795 2967 2797 2969
rect 2800 2967 2802 2969
rect 2805 2967 2807 2969
rect 2810 2967 2812 2969
rect 2815 2967 2817 2969
rect 2820 2967 2822 2969
rect 2825 2967 2827 2969
rect 2830 2967 2832 2969
rect 2835 2967 2837 2969
rect 2840 2967 2842 2969
rect 2845 2967 2847 2969
rect 2850 2967 2852 2969
rect 2855 2967 2857 2969
rect 2860 2967 2862 2969
rect 2865 2967 2867 2969
rect 2870 2967 2872 2969
rect 2875 2967 2877 2969
rect 2880 2967 2882 2969
rect 2885 2967 2887 2969
rect -620 2963 -618 2965
rect -615 2963 -613 2965
rect -610 2963 -608 2965
rect -605 2963 -603 2965
rect -600 2963 -598 2965
rect -595 2963 -593 2965
rect -590 2963 -588 2965
rect -585 2963 -583 2965
rect -580 2963 -578 2965
rect -575 2963 -573 2965
rect -570 2963 -568 2965
rect -565 2963 -563 2965
rect -560 2963 -558 2965
rect -555 2963 -553 2965
rect -550 2963 -548 2965
rect -545 2963 -543 2965
rect -540 2963 -538 2965
rect -535 2963 -533 2965
rect -530 2963 -528 2965
rect -525 2963 -523 2965
rect -520 2963 -518 2965
rect -515 2963 -513 2965
rect -510 2963 -508 2965
rect -505 2963 -503 2965
rect -500 2963 -498 2965
rect -495 2963 -493 2965
rect -490 2963 -488 2965
rect -485 2963 -483 2965
rect -480 2963 -478 2965
rect -475 2963 -473 2965
rect -470 2963 -468 2965
rect -465 2963 -463 2965
rect -460 2963 -458 2965
rect -455 2963 -453 2965
rect -450 2963 -448 2965
rect -445 2963 -443 2965
rect -440 2963 -438 2965
rect -435 2963 -433 2965
rect -430 2963 -428 2965
rect -425 2963 -423 2965
rect -420 2963 -418 2965
rect -415 2963 -413 2965
rect -410 2963 -408 2965
rect -405 2963 -403 2965
rect -400 2963 -398 2965
rect -395 2963 -393 2965
rect -390 2963 -388 2965
rect -385 2963 -383 2965
rect -380 2963 -378 2965
rect -375 2963 -373 2965
rect 622 2962 624 2964
rect 638 2963 640 2965
rect 654 2963 656 2965
rect 678 2963 680 2965
rect 694 2963 696 2965
rect 710 2963 712 2965
rect 726 2963 728 2965
rect 2620 2962 2622 2964
rect 2625 2962 2627 2964
rect 2630 2962 2632 2964
rect 2635 2962 2637 2964
rect 2640 2962 2642 2964
rect 2645 2962 2647 2964
rect 2650 2962 2652 2964
rect 2655 2962 2657 2964
rect 2660 2962 2662 2964
rect 2665 2962 2667 2964
rect 2670 2962 2672 2964
rect 2675 2962 2677 2964
rect 2680 2962 2682 2964
rect 2685 2962 2687 2964
rect 2690 2962 2692 2964
rect 2695 2962 2697 2964
rect 2700 2962 2702 2964
rect 2705 2962 2707 2964
rect 2710 2962 2712 2964
rect 2715 2962 2717 2964
rect 2720 2962 2722 2964
rect 2725 2962 2727 2964
rect 2730 2962 2732 2964
rect 2735 2962 2737 2964
rect 2740 2962 2742 2964
rect 2745 2962 2747 2964
rect 2750 2962 2752 2964
rect 2755 2962 2757 2964
rect 2760 2962 2762 2964
rect 2765 2962 2767 2964
rect 2770 2962 2772 2964
rect 2775 2962 2777 2964
rect 2780 2962 2782 2964
rect 2785 2962 2787 2964
rect 2790 2962 2792 2964
rect 2795 2962 2797 2964
rect 2800 2962 2802 2964
rect 2805 2962 2807 2964
rect 2810 2962 2812 2964
rect 2815 2962 2817 2964
rect 2820 2962 2822 2964
rect 2825 2962 2827 2964
rect 2830 2962 2832 2964
rect 2835 2962 2837 2964
rect 2840 2962 2842 2964
rect 2845 2962 2847 2964
rect 2850 2962 2852 2964
rect 2855 2962 2857 2964
rect 2860 2962 2862 2964
rect 2865 2962 2867 2964
rect 2870 2962 2872 2964
rect 2875 2962 2877 2964
rect 2880 2962 2882 2964
rect 2885 2962 2887 2964
rect -620 2958 -618 2960
rect -615 2958 -613 2960
rect -610 2958 -608 2960
rect -605 2958 -603 2960
rect -600 2958 -598 2960
rect -595 2958 -593 2960
rect -590 2958 -588 2960
rect -585 2958 -583 2960
rect -580 2958 -578 2960
rect -575 2958 -573 2960
rect -570 2958 -568 2960
rect -565 2958 -563 2960
rect -560 2958 -558 2960
rect -555 2958 -553 2960
rect -550 2958 -548 2960
rect -545 2958 -543 2960
rect -540 2958 -538 2960
rect -535 2958 -533 2960
rect -530 2958 -528 2960
rect -525 2958 -523 2960
rect -520 2958 -518 2960
rect -515 2958 -513 2960
rect -510 2958 -508 2960
rect -505 2958 -503 2960
rect -500 2958 -498 2960
rect -495 2958 -493 2960
rect -490 2958 -488 2960
rect -485 2958 -483 2960
rect -480 2958 -478 2960
rect -475 2958 -473 2960
rect -470 2958 -468 2960
rect -465 2958 -463 2960
rect -460 2958 -458 2960
rect -455 2958 -453 2960
rect -450 2958 -448 2960
rect -445 2958 -443 2960
rect -440 2958 -438 2960
rect -435 2958 -433 2960
rect -430 2958 -428 2960
rect -425 2958 -423 2960
rect -420 2958 -418 2960
rect -415 2958 -413 2960
rect -410 2958 -408 2960
rect -405 2958 -403 2960
rect -400 2958 -398 2960
rect -395 2958 -393 2960
rect -390 2958 -388 2960
rect -385 2958 -383 2960
rect -380 2958 -378 2960
rect -375 2958 -373 2960
rect 622 2957 624 2959
rect 638 2958 640 2960
rect 654 2958 656 2960
rect 678 2958 680 2960
rect 694 2958 696 2960
rect 710 2958 712 2960
rect 726 2958 728 2960
rect 2620 2957 2622 2959
rect 2625 2957 2627 2959
rect 2630 2957 2632 2959
rect 2635 2957 2637 2959
rect 2640 2957 2642 2959
rect 2645 2957 2647 2959
rect 2650 2957 2652 2959
rect 2655 2957 2657 2959
rect 2660 2957 2662 2959
rect 2665 2957 2667 2959
rect 2670 2957 2672 2959
rect 2675 2957 2677 2959
rect 2680 2957 2682 2959
rect 2685 2957 2687 2959
rect 2690 2957 2692 2959
rect 2695 2957 2697 2959
rect 2700 2957 2702 2959
rect 2705 2957 2707 2959
rect 2710 2957 2712 2959
rect 2715 2957 2717 2959
rect 2720 2957 2722 2959
rect 2725 2957 2727 2959
rect 2730 2957 2732 2959
rect 2735 2957 2737 2959
rect 2740 2957 2742 2959
rect 2745 2957 2747 2959
rect 2750 2957 2752 2959
rect 2755 2957 2757 2959
rect 2760 2957 2762 2959
rect 2765 2957 2767 2959
rect 2770 2957 2772 2959
rect 2775 2957 2777 2959
rect 2780 2957 2782 2959
rect 2785 2957 2787 2959
rect 2790 2957 2792 2959
rect 2795 2957 2797 2959
rect 2800 2957 2802 2959
rect 2805 2957 2807 2959
rect 2810 2957 2812 2959
rect 2815 2957 2817 2959
rect 2820 2957 2822 2959
rect 2825 2957 2827 2959
rect 2830 2957 2832 2959
rect 2835 2957 2837 2959
rect 2840 2957 2842 2959
rect 2845 2957 2847 2959
rect 2850 2957 2852 2959
rect 2855 2957 2857 2959
rect 2860 2957 2862 2959
rect 2865 2957 2867 2959
rect 2870 2957 2872 2959
rect 2875 2957 2877 2959
rect 2880 2957 2882 2959
rect 2885 2957 2887 2959
rect -620 2953 -618 2955
rect -615 2953 -613 2955
rect -610 2953 -608 2955
rect -605 2953 -603 2955
rect -600 2953 -598 2955
rect -595 2953 -593 2955
rect -590 2953 -588 2955
rect -585 2953 -583 2955
rect -580 2953 -578 2955
rect -575 2953 -573 2955
rect -570 2953 -568 2955
rect -565 2953 -563 2955
rect -560 2953 -558 2955
rect -555 2953 -553 2955
rect -550 2953 -548 2955
rect -545 2953 -543 2955
rect -540 2953 -538 2955
rect -535 2953 -533 2955
rect -530 2953 -528 2955
rect -525 2953 -523 2955
rect -520 2953 -518 2955
rect -515 2953 -513 2955
rect -510 2953 -508 2955
rect -505 2953 -503 2955
rect -500 2953 -498 2955
rect -495 2953 -493 2955
rect -490 2953 -488 2955
rect -485 2953 -483 2955
rect -480 2953 -478 2955
rect -475 2953 -473 2955
rect -470 2953 -468 2955
rect -465 2953 -463 2955
rect -460 2953 -458 2955
rect -455 2953 -453 2955
rect -450 2953 -448 2955
rect -445 2953 -443 2955
rect -440 2953 -438 2955
rect -435 2953 -433 2955
rect -430 2953 -428 2955
rect -425 2953 -423 2955
rect -420 2953 -418 2955
rect -415 2953 -413 2955
rect -410 2953 -408 2955
rect -405 2953 -403 2955
rect -400 2953 -398 2955
rect -395 2953 -393 2955
rect -390 2953 -388 2955
rect -385 2953 -383 2955
rect -380 2953 -378 2955
rect -375 2953 -373 2955
rect 622 2952 624 2954
rect 638 2953 640 2955
rect 654 2953 656 2955
rect 678 2953 680 2955
rect 694 2953 696 2955
rect 710 2953 712 2955
rect 726 2953 728 2955
rect 2620 2952 2622 2954
rect 2625 2952 2627 2954
rect 2630 2952 2632 2954
rect 2635 2952 2637 2954
rect 2640 2952 2642 2954
rect 2645 2952 2647 2954
rect 2650 2952 2652 2954
rect 2655 2952 2657 2954
rect 2660 2952 2662 2954
rect 2665 2952 2667 2954
rect 2670 2952 2672 2954
rect 2675 2952 2677 2954
rect 2680 2952 2682 2954
rect 2685 2952 2687 2954
rect 2690 2952 2692 2954
rect 2695 2952 2697 2954
rect 2700 2952 2702 2954
rect 2705 2952 2707 2954
rect 2710 2952 2712 2954
rect 2715 2952 2717 2954
rect 2720 2952 2722 2954
rect 2725 2952 2727 2954
rect 2730 2952 2732 2954
rect 2735 2952 2737 2954
rect 2740 2952 2742 2954
rect 2745 2952 2747 2954
rect 2750 2952 2752 2954
rect 2755 2952 2757 2954
rect 2760 2952 2762 2954
rect 2765 2952 2767 2954
rect 2770 2952 2772 2954
rect 2775 2952 2777 2954
rect 2780 2952 2782 2954
rect 2785 2952 2787 2954
rect 2790 2952 2792 2954
rect 2795 2952 2797 2954
rect 2800 2952 2802 2954
rect 2805 2952 2807 2954
rect 2810 2952 2812 2954
rect 2815 2952 2817 2954
rect 2820 2952 2822 2954
rect 2825 2952 2827 2954
rect 2830 2952 2832 2954
rect 2835 2952 2837 2954
rect 2840 2952 2842 2954
rect 2845 2952 2847 2954
rect 2850 2952 2852 2954
rect 2855 2952 2857 2954
rect 2860 2952 2862 2954
rect 2865 2952 2867 2954
rect 2870 2952 2872 2954
rect 2875 2952 2877 2954
rect 2880 2952 2882 2954
rect 2885 2952 2887 2954
rect -620 2948 -618 2950
rect -615 2948 -613 2950
rect -610 2948 -608 2950
rect -605 2948 -603 2950
rect -600 2948 -598 2950
rect -595 2948 -593 2950
rect -590 2948 -588 2950
rect -585 2948 -583 2950
rect -580 2948 -578 2950
rect -575 2948 -573 2950
rect -570 2948 -568 2950
rect -565 2948 -563 2950
rect -560 2948 -558 2950
rect -555 2948 -553 2950
rect -550 2948 -548 2950
rect -545 2948 -543 2950
rect -540 2948 -538 2950
rect -535 2948 -533 2950
rect -530 2948 -528 2950
rect -525 2948 -523 2950
rect -520 2948 -518 2950
rect -515 2948 -513 2950
rect -510 2948 -508 2950
rect -505 2948 -503 2950
rect -500 2948 -498 2950
rect -495 2948 -493 2950
rect -490 2948 -488 2950
rect -485 2948 -483 2950
rect -480 2948 -478 2950
rect -475 2948 -473 2950
rect -470 2948 -468 2950
rect -465 2948 -463 2950
rect -460 2948 -458 2950
rect -455 2948 -453 2950
rect -450 2948 -448 2950
rect -445 2948 -443 2950
rect -440 2948 -438 2950
rect -435 2948 -433 2950
rect -430 2948 -428 2950
rect -425 2948 -423 2950
rect -420 2948 -418 2950
rect -415 2948 -413 2950
rect -410 2948 -408 2950
rect -405 2948 -403 2950
rect -400 2948 -398 2950
rect -395 2948 -393 2950
rect -390 2948 -388 2950
rect -385 2948 -383 2950
rect -380 2948 -378 2950
rect -375 2948 -373 2950
rect 622 2947 624 2949
rect 638 2948 640 2950
rect 654 2948 656 2950
rect 678 2948 680 2950
rect 694 2948 696 2950
rect 710 2948 712 2950
rect 726 2948 728 2950
rect 2620 2947 2622 2949
rect 2625 2947 2627 2949
rect 2630 2947 2632 2949
rect 2635 2947 2637 2949
rect 2640 2947 2642 2949
rect 2645 2947 2647 2949
rect 2650 2947 2652 2949
rect 2655 2947 2657 2949
rect 2660 2947 2662 2949
rect 2665 2947 2667 2949
rect 2670 2947 2672 2949
rect 2675 2947 2677 2949
rect 2680 2947 2682 2949
rect 2685 2947 2687 2949
rect 2690 2947 2692 2949
rect 2695 2947 2697 2949
rect 2700 2947 2702 2949
rect 2705 2947 2707 2949
rect 2710 2947 2712 2949
rect 2715 2947 2717 2949
rect 2720 2947 2722 2949
rect 2725 2947 2727 2949
rect 2730 2947 2732 2949
rect 2735 2947 2737 2949
rect 2740 2947 2742 2949
rect 2745 2947 2747 2949
rect 2750 2947 2752 2949
rect 2755 2947 2757 2949
rect 2760 2947 2762 2949
rect 2765 2947 2767 2949
rect 2770 2947 2772 2949
rect 2775 2947 2777 2949
rect 2780 2947 2782 2949
rect 2785 2947 2787 2949
rect 2790 2947 2792 2949
rect 2795 2947 2797 2949
rect 2800 2947 2802 2949
rect 2805 2947 2807 2949
rect 2810 2947 2812 2949
rect 2815 2947 2817 2949
rect 2820 2947 2822 2949
rect 2825 2947 2827 2949
rect 2830 2947 2832 2949
rect 2835 2947 2837 2949
rect 2840 2947 2842 2949
rect 2845 2947 2847 2949
rect 2850 2947 2852 2949
rect 2855 2947 2857 2949
rect 2860 2947 2862 2949
rect 2865 2947 2867 2949
rect 2870 2947 2872 2949
rect 2875 2947 2877 2949
rect 2880 2947 2882 2949
rect 2885 2947 2887 2949
rect -620 2943 -618 2945
rect -615 2943 -613 2945
rect -610 2943 -608 2945
rect -605 2943 -603 2945
rect -600 2943 -598 2945
rect -595 2943 -593 2945
rect -590 2943 -588 2945
rect -585 2943 -583 2945
rect -580 2943 -578 2945
rect -575 2943 -573 2945
rect -570 2943 -568 2945
rect -565 2943 -563 2945
rect -560 2943 -558 2945
rect -555 2943 -553 2945
rect -550 2943 -548 2945
rect -545 2943 -543 2945
rect -540 2943 -538 2945
rect -535 2943 -533 2945
rect -530 2943 -528 2945
rect -525 2943 -523 2945
rect -520 2943 -518 2945
rect -515 2943 -513 2945
rect -510 2943 -508 2945
rect -505 2943 -503 2945
rect -500 2943 -498 2945
rect -495 2943 -493 2945
rect -490 2943 -488 2945
rect -485 2943 -483 2945
rect -480 2943 -478 2945
rect -475 2943 -473 2945
rect -470 2943 -468 2945
rect -465 2943 -463 2945
rect -460 2943 -458 2945
rect -455 2943 -453 2945
rect -450 2943 -448 2945
rect -445 2943 -443 2945
rect -440 2943 -438 2945
rect -435 2943 -433 2945
rect -430 2943 -428 2945
rect -425 2943 -423 2945
rect -420 2943 -418 2945
rect -415 2943 -413 2945
rect -410 2943 -408 2945
rect -405 2943 -403 2945
rect -400 2943 -398 2945
rect -395 2943 -393 2945
rect -390 2943 -388 2945
rect -385 2943 -383 2945
rect -380 2943 -378 2945
rect -375 2943 -373 2945
rect 622 2942 624 2944
rect 638 2943 640 2945
rect 654 2943 656 2945
rect 678 2943 680 2945
rect 694 2943 696 2945
rect 710 2943 712 2945
rect 726 2943 728 2945
rect 2620 2942 2622 2944
rect 2625 2942 2627 2944
rect 2630 2942 2632 2944
rect 2635 2942 2637 2944
rect 2640 2942 2642 2944
rect 2645 2942 2647 2944
rect 2650 2942 2652 2944
rect 2655 2942 2657 2944
rect 2660 2942 2662 2944
rect 2665 2942 2667 2944
rect 2670 2942 2672 2944
rect 2675 2942 2677 2944
rect 2680 2942 2682 2944
rect 2685 2942 2687 2944
rect 2690 2942 2692 2944
rect 2695 2942 2697 2944
rect 2700 2942 2702 2944
rect 2705 2942 2707 2944
rect 2710 2942 2712 2944
rect 2715 2942 2717 2944
rect 2720 2942 2722 2944
rect 2725 2942 2727 2944
rect 2730 2942 2732 2944
rect 2735 2942 2737 2944
rect 2740 2942 2742 2944
rect 2745 2942 2747 2944
rect 2750 2942 2752 2944
rect 2755 2942 2757 2944
rect 2760 2942 2762 2944
rect 2765 2942 2767 2944
rect 2770 2942 2772 2944
rect 2775 2942 2777 2944
rect 2780 2942 2782 2944
rect 2785 2942 2787 2944
rect 2790 2942 2792 2944
rect 2795 2942 2797 2944
rect 2800 2942 2802 2944
rect 2805 2942 2807 2944
rect 2810 2942 2812 2944
rect 2815 2942 2817 2944
rect 2820 2942 2822 2944
rect 2825 2942 2827 2944
rect 2830 2942 2832 2944
rect 2835 2942 2837 2944
rect 2840 2942 2842 2944
rect 2845 2942 2847 2944
rect 2850 2942 2852 2944
rect 2855 2942 2857 2944
rect 2860 2942 2862 2944
rect 2865 2942 2867 2944
rect 2870 2942 2872 2944
rect 2875 2942 2877 2944
rect 2880 2942 2882 2944
rect 2885 2942 2887 2944
rect -620 2938 -618 2940
rect -615 2938 -613 2940
rect -610 2938 -608 2940
rect -605 2938 -603 2940
rect -600 2938 -598 2940
rect -595 2938 -593 2940
rect -590 2938 -588 2940
rect -585 2938 -583 2940
rect -580 2938 -578 2940
rect -575 2938 -573 2940
rect -570 2938 -568 2940
rect -565 2938 -563 2940
rect -560 2938 -558 2940
rect -555 2938 -553 2940
rect -550 2938 -548 2940
rect -545 2938 -543 2940
rect -540 2938 -538 2940
rect -535 2938 -533 2940
rect -530 2938 -528 2940
rect -525 2938 -523 2940
rect -520 2938 -518 2940
rect -515 2938 -513 2940
rect -510 2938 -508 2940
rect -505 2938 -503 2940
rect -500 2938 -498 2940
rect -495 2938 -493 2940
rect -490 2938 -488 2940
rect -485 2938 -483 2940
rect -480 2938 -478 2940
rect -475 2938 -473 2940
rect -470 2938 -468 2940
rect -465 2938 -463 2940
rect -460 2938 -458 2940
rect -455 2938 -453 2940
rect -450 2938 -448 2940
rect -445 2938 -443 2940
rect -440 2938 -438 2940
rect -435 2938 -433 2940
rect -430 2938 -428 2940
rect -425 2938 -423 2940
rect -420 2938 -418 2940
rect -415 2938 -413 2940
rect -410 2938 -408 2940
rect -405 2938 -403 2940
rect -400 2938 -398 2940
rect -395 2938 -393 2940
rect -390 2938 -388 2940
rect -385 2938 -383 2940
rect -380 2938 -378 2940
rect -375 2938 -373 2940
rect 622 2937 624 2939
rect 638 2938 640 2940
rect 654 2938 656 2940
rect 678 2938 680 2940
rect 694 2938 696 2940
rect 710 2938 712 2940
rect 726 2938 728 2940
rect 2620 2937 2622 2939
rect 2625 2937 2627 2939
rect 2630 2937 2632 2939
rect 2635 2937 2637 2939
rect 2640 2937 2642 2939
rect 2645 2937 2647 2939
rect 2650 2937 2652 2939
rect 2655 2937 2657 2939
rect 2660 2937 2662 2939
rect 2665 2937 2667 2939
rect 2670 2937 2672 2939
rect 2675 2937 2677 2939
rect 2680 2937 2682 2939
rect 2685 2937 2687 2939
rect 2690 2937 2692 2939
rect 2695 2937 2697 2939
rect 2700 2937 2702 2939
rect 2705 2937 2707 2939
rect 2710 2937 2712 2939
rect 2715 2937 2717 2939
rect 2720 2937 2722 2939
rect 2725 2937 2727 2939
rect 2730 2937 2732 2939
rect 2735 2937 2737 2939
rect 2740 2937 2742 2939
rect 2745 2937 2747 2939
rect 2750 2937 2752 2939
rect 2755 2937 2757 2939
rect 2760 2937 2762 2939
rect 2765 2937 2767 2939
rect 2770 2937 2772 2939
rect 2775 2937 2777 2939
rect 2780 2937 2782 2939
rect 2785 2937 2787 2939
rect 2790 2937 2792 2939
rect 2795 2937 2797 2939
rect 2800 2937 2802 2939
rect 2805 2937 2807 2939
rect 2810 2937 2812 2939
rect 2815 2937 2817 2939
rect 2820 2937 2822 2939
rect 2825 2937 2827 2939
rect 2830 2937 2832 2939
rect 2835 2937 2837 2939
rect 2840 2937 2842 2939
rect 2845 2937 2847 2939
rect 2850 2937 2852 2939
rect 2855 2937 2857 2939
rect 2860 2937 2862 2939
rect 2865 2937 2867 2939
rect 2870 2937 2872 2939
rect 2875 2937 2877 2939
rect 2880 2937 2882 2939
rect 2885 2937 2887 2939
rect -620 2933 -618 2935
rect -615 2933 -613 2935
rect -610 2933 -608 2935
rect -605 2933 -603 2935
rect -600 2933 -598 2935
rect -595 2933 -593 2935
rect -590 2933 -588 2935
rect -585 2933 -583 2935
rect -580 2933 -578 2935
rect -575 2933 -573 2935
rect -570 2933 -568 2935
rect -565 2933 -563 2935
rect -560 2933 -558 2935
rect -555 2933 -553 2935
rect -550 2933 -548 2935
rect -545 2933 -543 2935
rect -540 2933 -538 2935
rect -535 2933 -533 2935
rect -530 2933 -528 2935
rect -525 2933 -523 2935
rect -520 2933 -518 2935
rect -515 2933 -513 2935
rect -510 2933 -508 2935
rect -505 2933 -503 2935
rect -500 2933 -498 2935
rect -495 2933 -493 2935
rect -490 2933 -488 2935
rect -485 2933 -483 2935
rect -480 2933 -478 2935
rect -475 2933 -473 2935
rect -470 2933 -468 2935
rect -465 2933 -463 2935
rect -460 2933 -458 2935
rect -455 2933 -453 2935
rect -450 2933 -448 2935
rect -445 2933 -443 2935
rect -440 2933 -438 2935
rect -435 2933 -433 2935
rect -430 2933 -428 2935
rect -425 2933 -423 2935
rect -420 2933 -418 2935
rect -415 2933 -413 2935
rect -410 2933 -408 2935
rect -405 2933 -403 2935
rect -400 2933 -398 2935
rect -395 2933 -393 2935
rect -390 2933 -388 2935
rect -385 2933 -383 2935
rect -380 2933 -378 2935
rect -375 2933 -373 2935
rect 622 2932 624 2934
rect 638 2933 640 2935
rect 654 2933 656 2935
rect 678 2933 680 2935
rect 694 2933 696 2935
rect 710 2933 712 2935
rect 726 2933 728 2935
rect 2620 2932 2622 2934
rect 2625 2932 2627 2934
rect 2630 2932 2632 2934
rect 2635 2932 2637 2934
rect 2640 2932 2642 2934
rect 2645 2932 2647 2934
rect 2650 2932 2652 2934
rect 2655 2932 2657 2934
rect 2660 2932 2662 2934
rect 2665 2932 2667 2934
rect 2670 2932 2672 2934
rect 2675 2932 2677 2934
rect 2680 2932 2682 2934
rect 2685 2932 2687 2934
rect 2690 2932 2692 2934
rect 2695 2932 2697 2934
rect 2700 2932 2702 2934
rect 2705 2932 2707 2934
rect 2710 2932 2712 2934
rect 2715 2932 2717 2934
rect 2720 2932 2722 2934
rect 2725 2932 2727 2934
rect 2730 2932 2732 2934
rect 2735 2932 2737 2934
rect 2740 2932 2742 2934
rect 2745 2932 2747 2934
rect 2750 2932 2752 2934
rect 2755 2932 2757 2934
rect 2760 2932 2762 2934
rect 2765 2932 2767 2934
rect 2770 2932 2772 2934
rect 2775 2932 2777 2934
rect 2780 2932 2782 2934
rect 2785 2932 2787 2934
rect 2790 2932 2792 2934
rect 2795 2932 2797 2934
rect 2800 2932 2802 2934
rect 2805 2932 2807 2934
rect 2810 2932 2812 2934
rect 2815 2932 2817 2934
rect 2820 2932 2822 2934
rect 2825 2932 2827 2934
rect 2830 2932 2832 2934
rect 2835 2932 2837 2934
rect 2840 2932 2842 2934
rect 2845 2932 2847 2934
rect 2850 2932 2852 2934
rect 2855 2932 2857 2934
rect 2860 2932 2862 2934
rect 2865 2932 2867 2934
rect 2870 2932 2872 2934
rect 2875 2932 2877 2934
rect 2880 2932 2882 2934
rect 2885 2932 2887 2934
rect -620 2928 -618 2930
rect -615 2928 -613 2930
rect -610 2928 -608 2930
rect -605 2928 -603 2930
rect -600 2928 -598 2930
rect -595 2928 -593 2930
rect -590 2928 -588 2930
rect -585 2928 -583 2930
rect -580 2928 -578 2930
rect -575 2928 -573 2930
rect -570 2928 -568 2930
rect -565 2928 -563 2930
rect -560 2928 -558 2930
rect -555 2928 -553 2930
rect -550 2928 -548 2930
rect -545 2928 -543 2930
rect -540 2928 -538 2930
rect -535 2928 -533 2930
rect -530 2928 -528 2930
rect -525 2928 -523 2930
rect -520 2928 -518 2930
rect -515 2928 -513 2930
rect -510 2928 -508 2930
rect -505 2928 -503 2930
rect -500 2928 -498 2930
rect -495 2928 -493 2930
rect -490 2928 -488 2930
rect -485 2928 -483 2930
rect -480 2928 -478 2930
rect -475 2928 -473 2930
rect -470 2928 -468 2930
rect -465 2928 -463 2930
rect -460 2928 -458 2930
rect -455 2928 -453 2930
rect -450 2928 -448 2930
rect -445 2928 -443 2930
rect -440 2928 -438 2930
rect -435 2928 -433 2930
rect -430 2928 -428 2930
rect -425 2928 -423 2930
rect -420 2928 -418 2930
rect -415 2928 -413 2930
rect -410 2928 -408 2930
rect -405 2928 -403 2930
rect -400 2928 -398 2930
rect -395 2928 -393 2930
rect -390 2928 -388 2930
rect -385 2928 -383 2930
rect -380 2928 -378 2930
rect -375 2928 -373 2930
rect 622 2927 624 2929
rect 638 2928 640 2930
rect 654 2928 656 2930
rect 678 2928 680 2930
rect 694 2928 696 2930
rect 710 2928 712 2930
rect 726 2928 728 2930
rect 748 2927 750 2929
rect 753 2927 755 2929
rect 764 2927 766 2929
rect 769 2927 771 2929
rect 780 2927 782 2929
rect 785 2927 787 2929
rect 796 2927 798 2929
rect 801 2927 803 2929
rect 812 2927 814 2929
rect 817 2927 819 2929
rect 828 2927 830 2929
rect 833 2927 835 2929
rect 844 2927 846 2929
rect 849 2927 851 2929
rect 860 2927 862 2929
rect 865 2927 867 2929
rect 876 2927 878 2929
rect 881 2927 883 2929
rect 892 2927 894 2929
rect 897 2927 899 2929
rect 2620 2927 2622 2929
rect 2625 2927 2627 2929
rect 2630 2927 2632 2929
rect 2635 2927 2637 2929
rect 2640 2927 2642 2929
rect 2645 2927 2647 2929
rect 2650 2927 2652 2929
rect 2655 2927 2657 2929
rect 2660 2927 2662 2929
rect 2665 2927 2667 2929
rect 2670 2927 2672 2929
rect 2675 2927 2677 2929
rect 2680 2927 2682 2929
rect 2685 2927 2687 2929
rect 2690 2927 2692 2929
rect 2695 2927 2697 2929
rect 2700 2927 2702 2929
rect 2705 2927 2707 2929
rect 2710 2927 2712 2929
rect 2715 2927 2717 2929
rect 2720 2927 2722 2929
rect 2725 2927 2727 2929
rect 2730 2927 2732 2929
rect 2735 2927 2737 2929
rect 2740 2927 2742 2929
rect 2745 2927 2747 2929
rect 2750 2927 2752 2929
rect 2755 2927 2757 2929
rect 2760 2927 2762 2929
rect 2765 2927 2767 2929
rect 2770 2927 2772 2929
rect 2775 2927 2777 2929
rect 2780 2927 2782 2929
rect 2785 2927 2787 2929
rect 2790 2927 2792 2929
rect 2795 2927 2797 2929
rect 2800 2927 2802 2929
rect 2805 2927 2807 2929
rect 2810 2927 2812 2929
rect 2815 2927 2817 2929
rect 2820 2927 2822 2929
rect 2825 2927 2827 2929
rect 2830 2927 2832 2929
rect 2835 2927 2837 2929
rect 2840 2927 2842 2929
rect 2845 2927 2847 2929
rect 2850 2927 2852 2929
rect 2855 2927 2857 2929
rect 2860 2927 2862 2929
rect 2865 2927 2867 2929
rect 2870 2927 2872 2929
rect 2875 2927 2877 2929
rect 2880 2927 2882 2929
rect 2885 2927 2887 2929
rect 1462 2925 1464 2927
rect 1518 2925 1520 2927
rect 1534 2925 1536 2927
rect 1598 2925 1600 2927
rect 1726 2925 1728 2927
rect 1894 2925 1896 2927
rect 2086 2925 2088 2927
rect -620 2923 -618 2925
rect -615 2923 -613 2925
rect -610 2923 -608 2925
rect -605 2923 -603 2925
rect -600 2923 -598 2925
rect -595 2923 -593 2925
rect -590 2923 -588 2925
rect -585 2923 -583 2925
rect -580 2923 -578 2925
rect -575 2923 -573 2925
rect -570 2923 -568 2925
rect -565 2923 -563 2925
rect -560 2923 -558 2925
rect -555 2923 -553 2925
rect -550 2923 -548 2925
rect -545 2923 -543 2925
rect -540 2923 -538 2925
rect -535 2923 -533 2925
rect -530 2923 -528 2925
rect -525 2923 -523 2925
rect -520 2923 -518 2925
rect -515 2923 -513 2925
rect -510 2923 -508 2925
rect -505 2923 -503 2925
rect -500 2923 -498 2925
rect -495 2923 -493 2925
rect -490 2923 -488 2925
rect -485 2923 -483 2925
rect -480 2923 -478 2925
rect -475 2923 -473 2925
rect -470 2923 -468 2925
rect -465 2923 -463 2925
rect -460 2923 -458 2925
rect -455 2923 -453 2925
rect -450 2923 -448 2925
rect -445 2923 -443 2925
rect -440 2923 -438 2925
rect -435 2923 -433 2925
rect -430 2923 -428 2925
rect -425 2923 -423 2925
rect -420 2923 -418 2925
rect -415 2923 -413 2925
rect -410 2923 -408 2925
rect -405 2923 -403 2925
rect -400 2923 -398 2925
rect -395 2923 -393 2925
rect -390 2923 -388 2925
rect -385 2923 -383 2925
rect -380 2923 -378 2925
rect -375 2923 -373 2925
rect 622 2922 624 2924
rect 638 2923 640 2925
rect 654 2923 656 2925
rect 678 2923 680 2925
rect 694 2923 696 2925
rect 710 2923 712 2925
rect 726 2923 728 2925
rect 748 2922 750 2924
rect 753 2922 755 2924
rect 764 2922 766 2924
rect 769 2922 771 2924
rect 780 2922 782 2924
rect 785 2922 787 2924
rect 796 2922 798 2924
rect 801 2922 803 2924
rect 812 2922 814 2924
rect 817 2922 819 2924
rect 828 2922 830 2924
rect 833 2922 835 2924
rect 844 2922 846 2924
rect 849 2922 851 2924
rect 860 2922 862 2924
rect 865 2922 867 2924
rect 876 2922 878 2924
rect 881 2922 883 2924
rect 892 2922 894 2924
rect 897 2922 899 2924
rect 2620 2922 2622 2924
rect 2625 2922 2627 2924
rect 2630 2922 2632 2924
rect 2635 2922 2637 2924
rect 2640 2922 2642 2924
rect 2645 2922 2647 2924
rect 2650 2922 2652 2924
rect 2655 2922 2657 2924
rect 2660 2922 2662 2924
rect 2665 2922 2667 2924
rect 2670 2922 2672 2924
rect 2675 2922 2677 2924
rect 2680 2922 2682 2924
rect 2685 2922 2687 2924
rect 2690 2922 2692 2924
rect 2695 2922 2697 2924
rect 2700 2922 2702 2924
rect 2705 2922 2707 2924
rect 2710 2922 2712 2924
rect 2715 2922 2717 2924
rect 2720 2922 2722 2924
rect 2725 2922 2727 2924
rect 2730 2922 2732 2924
rect 2735 2922 2737 2924
rect 2740 2922 2742 2924
rect 2745 2922 2747 2924
rect 2750 2922 2752 2924
rect 2755 2922 2757 2924
rect 2760 2922 2762 2924
rect 2765 2922 2767 2924
rect 2770 2922 2772 2924
rect 2775 2922 2777 2924
rect 2780 2922 2782 2924
rect 2785 2922 2787 2924
rect 2790 2922 2792 2924
rect 2795 2922 2797 2924
rect 2800 2922 2802 2924
rect 2805 2922 2807 2924
rect 2810 2922 2812 2924
rect 2815 2922 2817 2924
rect 2820 2922 2822 2924
rect 2825 2922 2827 2924
rect 2830 2922 2832 2924
rect 2835 2922 2837 2924
rect 2840 2922 2842 2924
rect 2845 2922 2847 2924
rect 2850 2922 2852 2924
rect 2855 2922 2857 2924
rect 2860 2922 2862 2924
rect 2865 2922 2867 2924
rect 2870 2922 2872 2924
rect 2875 2922 2877 2924
rect 2880 2922 2882 2924
rect 2885 2922 2887 2924
rect -620 2918 -618 2920
rect -615 2918 -613 2920
rect -610 2918 -608 2920
rect -605 2918 -603 2920
rect -600 2918 -598 2920
rect -595 2918 -593 2920
rect -590 2918 -588 2920
rect -585 2918 -583 2920
rect -580 2918 -578 2920
rect -575 2918 -573 2920
rect -570 2918 -568 2920
rect -565 2918 -563 2920
rect -560 2918 -558 2920
rect -555 2918 -553 2920
rect -550 2918 -548 2920
rect -545 2918 -543 2920
rect -540 2918 -538 2920
rect -535 2918 -533 2920
rect -530 2918 -528 2920
rect -525 2918 -523 2920
rect -520 2918 -518 2920
rect -515 2918 -513 2920
rect -510 2918 -508 2920
rect -505 2918 -503 2920
rect -500 2918 -498 2920
rect -495 2918 -493 2920
rect -490 2918 -488 2920
rect -485 2918 -483 2920
rect -480 2918 -478 2920
rect -475 2918 -473 2920
rect -470 2918 -468 2920
rect -465 2918 -463 2920
rect -460 2918 -458 2920
rect -455 2918 -453 2920
rect -450 2918 -448 2920
rect -445 2918 -443 2920
rect -440 2918 -438 2920
rect -435 2918 -433 2920
rect -430 2918 -428 2920
rect -425 2918 -423 2920
rect -420 2918 -418 2920
rect -415 2918 -413 2920
rect -410 2918 -408 2920
rect -405 2918 -403 2920
rect -400 2918 -398 2920
rect -395 2918 -393 2920
rect -390 2918 -388 2920
rect -385 2918 -383 2920
rect -380 2918 -378 2920
rect -375 2918 -373 2920
rect 2620 2917 2622 2919
rect 2625 2917 2627 2919
rect 2630 2917 2632 2919
rect 2635 2917 2637 2919
rect 2640 2917 2642 2919
rect 2645 2917 2647 2919
rect 2650 2917 2652 2919
rect 2655 2917 2657 2919
rect 2660 2917 2662 2919
rect 2665 2917 2667 2919
rect 2670 2917 2672 2919
rect 2675 2917 2677 2919
rect 2680 2917 2682 2919
rect 2685 2917 2687 2919
rect 2690 2917 2692 2919
rect 2695 2917 2697 2919
rect 2700 2917 2702 2919
rect 2705 2917 2707 2919
rect 2710 2917 2712 2919
rect 2715 2917 2717 2919
rect 2720 2917 2722 2919
rect 2725 2917 2727 2919
rect 2730 2917 2732 2919
rect 2735 2917 2737 2919
rect 2740 2917 2742 2919
rect 2745 2917 2747 2919
rect 2750 2917 2752 2919
rect 2755 2917 2757 2919
rect 2760 2917 2762 2919
rect 2765 2917 2767 2919
rect 2770 2917 2772 2919
rect 2775 2917 2777 2919
rect 2780 2917 2782 2919
rect 2785 2917 2787 2919
rect 2790 2917 2792 2919
rect 2795 2917 2797 2919
rect 2800 2917 2802 2919
rect 2805 2917 2807 2919
rect 2810 2917 2812 2919
rect 2815 2917 2817 2919
rect 2820 2917 2822 2919
rect 2825 2917 2827 2919
rect 2830 2917 2832 2919
rect 2835 2917 2837 2919
rect 2840 2917 2842 2919
rect 2845 2917 2847 2919
rect 2850 2917 2852 2919
rect 2855 2917 2857 2919
rect 2860 2917 2862 2919
rect 2865 2917 2867 2919
rect 2870 2917 2872 2919
rect 2875 2917 2877 2919
rect 2880 2917 2882 2919
rect 2885 2917 2887 2919
rect -620 2913 -618 2915
rect -615 2913 -613 2915
rect -610 2913 -608 2915
rect -605 2913 -603 2915
rect -600 2913 -598 2915
rect -595 2913 -593 2915
rect -590 2913 -588 2915
rect -585 2913 -583 2915
rect -580 2913 -578 2915
rect -575 2913 -573 2915
rect -570 2913 -568 2915
rect -565 2913 -563 2915
rect -560 2913 -558 2915
rect -555 2913 -553 2915
rect -550 2913 -548 2915
rect -545 2913 -543 2915
rect -540 2913 -538 2915
rect -535 2913 -533 2915
rect -530 2913 -528 2915
rect -525 2913 -523 2915
rect -520 2913 -518 2915
rect -515 2913 -513 2915
rect -510 2913 -508 2915
rect -505 2913 -503 2915
rect -500 2913 -498 2915
rect -495 2913 -493 2915
rect -490 2913 -488 2915
rect -485 2913 -483 2915
rect -480 2913 -478 2915
rect -475 2913 -473 2915
rect -470 2913 -468 2915
rect -465 2913 -463 2915
rect -460 2913 -458 2915
rect -455 2913 -453 2915
rect -450 2913 -448 2915
rect -445 2913 -443 2915
rect -440 2913 -438 2915
rect -435 2913 -433 2915
rect -430 2913 -428 2915
rect -425 2913 -423 2915
rect -420 2913 -418 2915
rect -415 2913 -413 2915
rect -410 2913 -408 2915
rect -405 2913 -403 2915
rect -400 2913 -398 2915
rect -395 2913 -393 2915
rect -390 2913 -388 2915
rect -385 2913 -383 2915
rect -380 2913 -378 2915
rect -375 2913 -373 2915
rect 2620 2912 2622 2914
rect 2625 2912 2627 2914
rect 2630 2912 2632 2914
rect 2635 2912 2637 2914
rect 2640 2912 2642 2914
rect 2645 2912 2647 2914
rect 2650 2912 2652 2914
rect 2655 2912 2657 2914
rect 2660 2912 2662 2914
rect 2665 2912 2667 2914
rect 2670 2912 2672 2914
rect 2675 2912 2677 2914
rect 2680 2912 2682 2914
rect 2685 2912 2687 2914
rect 2690 2912 2692 2914
rect 2695 2912 2697 2914
rect 2700 2912 2702 2914
rect 2705 2912 2707 2914
rect 2710 2912 2712 2914
rect 2715 2912 2717 2914
rect 2720 2912 2722 2914
rect 2725 2912 2727 2914
rect 2730 2912 2732 2914
rect 2735 2912 2737 2914
rect 2740 2912 2742 2914
rect 2745 2912 2747 2914
rect 2750 2912 2752 2914
rect 2755 2912 2757 2914
rect 2760 2912 2762 2914
rect 2765 2912 2767 2914
rect 2770 2912 2772 2914
rect 2775 2912 2777 2914
rect 2780 2912 2782 2914
rect 2785 2912 2787 2914
rect 2790 2912 2792 2914
rect 2795 2912 2797 2914
rect 2800 2912 2802 2914
rect 2805 2912 2807 2914
rect 2810 2912 2812 2914
rect 2815 2912 2817 2914
rect 2820 2912 2822 2914
rect 2825 2912 2827 2914
rect 2830 2912 2832 2914
rect 2835 2912 2837 2914
rect 2840 2912 2842 2914
rect 2845 2912 2847 2914
rect 2850 2912 2852 2914
rect 2855 2912 2857 2914
rect 2860 2912 2862 2914
rect 2865 2912 2867 2914
rect 2870 2912 2872 2914
rect 2875 2912 2877 2914
rect 2880 2912 2882 2914
rect 2885 2912 2887 2914
rect 3289 2912 3291 2914
rect -620 2908 -618 2910
rect -615 2908 -613 2910
rect -610 2908 -608 2910
rect -605 2908 -603 2910
rect -600 2908 -598 2910
rect -595 2908 -593 2910
rect -590 2908 -588 2910
rect -585 2908 -583 2910
rect -580 2908 -578 2910
rect -575 2908 -573 2910
rect -570 2908 -568 2910
rect -565 2908 -563 2910
rect -560 2908 -558 2910
rect -555 2908 -553 2910
rect -550 2908 -548 2910
rect -545 2908 -543 2910
rect -540 2908 -538 2910
rect -535 2908 -533 2910
rect -530 2908 -528 2910
rect -525 2908 -523 2910
rect -520 2908 -518 2910
rect -515 2908 -513 2910
rect -510 2908 -508 2910
rect -505 2908 -503 2910
rect -500 2908 -498 2910
rect -495 2908 -493 2910
rect -490 2908 -488 2910
rect -485 2908 -483 2910
rect -480 2908 -478 2910
rect -475 2908 -473 2910
rect -470 2908 -468 2910
rect -465 2908 -463 2910
rect -460 2908 -458 2910
rect -455 2908 -453 2910
rect -450 2908 -448 2910
rect -445 2908 -443 2910
rect -440 2908 -438 2910
rect -435 2908 -433 2910
rect -430 2908 -428 2910
rect -425 2908 -423 2910
rect -420 2908 -418 2910
rect -415 2908 -413 2910
rect -410 2908 -408 2910
rect -405 2908 -403 2910
rect -400 2908 -398 2910
rect -395 2908 -393 2910
rect -390 2908 -388 2910
rect -385 2908 -383 2910
rect -380 2908 -378 2910
rect -375 2908 -373 2910
rect 2620 2907 2622 2909
rect 2625 2907 2627 2909
rect 2630 2907 2632 2909
rect 2635 2907 2637 2909
rect 2640 2907 2642 2909
rect 2645 2907 2647 2909
rect 2650 2907 2652 2909
rect 2655 2907 2657 2909
rect 2660 2907 2662 2909
rect 2665 2907 2667 2909
rect 2670 2907 2672 2909
rect 2675 2907 2677 2909
rect 2680 2907 2682 2909
rect 2685 2907 2687 2909
rect 2690 2907 2692 2909
rect 2695 2907 2697 2909
rect 2700 2907 2702 2909
rect 2705 2907 2707 2909
rect 2710 2907 2712 2909
rect 2715 2907 2717 2909
rect 2720 2907 2722 2909
rect 2725 2907 2727 2909
rect 2730 2907 2732 2909
rect 2735 2907 2737 2909
rect 2740 2907 2742 2909
rect 2745 2907 2747 2909
rect 2750 2907 2752 2909
rect 2755 2907 2757 2909
rect 2760 2907 2762 2909
rect 2765 2907 2767 2909
rect 2770 2907 2772 2909
rect 2775 2907 2777 2909
rect 2780 2907 2782 2909
rect 2785 2907 2787 2909
rect 2790 2907 2792 2909
rect 2795 2907 2797 2909
rect 2800 2907 2802 2909
rect 2805 2907 2807 2909
rect 2810 2907 2812 2909
rect 2815 2907 2817 2909
rect 2820 2907 2822 2909
rect 2825 2907 2827 2909
rect 2830 2907 2832 2909
rect 2835 2907 2837 2909
rect 2840 2907 2842 2909
rect 2845 2907 2847 2909
rect 2850 2907 2852 2909
rect 2855 2907 2857 2909
rect 2860 2907 2862 2909
rect 2865 2907 2867 2909
rect 2870 2907 2872 2909
rect 2875 2907 2877 2909
rect 2880 2907 2882 2909
rect 2885 2907 2887 2909
rect -620 2903 -618 2905
rect -615 2903 -613 2905
rect -610 2903 -608 2905
rect -605 2903 -603 2905
rect -600 2903 -598 2905
rect -595 2903 -593 2905
rect -590 2903 -588 2905
rect -585 2903 -583 2905
rect -580 2903 -578 2905
rect -575 2903 -573 2905
rect -570 2903 -568 2905
rect -565 2903 -563 2905
rect -560 2903 -558 2905
rect -555 2903 -553 2905
rect -550 2903 -548 2905
rect -545 2903 -543 2905
rect -540 2903 -538 2905
rect -535 2903 -533 2905
rect -530 2903 -528 2905
rect -525 2903 -523 2905
rect -520 2903 -518 2905
rect -515 2903 -513 2905
rect -510 2903 -508 2905
rect -505 2903 -503 2905
rect -500 2903 -498 2905
rect -495 2903 -493 2905
rect -490 2903 -488 2905
rect -485 2903 -483 2905
rect -480 2903 -478 2905
rect -475 2903 -473 2905
rect -470 2903 -468 2905
rect -465 2903 -463 2905
rect -460 2903 -458 2905
rect -455 2903 -453 2905
rect -450 2903 -448 2905
rect -445 2903 -443 2905
rect -440 2903 -438 2905
rect -435 2903 -433 2905
rect -430 2903 -428 2905
rect -425 2903 -423 2905
rect -420 2903 -418 2905
rect -415 2903 -413 2905
rect -410 2903 -408 2905
rect -405 2903 -403 2905
rect -400 2903 -398 2905
rect -395 2903 -393 2905
rect -390 2903 -388 2905
rect -385 2903 -383 2905
rect -380 2903 -378 2905
rect -375 2903 -373 2905
rect 2620 2902 2622 2904
rect 2625 2902 2627 2904
rect 2630 2902 2632 2904
rect 2635 2902 2637 2904
rect 2640 2902 2642 2904
rect 2645 2902 2647 2904
rect 2650 2902 2652 2904
rect 2655 2902 2657 2904
rect 2660 2902 2662 2904
rect 2665 2902 2667 2904
rect 2670 2902 2672 2904
rect 2675 2902 2677 2904
rect 2680 2902 2682 2904
rect 2685 2902 2687 2904
rect 2690 2902 2692 2904
rect 2695 2902 2697 2904
rect 2700 2902 2702 2904
rect 2705 2902 2707 2904
rect 2710 2902 2712 2904
rect 2715 2902 2717 2904
rect 2720 2902 2722 2904
rect 2725 2902 2727 2904
rect 2730 2902 2732 2904
rect 2735 2902 2737 2904
rect 2740 2902 2742 2904
rect 2745 2902 2747 2904
rect 2750 2902 2752 2904
rect 2755 2902 2757 2904
rect 2760 2902 2762 2904
rect 2765 2902 2767 2904
rect 2770 2902 2772 2904
rect 2775 2902 2777 2904
rect 2780 2902 2782 2904
rect 2785 2902 2787 2904
rect 2790 2902 2792 2904
rect 2795 2902 2797 2904
rect 2800 2902 2802 2904
rect 2805 2902 2807 2904
rect 2810 2902 2812 2904
rect 2815 2902 2817 2904
rect 2820 2902 2822 2904
rect 2825 2902 2827 2904
rect 2830 2902 2832 2904
rect 2835 2902 2837 2904
rect 2840 2902 2842 2904
rect 2845 2902 2847 2904
rect 2850 2902 2852 2904
rect 2855 2902 2857 2904
rect 2860 2902 2862 2904
rect 2865 2902 2867 2904
rect 2870 2902 2872 2904
rect 2875 2902 2877 2904
rect 2880 2902 2882 2904
rect 2885 2902 2887 2904
rect -620 2898 -618 2900
rect -615 2898 -613 2900
rect -610 2898 -608 2900
rect -605 2898 -603 2900
rect -600 2898 -598 2900
rect -595 2898 -593 2900
rect -590 2898 -588 2900
rect -585 2898 -583 2900
rect -580 2898 -578 2900
rect -575 2898 -573 2900
rect -570 2898 -568 2900
rect -565 2898 -563 2900
rect -560 2898 -558 2900
rect -555 2898 -553 2900
rect -550 2898 -548 2900
rect -545 2898 -543 2900
rect -540 2898 -538 2900
rect -535 2898 -533 2900
rect -530 2898 -528 2900
rect -525 2898 -523 2900
rect -520 2898 -518 2900
rect -515 2898 -513 2900
rect -510 2898 -508 2900
rect -505 2898 -503 2900
rect -500 2898 -498 2900
rect -495 2898 -493 2900
rect -490 2898 -488 2900
rect -485 2898 -483 2900
rect -480 2898 -478 2900
rect -475 2898 -473 2900
rect -470 2898 -468 2900
rect -465 2898 -463 2900
rect -460 2898 -458 2900
rect -455 2898 -453 2900
rect -450 2898 -448 2900
rect -445 2898 -443 2900
rect -440 2898 -438 2900
rect -435 2898 -433 2900
rect -430 2898 -428 2900
rect -425 2898 -423 2900
rect -420 2898 -418 2900
rect -415 2898 -413 2900
rect -410 2898 -408 2900
rect -405 2898 -403 2900
rect -400 2898 -398 2900
rect -395 2898 -393 2900
rect -390 2898 -388 2900
rect -385 2898 -383 2900
rect -380 2898 -378 2900
rect -375 2898 -373 2900
rect 2620 2897 2622 2899
rect 2625 2897 2627 2899
rect 2630 2897 2632 2899
rect 2635 2897 2637 2899
rect 2640 2897 2642 2899
rect 2645 2897 2647 2899
rect 2650 2897 2652 2899
rect 2655 2897 2657 2899
rect 2660 2897 2662 2899
rect 2665 2897 2667 2899
rect 2670 2897 2672 2899
rect 2675 2897 2677 2899
rect 2680 2897 2682 2899
rect 2685 2897 2687 2899
rect 2690 2897 2692 2899
rect 2695 2897 2697 2899
rect 2700 2897 2702 2899
rect 2705 2897 2707 2899
rect 2710 2897 2712 2899
rect 2715 2897 2717 2899
rect 2720 2897 2722 2899
rect 2725 2897 2727 2899
rect 2730 2897 2732 2899
rect 2735 2897 2737 2899
rect 2740 2897 2742 2899
rect 2745 2897 2747 2899
rect 2750 2897 2752 2899
rect 2755 2897 2757 2899
rect 2760 2897 2762 2899
rect 2765 2897 2767 2899
rect 2770 2897 2772 2899
rect 2775 2897 2777 2899
rect 2780 2897 2782 2899
rect 2785 2897 2787 2899
rect 2790 2897 2792 2899
rect 2795 2897 2797 2899
rect 2800 2897 2802 2899
rect 2805 2897 2807 2899
rect 2810 2897 2812 2899
rect 2815 2897 2817 2899
rect 2820 2897 2822 2899
rect 2825 2897 2827 2899
rect 2830 2897 2832 2899
rect 2835 2897 2837 2899
rect 2840 2897 2842 2899
rect 2845 2897 2847 2899
rect 2850 2897 2852 2899
rect 2855 2897 2857 2899
rect 2860 2897 2862 2899
rect 2865 2897 2867 2899
rect 2870 2897 2872 2899
rect 2875 2897 2877 2899
rect 2880 2897 2882 2899
rect 2885 2897 2887 2899
rect 3289 2612 3291 2614
rect 3266 2550 3268 2552
rect 3271 2550 3273 2552
rect 3276 2550 3278 2552
rect 3281 2550 3283 2552
rect 3266 2545 3268 2547
rect 3271 2545 3273 2547
rect 3276 2545 3278 2547
rect 3281 2545 3283 2547
rect 3262 2463 3264 2465
rect 3267 2463 3269 2465
rect 3272 2463 3274 2465
rect 3277 2463 3279 2465
rect 3282 2463 3284 2465
rect 3262 2458 3264 2460
rect 3267 2458 3269 2460
rect 3272 2458 3274 2460
rect 3277 2458 3279 2460
rect 3282 2458 3284 2460
rect 3289 2312 3291 2314
rect 3267 2163 3269 2165
rect 3272 2163 3274 2165
rect 3277 2163 3279 2165
rect 3267 2158 3269 2160
rect 3272 2158 3274 2160
rect 3277 2158 3279 2160
rect 3009 2151 3011 2153
rect 3009 2121 3011 2123
rect 3009 2101 3011 2103
rect -1487 2094 -1485 2096
rect -1482 2094 -1480 2096
rect -1487 2089 -1485 2091
rect -1482 2089 -1480 2091
rect -1487 2084 -1485 2086
rect -1482 2084 -1480 2086
rect -1487 2079 -1485 2081
rect -1482 2079 -1480 2081
rect -1487 2074 -1485 2076
rect -1482 2074 -1480 2076
rect -1487 2069 -1485 2071
rect -1482 2069 -1480 2071
rect -1487 2064 -1485 2066
rect -1482 2064 -1480 2066
rect -1487 2059 -1485 2061
rect -1482 2059 -1480 2061
rect -1487 2054 -1485 2056
rect -1482 2054 -1480 2056
rect -1487 2049 -1485 2051
rect -1482 2049 -1480 2051
rect -1487 2044 -1485 2046
rect -1482 2044 -1480 2046
rect -1487 2039 -1485 2041
rect -1482 2039 -1480 2041
rect -1487 2034 -1485 2036
rect -1482 2034 -1480 2036
rect -1487 2029 -1485 2031
rect -1482 2029 -1480 2031
rect -1487 2024 -1485 2026
rect -1482 2024 -1480 2026
rect -1487 2019 -1485 2021
rect -1482 2019 -1480 2021
rect -1487 2014 -1485 2016
rect -1482 2014 -1480 2016
rect 3289 2012 3291 2014
rect -1487 2009 -1485 2011
rect -1482 2009 -1480 2011
rect -1487 2004 -1485 2006
rect -1482 2004 -1480 2006
rect 3279 1794 3281 1796
rect 3284 1794 3286 1796
rect 3279 1789 3281 1791
rect 3284 1789 3286 1791
rect 3279 1784 3281 1786
rect 3284 1784 3286 1786
rect 3279 1779 3281 1781
rect 3284 1779 3286 1781
rect 3279 1774 3281 1776
rect 3284 1774 3286 1776
rect 3279 1769 3281 1771
rect 3284 1769 3286 1771
rect 3279 1764 3281 1766
rect 3284 1764 3286 1766
rect 3279 1759 3281 1761
rect 3284 1759 3286 1761
rect 3279 1754 3281 1756
rect 3284 1754 3286 1756
rect 3279 1749 3281 1751
rect 3284 1749 3286 1751
rect 3279 1744 3281 1746
rect 3284 1744 3286 1746
rect 3279 1739 3281 1741
rect 3284 1739 3286 1741
rect 3279 1734 3281 1736
rect 3284 1734 3286 1736
rect 3279 1729 3281 1731
rect 3284 1729 3286 1731
rect 3279 1724 3281 1726
rect 3284 1724 3286 1726
rect 3279 1719 3281 1721
rect 3284 1719 3286 1721
rect 3279 1714 3281 1716
rect 3284 1714 3286 1716
rect 3279 1709 3281 1711
rect 3284 1709 3286 1711
rect 3279 1704 3281 1706
rect 3284 1704 3286 1706
rect 3289 1412 3291 1414
rect 3267 1350 3269 1352
rect 3272 1350 3274 1352
rect 3277 1350 3279 1352
rect 3267 1345 3269 1347
rect 3272 1345 3274 1347
rect 3277 1345 3279 1347
rect -1486 1263 -1484 1265
rect -1486 1258 -1484 1260
rect -1491 1112 -1489 1114
rect -1226 1111 -1224 1113
rect 3289 1112 3291 1114
rect 3268 1050 3270 1052
rect 3273 1050 3275 1052
rect 3278 1050 3280 1052
rect 3268 1045 3270 1047
rect 3273 1045 3275 1047
rect 3278 1045 3280 1047
rect 3289 812 3291 814
rect 3267 750 3269 752
rect 3272 750 3274 752
rect 3277 750 3279 752
rect 3267 745 3269 747
rect 3272 745 3274 747
rect 3277 745 3279 747
rect 3289 512 3291 514
rect 3267 450 3269 452
rect 3272 450 3274 452
rect 3277 450 3279 452
rect 3267 445 3269 447
rect 3272 445 3274 447
rect 3277 445 3279 447
rect -1488 294 -1486 296
rect -1483 294 -1481 296
rect -1488 289 -1486 291
rect -1483 289 -1481 291
rect -1488 284 -1486 286
rect -1483 284 -1481 286
rect -1488 279 -1486 281
rect -1483 279 -1481 281
rect -1488 274 -1486 276
rect -1483 274 -1481 276
rect -1488 269 -1486 271
rect -1483 269 -1481 271
rect -1488 264 -1486 266
rect -1483 264 -1481 266
rect -1488 259 -1486 261
rect -1483 259 -1481 261
rect -1488 254 -1486 256
rect -1483 254 -1481 256
rect -1488 249 -1486 251
rect -1483 249 -1481 251
rect -1488 244 -1486 246
rect -1483 244 -1481 246
rect -1488 239 -1486 241
rect -1483 239 -1481 241
rect -1488 234 -1486 236
rect -1483 234 -1481 236
rect -1488 229 -1486 231
rect -1483 229 -1481 231
rect -1488 224 -1486 226
rect -1483 224 -1481 226
rect -1488 219 -1486 221
rect -1483 219 -1481 221
rect -1488 214 -1486 216
rect -1483 214 -1481 216
rect 3289 212 3291 214
rect -1488 209 -1486 211
rect -1483 209 -1481 211
rect -1488 204 -1486 206
rect -1483 204 -1481 206
rect 3267 150 3269 152
rect 3272 150 3274 152
rect 3277 150 3279 152
rect 3267 145 3269 147
rect 3272 145 3274 147
rect 3277 145 3279 147
rect 3285 -6 3287 -4
rect 3285 -11 3287 -9
rect 3285 -16 3287 -14
rect 3285 -21 3287 -19
rect 3285 -26 3287 -24
rect 3285 -31 3287 -29
rect 3285 -36 3287 -34
rect 3285 -41 3287 -39
rect 3285 -46 3287 -44
rect 3285 -51 3287 -49
rect 3285 -56 3287 -54
rect 3285 -61 3287 -59
rect 3285 -66 3287 -64
rect 3285 -71 3287 -69
rect 3285 -76 3287 -74
rect 3285 -81 3287 -79
rect 3285 -86 3287 -84
rect 3285 -91 3287 -89
rect 3285 -96 3287 -94
rect 3289 -388 3291 -386
rect 3268 -450 3270 -448
rect 3273 -450 3275 -448
rect 3278 -450 3280 -448
rect 3268 -455 3270 -453
rect 3273 -455 3275 -453
rect 3278 -455 3280 -453
rect 3289 -688 3291 -686
rect 3267 -750 3269 -748
rect 3272 -750 3274 -748
rect 3277 -750 3279 -748
rect 3267 -755 3269 -753
rect 3272 -755 3274 -753
rect 3277 -755 3279 -753
rect -196 -1372 -194 -1370
rect -191 -1372 -189 -1370
rect -186 -1372 -184 -1370
rect -181 -1372 -179 -1370
rect -176 -1372 -174 -1370
rect -171 -1372 -169 -1370
rect -166 -1372 -164 -1370
rect -161 -1372 -159 -1370
rect -156 -1372 -154 -1370
rect -151 -1372 -149 -1370
rect -146 -1372 -144 -1370
rect -141 -1372 -139 -1370
rect -136 -1372 -134 -1370
rect -131 -1372 -129 -1370
rect -126 -1372 -124 -1370
rect -121 -1372 -119 -1370
rect -116 -1372 -114 -1370
rect -111 -1372 -109 -1370
rect -106 -1372 -104 -1370
rect -196 -1377 -194 -1375
rect -191 -1377 -189 -1375
rect -186 -1377 -184 -1375
rect -181 -1377 -179 -1375
rect -176 -1377 -174 -1375
rect -171 -1377 -169 -1375
rect -166 -1377 -164 -1375
rect -161 -1377 -159 -1375
rect -156 -1377 -154 -1375
rect -151 -1377 -149 -1375
rect -146 -1377 -144 -1375
rect -141 -1377 -139 -1375
rect -136 -1377 -134 -1375
rect -131 -1377 -129 -1375
rect -126 -1377 -124 -1375
rect -121 -1377 -119 -1375
rect -116 -1377 -114 -1375
rect -111 -1377 -109 -1375
rect -106 -1377 -104 -1375
rect 1604 -1378 1606 -1376
rect 1609 -1378 1611 -1376
rect 1614 -1378 1616 -1376
rect 1619 -1378 1621 -1376
rect 1624 -1378 1626 -1376
rect 1629 -1378 1631 -1376
rect 1634 -1378 1636 -1376
rect 1639 -1378 1641 -1376
rect 1644 -1378 1646 -1376
rect 1649 -1378 1651 -1376
rect 1654 -1378 1656 -1376
rect 1659 -1378 1661 -1376
rect 1664 -1378 1666 -1376
rect 1669 -1378 1671 -1376
rect 1674 -1378 1676 -1376
rect 1679 -1378 1681 -1376
rect 1684 -1378 1686 -1376
rect 1689 -1378 1691 -1376
rect 1694 -1378 1696 -1376
rect -196 -1382 -194 -1380
rect -191 -1382 -189 -1380
rect -186 -1382 -184 -1380
rect -181 -1382 -179 -1380
rect -176 -1382 -174 -1380
rect -171 -1382 -169 -1380
rect -166 -1382 -164 -1380
rect -161 -1382 -159 -1380
rect -156 -1382 -154 -1380
rect -151 -1382 -149 -1380
rect -146 -1382 -144 -1380
rect -141 -1382 -139 -1380
rect -136 -1382 -134 -1380
rect -131 -1382 -129 -1380
rect -126 -1382 -124 -1380
rect -121 -1382 -119 -1380
rect -116 -1382 -114 -1380
rect -111 -1382 -109 -1380
rect -106 -1382 -104 -1380
rect 1604 -1383 1606 -1381
rect 1609 -1383 1611 -1381
rect 1614 -1383 1616 -1381
rect 1619 -1383 1621 -1381
rect 1624 -1383 1626 -1381
rect 1629 -1383 1631 -1381
rect 1634 -1383 1636 -1381
rect 1639 -1383 1641 -1381
rect 1644 -1383 1646 -1381
rect 1649 -1383 1651 -1381
rect 1654 -1383 1656 -1381
rect 1659 -1383 1661 -1381
rect 1664 -1383 1666 -1381
rect 1669 -1383 1671 -1381
rect 1674 -1383 1676 -1381
rect 1679 -1383 1681 -1381
rect 1684 -1383 1686 -1381
rect 1689 -1383 1691 -1381
rect 1694 -1383 1696 -1381
rect -196 -1387 -194 -1385
rect -191 -1387 -189 -1385
rect -186 -1387 -184 -1385
rect -181 -1387 -179 -1385
rect -176 -1387 -174 -1385
rect -171 -1387 -169 -1385
rect -166 -1387 -164 -1385
rect -161 -1387 -159 -1385
rect -156 -1387 -154 -1385
rect -151 -1387 -149 -1385
rect -146 -1387 -144 -1385
rect -141 -1387 -139 -1385
rect -136 -1387 -134 -1385
rect -131 -1387 -129 -1385
rect -126 -1387 -124 -1385
rect -121 -1387 -119 -1385
rect -116 -1387 -114 -1385
rect -111 -1387 -109 -1385
rect -106 -1387 -104 -1385
rect 1604 -1388 1606 -1386
rect 1609 -1388 1611 -1386
rect 1614 -1388 1616 -1386
rect 1619 -1388 1621 -1386
rect 1624 -1388 1626 -1386
rect 1629 -1388 1631 -1386
rect 1634 -1388 1636 -1386
rect 1639 -1388 1641 -1386
rect 1644 -1388 1646 -1386
rect 1649 -1388 1651 -1386
rect 1654 -1388 1656 -1386
rect 1659 -1388 1661 -1386
rect 1664 -1388 1666 -1386
rect 1669 -1388 1671 -1386
rect 1674 -1388 1676 -1386
rect 1679 -1388 1681 -1386
rect 1684 -1388 1686 -1386
rect 1689 -1388 1691 -1386
rect 1694 -1388 1696 -1386
<< metal3 >>
rect -1478 3341 -1470 3385
rect -1407 3341 -1399 3393
rect -1178 3341 -1170 3384
rect -1106 3341 -1100 3393
rect -878 3341 -870 3384
rect -806 3341 -800 3393
rect -578 3341 -570 3385
rect -506 3341 -500 3393
rect -278 3341 -270 3384
rect -206 3341 -200 3393
rect 22 3341 30 3384
rect 94 3341 100 3393
rect 622 3341 630 3384
rect 694 3341 700 3395
rect 922 3341 930 3384
rect 994 3341 1000 3393
rect 1222 3341 1230 3385
rect 1294 3341 1300 3393
rect 1522 3341 1530 3385
rect 1594 3341 1600 3383
rect 1822 3341 1830 3385
rect 1894 3341 1900 3389
rect 2122 3341 2130 3384
rect 2194 3341 2200 3393
rect 2722 3341 2730 3385
rect 2794 3341 2800 3391
rect 3022 3341 3030 3384
rect 3094 3341 3100 3391
rect -1478 3334 3246 3341
rect -1454 3289 3246 3334
rect -1454 3288 -1293 3289
rect -1454 3201 -1396 3288
rect -1313 3201 -1299 3288
rect -1493 3193 -1299 3201
rect 3175 3200 3246 3289
rect 3175 3194 3293 3200
rect -1454 3130 -1396 3193
rect -1484 3122 -1396 3130
rect -1454 2830 -1396 3122
rect -1483 2822 -1396 2830
rect -1454 2530 -1396 2822
rect -1483 2522 -1396 2530
rect -1454 2230 -1396 2522
rect -1483 2222 -1396 2230
rect -1454 2099 -1396 2222
rect 3175 3130 3246 3194
rect 3175 3122 3284 3130
rect 3175 2900 3246 3122
rect 3175 2894 3293 2900
rect 3175 2830 3246 2894
rect 3175 2822 3283 2830
rect 3175 2600 3246 2822
rect 3175 2594 3293 2600
rect 3175 2300 3246 2594
rect 3175 2294 3293 2300
rect 3175 2230 3246 2294
rect 3175 2222 3283 2230
rect 3000 2149 3007 2156
rect 3000 2119 3007 2126
rect 3000 2099 3007 2106
rect -1479 2001 -1396 2099
rect -1454 1100 -1396 2001
rect 3175 2000 3246 2222
rect 3175 1994 3293 2000
rect 3175 1930 3246 1994
rect 3175 1922 3283 1930
rect 3175 1799 3246 1922
rect 3175 1752 3277 1799
rect 2948 1701 3277 1752
rect 2948 1665 3246 1701
rect 3175 1400 3246 1665
rect 3175 1394 3293 1400
rect -1221 1109 -1214 1116
rect -1493 1094 -1396 1100
rect -1454 1030 -1396 1094
rect -1484 1022 -1396 1030
rect -1454 730 -1396 1022
rect -1484 722 -1396 730
rect -1454 430 -1396 722
rect -1484 422 -1396 430
rect -1454 299 -1396 422
rect -1481 201 -1396 299
rect -1454 78 -1396 201
rect -1483 70 -1396 78
rect -1454 -470 -1396 70
rect 3175 1100 3246 1394
rect 3175 1094 3293 1100
rect 3175 800 3246 1094
rect 3175 794 3293 800
rect 3175 500 3246 794
rect 3175 494 3293 500
rect 3175 200 3246 494
rect 3175 194 3293 200
rect 3175 -1 3246 194
rect 3175 -49 3284 -1
rect 2947 -99 3284 -49
rect 2947 -137 3246 -99
rect -1483 -478 -1396 -470
rect -1454 -770 -1396 -478
rect -1484 -778 -1396 -770
rect -1454 -1070 -1396 -778
rect -1484 -1078 -1396 -1070
rect -1454 -1294 -1396 -1078
rect 3175 -400 3246 -137
rect 3175 -406 3293 -400
rect 3175 -700 3246 -406
rect 3175 -706 3293 -700
rect 3175 -1070 3246 -706
rect 3175 -1078 3283 -1070
rect 3175 -1294 3246 -1078
rect -1454 -1351 3246 -1294
rect -1444 -1370 -1439 -1351
rect -1483 -1375 -1439 -1370
rect -1483 -1383 -1470 -1375
rect -1178 -1383 -1170 -1351
rect -878 -1383 -870 -1351
rect -578 -1383 -570 -1351
rect 22 -1383 30 -1351
rect 322 -1383 330 -1351
rect 622 -1383 630 -1351
rect 922 -1383 930 -1351
rect 1222 -1383 1230 -1351
rect 1822 -1383 1830 -1351
rect 2122 -1383 2130 -1351
rect 2422 -1383 2430 -1351
rect 2722 -1383 2730 -1351
rect 3022 -1383 3030 -1351
rect 3237 -1370 3246 -1351
rect 3237 -1378 3284 -1370
<< gv2 >>
rect -1404 3389 -1402 3391
rect -1104 3389 -1102 3391
rect -804 3389 -802 3391
rect -504 3388 -502 3390
rect -204 3389 -202 3391
rect 96 3389 98 3391
rect 696 3389 698 3391
rect 996 3389 998 3391
rect 1296 3389 1298 3391
rect 2196 3389 2198 3391
rect 2796 3387 2798 3389
rect 3096 3387 3098 3389
rect 1896 3385 1898 3387
rect -1475 3380 -1473 3382
rect -1175 3379 -1173 3381
rect -875 3379 -873 3381
rect -575 3380 -573 3382
rect -275 3379 -273 3381
rect 25 3379 27 3381
rect 625 3379 627 3381
rect 925 3379 927 3381
rect 1225 3380 1227 3382
rect 1525 3379 1527 3381
rect 1825 3380 1827 3382
rect 1596 3378 1598 3380
rect 2125 3379 2127 3381
rect 2725 3379 2727 3381
rect 3025 3379 3027 3381
rect -1491 3196 -1489 3198
rect 3289 3196 3291 3198
rect -1482 3125 -1480 3127
rect 3279 3125 3281 3127
rect 3289 2896 3291 2898
rect -1480 2825 -1478 2827
rect 3278 2825 3280 2827
rect 3289 2596 3291 2598
rect -1480 2525 -1478 2527
rect 3289 2296 3291 2298
rect -1480 2225 -1478 2227
rect 3278 2225 3280 2227
rect 3002 2151 3004 2153
rect 3002 2121 3004 2123
rect 3002 2101 3004 2103
rect -1476 2094 -1474 2096
rect -1471 2094 -1469 2096
rect -1476 2089 -1474 2091
rect -1471 2089 -1469 2091
rect -1476 2084 -1474 2086
rect -1471 2084 -1469 2086
rect -1476 2079 -1474 2081
rect -1471 2079 -1469 2081
rect -1476 2074 -1474 2076
rect -1471 2074 -1469 2076
rect -1476 2069 -1474 2071
rect -1471 2069 -1469 2071
rect -1476 2064 -1474 2066
rect -1471 2064 -1469 2066
rect -1476 2059 -1474 2061
rect -1471 2059 -1469 2061
rect -1476 2054 -1474 2056
rect -1471 2054 -1469 2056
rect -1476 2049 -1474 2051
rect -1471 2049 -1469 2051
rect -1476 2044 -1474 2046
rect -1471 2044 -1469 2046
rect -1476 2039 -1474 2041
rect -1471 2039 -1469 2041
rect -1476 2034 -1474 2036
rect -1471 2034 -1469 2036
rect -1476 2029 -1474 2031
rect -1471 2029 -1469 2031
rect -1476 2024 -1474 2026
rect -1471 2024 -1469 2026
rect -1476 2019 -1474 2021
rect -1471 2019 -1469 2021
rect -1476 2014 -1474 2016
rect -1471 2014 -1469 2016
rect -1476 2009 -1474 2011
rect -1471 2009 -1469 2011
rect -1476 2004 -1474 2006
rect -1471 2004 -1469 2006
rect 3289 1996 3291 1998
rect 3278 1925 3280 1927
rect 3257 1794 3259 1796
rect 3262 1794 3264 1796
rect 3267 1794 3269 1796
rect 3272 1794 3274 1796
rect 3257 1789 3259 1791
rect 3262 1789 3264 1791
rect 3267 1789 3269 1791
rect 3272 1789 3274 1791
rect 3257 1784 3259 1786
rect 3262 1784 3264 1786
rect 3267 1784 3269 1786
rect 3272 1784 3274 1786
rect 3257 1779 3259 1781
rect 3262 1779 3264 1781
rect 3267 1779 3269 1781
rect 3272 1779 3274 1781
rect 3257 1774 3259 1776
rect 3262 1774 3264 1776
rect 3267 1774 3269 1776
rect 3272 1774 3274 1776
rect 3257 1769 3259 1771
rect 3262 1769 3264 1771
rect 3267 1769 3269 1771
rect 3272 1769 3274 1771
rect 3257 1764 3259 1766
rect 3262 1764 3264 1766
rect 3267 1764 3269 1766
rect 3272 1764 3274 1766
rect 3257 1759 3259 1761
rect 3262 1759 3264 1761
rect 3267 1759 3269 1761
rect 3272 1759 3274 1761
rect 3257 1754 3259 1756
rect 3262 1754 3264 1756
rect 3267 1754 3269 1756
rect 3272 1754 3274 1756
rect 3257 1749 3259 1751
rect 3262 1749 3264 1751
rect 3267 1749 3269 1751
rect 3272 1749 3274 1751
rect 2951 1747 2953 1749
rect 2956 1747 2958 1749
rect 2961 1747 2963 1749
rect 3257 1744 3259 1746
rect 3262 1744 3264 1746
rect 3267 1744 3269 1746
rect 3272 1744 3274 1746
rect 2951 1742 2953 1744
rect 2956 1742 2958 1744
rect 2961 1742 2963 1744
rect 3257 1739 3259 1741
rect 3262 1739 3264 1741
rect 3267 1739 3269 1741
rect 3272 1739 3274 1741
rect 2951 1737 2953 1739
rect 2956 1737 2958 1739
rect 2961 1737 2963 1739
rect 3257 1734 3259 1736
rect 3262 1734 3264 1736
rect 3267 1734 3269 1736
rect 3272 1734 3274 1736
rect 2951 1732 2953 1734
rect 2956 1732 2958 1734
rect 2961 1732 2963 1734
rect 3257 1729 3259 1731
rect 3262 1729 3264 1731
rect 3267 1729 3269 1731
rect 3272 1729 3274 1731
rect 2951 1727 2953 1729
rect 2956 1727 2958 1729
rect 2961 1727 2963 1729
rect 3257 1724 3259 1726
rect 3262 1724 3264 1726
rect 3267 1724 3269 1726
rect 3272 1724 3274 1726
rect 2951 1722 2953 1724
rect 2956 1722 2958 1724
rect 2961 1722 2963 1724
rect 3257 1719 3259 1721
rect 3262 1719 3264 1721
rect 3267 1719 3269 1721
rect 3272 1719 3274 1721
rect 2951 1717 2953 1719
rect 2956 1717 2958 1719
rect 2961 1717 2963 1719
rect 3257 1714 3259 1716
rect 3262 1714 3264 1716
rect 3267 1714 3269 1716
rect 3272 1714 3274 1716
rect 2951 1712 2953 1714
rect 2956 1712 2958 1714
rect 2961 1712 2963 1714
rect 3257 1709 3259 1711
rect 3262 1709 3264 1711
rect 3267 1709 3269 1711
rect 3272 1709 3274 1711
rect 2951 1707 2953 1709
rect 2956 1707 2958 1709
rect 2961 1707 2963 1709
rect 3257 1704 3259 1706
rect 3262 1704 3264 1706
rect 3267 1704 3269 1706
rect 3272 1704 3274 1706
rect 2951 1702 2953 1704
rect 2956 1702 2958 1704
rect 2961 1702 2963 1704
rect 2951 1697 2953 1699
rect 2956 1697 2958 1699
rect 2961 1697 2963 1699
rect 2951 1692 2953 1694
rect 2956 1692 2958 1694
rect 2961 1692 2963 1694
rect 2951 1687 2953 1689
rect 2956 1687 2958 1689
rect 2961 1687 2963 1689
rect 2951 1682 2953 1684
rect 2956 1682 2958 1684
rect 2961 1682 2963 1684
rect 2951 1677 2953 1679
rect 2956 1677 2958 1679
rect 2961 1677 2963 1679
rect 2951 1672 2953 1674
rect 2956 1672 2958 1674
rect 2961 1672 2963 1674
rect 2951 1667 2953 1669
rect 2956 1667 2958 1669
rect 2961 1667 2963 1669
rect 3289 1396 3291 1398
rect -1219 1111 -1217 1113
rect -1491 1096 -1489 1098
rect 3289 1096 3291 1098
rect -1482 1025 -1480 1027
rect 3289 796 3291 798
rect -1482 725 -1480 727
rect 3289 496 3291 498
rect -1482 425 -1480 427
rect -1479 294 -1477 296
rect -1474 294 -1472 296
rect -1479 289 -1477 291
rect -1474 289 -1472 291
rect -1479 284 -1477 286
rect -1474 284 -1472 286
rect -1479 279 -1477 281
rect -1474 279 -1472 281
rect -1479 274 -1477 276
rect -1474 274 -1472 276
rect -1479 269 -1477 271
rect -1474 269 -1472 271
rect -1479 264 -1477 266
rect -1474 264 -1472 266
rect -1479 259 -1477 261
rect -1474 259 -1472 261
rect -1479 254 -1477 256
rect -1474 254 -1472 256
rect -1479 249 -1477 251
rect -1474 249 -1472 251
rect -1479 244 -1477 246
rect -1474 244 -1472 246
rect -1479 239 -1477 241
rect -1474 239 -1472 241
rect -1479 234 -1477 236
rect -1474 234 -1472 236
rect -1479 229 -1477 231
rect -1474 229 -1472 231
rect -1479 224 -1477 226
rect -1474 224 -1472 226
rect -1479 219 -1477 221
rect -1474 219 -1472 221
rect -1479 214 -1477 216
rect -1474 214 -1472 216
rect -1479 209 -1477 211
rect -1474 209 -1472 211
rect -1479 204 -1477 206
rect -1474 204 -1472 206
rect 3289 196 3291 198
rect -1480 73 -1478 75
rect 3279 -6 3281 -4
rect 3279 -11 3281 -9
rect 3279 -16 3281 -14
rect 3279 -21 3281 -19
rect 3279 -26 3281 -24
rect 3279 -31 3281 -29
rect 3279 -36 3281 -34
rect 3279 -41 3281 -39
rect 3279 -46 3281 -44
rect 3279 -51 3281 -49
rect 2951 -54 2953 -52
rect 2956 -54 2958 -52
rect 2961 -54 2963 -52
rect 3279 -56 3281 -54
rect 2951 -59 2953 -57
rect 2956 -59 2958 -57
rect 2961 -59 2963 -57
rect 3279 -61 3281 -59
rect 2951 -64 2953 -62
rect 2956 -64 2958 -62
rect 2961 -64 2963 -62
rect 3279 -66 3281 -64
rect 2951 -69 2953 -67
rect 2956 -69 2958 -67
rect 2961 -69 2963 -67
rect 3279 -71 3281 -69
rect 2951 -74 2953 -72
rect 2956 -74 2958 -72
rect 2961 -74 2963 -72
rect 3279 -76 3281 -74
rect 2951 -79 2953 -77
rect 2956 -79 2958 -77
rect 2961 -79 2963 -77
rect 3279 -81 3281 -79
rect 2951 -84 2953 -82
rect 2956 -84 2958 -82
rect 2961 -84 2963 -82
rect 3279 -86 3281 -84
rect 2951 -89 2953 -87
rect 2956 -89 2958 -87
rect 2961 -89 2963 -87
rect 3279 -91 3281 -89
rect 2951 -94 2953 -92
rect 2956 -94 2958 -92
rect 2961 -94 2963 -92
rect 3279 -96 3281 -94
rect 2951 -99 2953 -97
rect 2956 -99 2958 -97
rect 2961 -99 2963 -97
rect 2951 -104 2953 -102
rect 2956 -104 2958 -102
rect 2961 -104 2963 -102
rect 2951 -109 2953 -107
rect 2956 -109 2958 -107
rect 2961 -109 2963 -107
rect 2951 -114 2953 -112
rect 2956 -114 2958 -112
rect 2961 -114 2963 -112
rect 2951 -119 2953 -117
rect 2956 -119 2958 -117
rect 2961 -119 2963 -117
rect 2951 -124 2953 -122
rect 2956 -124 2958 -122
rect 2961 -124 2963 -122
rect 2951 -129 2953 -127
rect 2956 -129 2958 -127
rect 2961 -129 2963 -127
rect 2951 -134 2953 -132
rect 2956 -134 2958 -132
rect 2961 -134 2963 -132
rect 3289 -404 3291 -402
rect -1480 -475 -1478 -473
rect 3289 -704 3291 -702
rect -1481 -775 -1479 -773
rect -1481 -1075 -1479 -1073
rect 3278 -1075 3280 -1073
rect -1480 -1375 -1478 -1373
rect -1475 -1375 -1473 -1373
rect 3279 -1375 3281 -1373
rect -1480 -1380 -1478 -1378
rect -1475 -1380 -1473 -1378
rect -1175 -1380 -1173 -1378
rect -875 -1380 -873 -1378
rect -575 -1380 -573 -1378
rect 25 -1380 27 -1378
rect 325 -1380 327 -1378
rect 625 -1380 627 -1378
rect 925 -1380 927 -1378
rect 1225 -1380 1227 -1378
rect 1825 -1380 1827 -1378
rect 2125 -1380 2127 -1378
rect 2425 -1380 2427 -1378
rect 2725 -1380 2727 -1378
rect 3025 -1380 3027 -1378
use top_level  top_level_0
timestamp 1682896469
transform 1 0 -1220 0 1 -1212
box 0 12 4226 4140
use PadFrame64  PadFrame64_0
timestamp 1682896469
transform 1 0 0 0 1 0
box -2500 -2400 4300 4400
<< labels >>
rlabel metal2 3282 3361 3282 3361 6 17_17_DI
rlabel metal2 3282 3348 3282 3348 6 17_17_DIB
rlabel metal1 -2206 249 -2206 249 4 Gnd!
rlabel metal1 447 4108 447 4108 6 Vdd!
rlabel metal1 -2207 2051 -2207 2051 4 Gnd!
rlabel metal1 -2212 1154 -2212 1154 4 p_clkb
rlabel metal1 -2212 3250 -2212 3250 4 p_load[8]
rlabel metal1 -1352 4113 -1352 4113 4 p_load[0]
rlabel metal1 -1047 4106 -1047 4106 4 p_load[14]
rlabel metal1 -753 4109 -753 4109 4 p_load[12]
rlabel metal1 -448 4112 -448 4112 4 p_load[13]
rlabel metal1 -145 4112 -145 4112 4 p_load[9]
rlabel metal1 153 4115 153 4115 6 p_load[7]
rlabel metal1 754 4109 754 4109 6 p_load[3]
rlabel metal1 1055 4112 1055 4112 6 p_load[10]
rlabel metal1 1353 4109 1353 4109 6 p_load[5]
rlabel metal1 1660 4112 1660 4112 6 p_load[11]
rlabel metal1 1952 4114 1952 4114 6 p_load[6]
rlabel metal1 2254 4113 2254 4113 6 p_load[15]
rlabel metal1 2549 4110 2549 4110 6 Vdd!
rlabel metal1 2846 4106 2846 4106 6 p_load[2]
rlabel metal1 3145 4106 3145 4106 6 p_load[1]
rlabel metal1 4006 3244 4006 3244 6 p_we_ins
rlabel metal1 4001 2946 4001 2946 6 p_load[4]
rlabel metal1 4010 2655 4010 2655 6 p_reg_0_out[7]
rlabel metal1 4011 2345 4011 2345 6 p_clka
rlabel metal1 4015 2053 4015 2053 6 p_reset
rlabel metal1 4013 1453 4013 1453 6 p_reg_0_out[1]
rlabel metal1 4007 1757 4007 1757 6 Gnd!
rlabel metal1 4013 1151 4013 1151 6 p_reg_0_out[0]
rlabel metal1 4008 848 4008 848 6 p_reg_0_out[6]
rlabel metal1 4008 557 4008 557 6 p_reg_0_out[2]
rlabel metal1 4007 253 4007 253 6 p_reg_0_out[3]
rlabel metal1 4008 -350 4008 -350 8 p_reg_0_out[5]
rlabel metal1 4009 -645 4009 -645 8 p_reg_0_out[4]
rlabel metal1 4002 -48 4002 -48 8 Gnd!
<< end >>

magic
tech scmos
timestamp 1680363874
<< nwell >>
rect -5 48 126 105
rect 23 46 100 48
rect 65 39 100 46
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
rect 31 6 33 26
rect 36 6 38 26
rect 44 6 46 26
rect 52 6 54 26
rect 60 6 62 26
rect 68 6 70 26
rect 77 6 79 26
rect 82 6 84 26
rect 87 6 89 26
rect 95 6 97 16
rect 111 6 113 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
rect 36 54 38 94
rect 44 54 46 94
rect 52 58 54 94
rect 60 58 62 94
rect 68 58 70 94
rect 77 46 79 94
rect 82 46 84 94
rect 87 46 89 94
rect 95 74 97 94
rect 111 74 113 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 20 15 26
rect 9 6 10 20
rect 14 6 15 20
rect 17 25 23 26
rect 17 6 18 25
rect 22 6 23 25
rect 25 21 31 26
rect 25 7 26 21
rect 30 7 31 21
rect 25 6 31 7
rect 33 6 36 26
rect 38 22 44 26
rect 38 8 39 22
rect 43 8 44 22
rect 38 6 44 8
rect 46 25 52 26
rect 46 6 47 25
rect 51 6 52 25
rect 54 17 60 26
rect 54 8 55 17
rect 59 8 60 17
rect 54 6 60 8
rect 62 25 68 26
rect 62 6 63 25
rect 67 6 68 25
rect 70 20 77 26
rect 70 6 71 20
rect 75 6 77 20
rect 79 6 82 26
rect 84 6 87 26
rect 89 25 94 26
rect 89 6 90 25
rect 94 6 95 16
rect 97 15 102 16
rect 97 6 98 15
rect 106 15 111 16
rect 110 6 111 15
rect 113 15 118 16
rect 113 6 114 15
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 60 10 94
rect 14 60 15 94
rect 9 54 15 60
rect 17 93 23 94
rect 17 54 18 93
rect 22 54 23 93
rect 25 93 31 94
rect 25 59 26 93
rect 30 59 31 93
rect 25 54 31 59
rect 33 54 36 94
rect 38 93 44 94
rect 38 54 39 93
rect 43 54 44 93
rect 46 93 52 94
rect 46 54 47 93
rect 51 58 52 93
rect 54 93 60 94
rect 54 64 55 93
rect 59 64 60 93
rect 54 58 60 64
rect 62 93 68 94
rect 62 59 63 93
rect 67 59 68 93
rect 62 58 68 59
rect 70 92 77 94
rect 70 58 71 92
rect 75 53 77 92
rect 71 51 77 53
rect 72 47 77 51
rect 74 46 77 47
rect 79 46 82 94
rect 84 46 87 94
rect 89 92 95 94
rect 89 48 90 92
rect 94 74 95 92
rect 97 93 102 94
rect 97 74 98 93
rect 106 93 111 94
rect 110 74 111 93
rect 113 93 118 94
rect 113 74 114 93
rect 89 46 94 48
<< ndcontact >>
rect 2 6 6 25
rect 10 6 14 20
rect 18 6 22 25
rect 26 7 30 21
rect 39 8 43 22
rect 47 6 51 25
rect 55 8 59 17
rect 63 6 67 25
rect 71 6 75 20
rect 90 6 94 25
rect 98 6 102 15
rect 106 6 110 15
rect 114 6 118 15
<< pdcontact >>
rect 2 54 6 93
rect 10 60 14 94
rect 18 54 22 93
rect 26 59 30 93
rect 39 54 43 93
rect 47 54 51 93
rect 55 64 59 93
rect 63 59 67 93
rect 71 53 75 92
rect 90 48 94 92
rect 98 74 102 93
rect 106 74 110 93
rect 114 74 118 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
rect 94 -2 98 2
rect 110 -2 114 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
rect 94 98 98 102
rect 110 98 114 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 36 94 38 96
rect 44 94 46 96
rect 52 94 54 96
rect 60 94 62 96
rect 68 94 70 96
rect 77 94 79 96
rect 82 94 84 96
rect 87 94 89 96
rect 95 94 97 96
rect 111 94 113 96
rect 7 33 9 54
rect 15 39 17 54
rect 23 47 25 54
rect 7 26 9 29
rect 15 26 17 35
rect 23 26 25 43
rect 31 39 33 54
rect 36 53 38 54
rect 44 53 46 54
rect 52 53 54 58
rect 60 57 62 58
rect 68 57 70 58
rect 36 51 46 53
rect 49 51 54 53
rect 57 55 62 57
rect 66 55 70 57
rect 31 26 33 35
rect 37 32 39 51
rect 49 38 51 51
rect 57 45 59 55
rect 66 51 68 55
rect 51 34 54 36
rect 36 28 37 29
rect 41 28 46 29
rect 36 27 46 28
rect 36 26 38 27
rect 44 26 46 27
rect 52 26 54 34
rect 57 29 59 41
rect 66 29 68 47
rect 95 73 97 74
rect 95 71 99 73
rect 77 44 79 46
rect 76 42 79 44
rect 74 29 76 40
rect 82 38 84 46
rect 87 44 89 46
rect 87 42 91 44
rect 57 27 62 29
rect 66 27 70 29
rect 74 27 79 29
rect 60 26 62 27
rect 68 26 70 27
rect 77 26 79 27
rect 82 26 84 34
rect 89 38 91 42
rect 97 39 99 71
rect 111 57 113 74
rect 112 53 113 57
rect 89 30 91 34
rect 87 28 91 30
rect 87 26 89 28
rect 97 25 99 35
rect 95 23 99 25
rect 95 16 97 23
rect 111 16 113 53
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
rect 36 4 38 6
rect 44 4 46 6
rect 52 4 54 6
rect 60 4 62 6
rect 68 4 70 6
rect 77 4 79 6
rect 82 4 84 6
rect 87 4 89 6
rect 95 4 97 6
rect 111 4 113 6
<< polycontact >>
rect 22 43 26 47
rect 14 35 18 39
rect 6 29 10 33
rect 29 35 33 39
rect 64 47 68 51
rect 55 41 59 45
rect 47 34 51 38
rect 37 28 41 32
rect 72 40 76 44
rect 80 34 84 38
rect 108 53 112 57
rect 89 34 93 38
rect 97 35 101 39
<< metal1 >>
rect -2 102 122 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 62 102
rect 66 98 78 102
rect 82 98 94 102
rect 98 98 110 102
rect 114 98 122 102
rect -2 97 122 98
rect 10 94 14 97
rect 2 93 6 94
rect 18 93 22 94
rect 6 54 18 57
rect 26 93 30 94
rect 26 58 30 59
rect 39 93 43 97
rect 47 93 51 94
rect 55 93 59 97
rect 63 93 67 94
rect 51 59 63 61
rect 51 58 67 59
rect 71 92 76 94
rect 75 53 76 92
rect 71 51 76 53
rect 90 92 94 97
rect 98 93 102 94
rect 10 43 14 47
rect 18 43 22 47
rect 90 46 94 48
rect 97 74 98 77
rect 106 93 110 97
rect 114 93 118 94
rect 97 49 100 74
rect 97 46 107 49
rect 26 43 55 46
rect 2 33 6 37
rect 11 36 14 43
rect 52 41 55 43
rect 59 41 72 44
rect 18 35 29 38
rect 33 35 47 38
rect 51 34 80 37
rect 3 30 6 33
rect 10 29 37 32
rect 89 31 92 34
rect 41 28 92 31
rect 104 27 107 46
rect 115 37 118 74
rect 114 33 118 37
rect 2 25 22 26
rect 6 23 18 25
rect 26 21 30 22
rect 26 6 30 7
rect 39 22 43 24
rect 10 3 14 6
rect 39 3 43 8
rect 51 22 63 25
rect 55 17 59 19
rect 55 3 59 8
rect 71 20 76 21
rect 75 6 76 20
rect 104 23 110 27
rect 104 22 107 23
rect 99 19 107 22
rect 99 16 102 19
rect 115 16 118 33
rect 98 15 102 16
rect 106 15 110 16
rect 114 15 118 16
rect 90 3 94 6
rect 106 3 110 6
rect -2 2 122 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 62 2
rect 66 -2 78 2
rect 82 -2 94 2
rect 98 -2 110 2
rect 114 -2 122 2
rect -2 -3 122 -2
<< m2contact >>
rect 26 54 30 58
rect 60 48 64 52
rect 72 47 76 51
rect 104 53 108 57
rect 97 39 101 43
rect 26 22 30 26
rect 72 21 76 25
<< metal2 >>
rect 30 54 104 57
rect 27 26 30 54
rect 60 52 64 54
rect 73 42 76 47
rect 73 39 97 42
rect 73 25 76 39
<< m1p >>
rect 10 43 14 47
rect 18 43 22 47
rect 2 33 6 37
rect 114 33 118 37
rect 106 23 110 27
<< labels >>
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 35 4 35 4 A
rlabel metal1 12 45 12 45 4 B
rlabel metal1 20 45 20 45 4 C
rlabel metal1 116 35 116 35 4 YC
rlabel metal1 108 25 108 25 4 YS
<< end >>

magic
tech scmos
timestamp 1677677812
<< m2contact >>
rect -2 -2 2 2
<< end >>

module pc (
    clka,
    clkb,
    pc_lat_clk,
    reset_in,
    immed_in,
    sr1_out_in,
    pc_out
);
input wire clka, clkb, pc_lat_clk, reset_in;
input wire [5:0] immed_in;
input wire [7:0] sr1_out_in;
output reg [5:0] pc_out;

// TODO: need to fill in

    
endmodule
magic
tech scmos
timestamp 1680363874
<< m2contact >>
rect -2 -2 2 2
<< end >>

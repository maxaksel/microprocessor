magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
rect 20 6 22 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 12 26
rect 14 6 20 26
rect 22 6 27 26
<< pdiffusion >>
rect 2 74 7 94
rect 9 74 15 94
rect 17 74 23 94
rect 18 56 23 74
rect 20 54 23 56
rect 25 54 30 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 73 9 74
rect 5 71 9 73
rect 5 41 7 71
rect 2 37 7 41
rect 15 39 17 74
rect 5 30 7 37
rect 12 37 17 39
rect 12 35 16 37
rect 5 28 9 30
rect 7 26 9 28
rect 12 26 14 35
rect 23 33 25 54
rect 20 31 25 33
rect 20 29 24 31
rect 20 26 22 29
rect 7 4 9 6
rect 12 4 14 6
rect 20 4 22 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 11 90 13 92
rect 19 89 21 91
rect 27 90 29 92
rect 3 85 5 87
rect 11 85 13 87
rect 19 84 21 86
rect 27 85 29 87
rect 3 80 5 82
rect 11 80 13 82
rect 19 79 21 81
rect 27 80 29 82
rect 3 75 5 77
rect 11 75 13 77
rect 19 74 21 76
rect 27 75 29 77
rect 19 69 21 71
rect 27 70 29 72
rect 19 64 21 66
rect 27 65 29 67
rect 19 59 21 61
rect 27 60 29 62
rect 27 55 29 57
rect 3 38 5 40
rect 13 36 15 38
rect 21 30 23 32
rect 3 22 5 24
rect 16 22 18 24
rect 24 22 26 24
rect 3 17 5 19
rect 16 17 18 19
rect 24 17 26 19
rect 3 12 5 14
rect 16 12 18 14
rect 24 12 26 14
rect 3 7 5 9
rect 16 7 18 9
rect 24 7 26 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 34 103
rect 2 74 6 97
rect 10 74 14 94
rect 11 53 14 74
rect 18 56 22 97
rect 26 54 30 94
rect 11 50 23 53
rect 10 43 14 47
rect 2 33 6 41
rect 11 39 14 43
rect 11 36 16 39
rect 12 35 16 36
rect 20 33 23 50
rect 27 47 30 54
rect 26 43 30 47
rect 20 32 24 33
rect 9 30 24 32
rect 3 29 24 30
rect 3 27 12 29
rect 3 26 6 27
rect 27 26 30 43
rect 2 6 6 26
rect 15 3 19 25
rect 23 21 30 26
rect 23 6 27 21
rect -2 -3 34 3
<< m1p >>
rect 10 43 14 47
rect 26 43 30 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 35 4 35 6 A
rlabel metal1 12 45 12 45 6 B
rlabel metal1 28 45 28 45 6 Y
<< end >>

magic
tech scmos
timestamp 1680363874
<< metal1 >>
rect 14 4707 4861 4727
rect 38 4683 4837 4703
rect 14 4667 4861 4673
rect 66 4613 84 4616
rect 228 4613 253 4616
rect 284 4613 301 4616
rect 380 4613 405 4616
rect 436 4613 445 4616
rect 452 4613 461 4616
rect 588 4613 597 4616
rect 604 4613 621 4616
rect 748 4613 765 4616
rect 804 4613 829 4616
rect 860 4613 877 4616
rect 884 4613 908 4616
rect 980 4613 1005 4616
rect 1036 4613 1045 4616
rect 1052 4613 1092 4616
rect 1322 4613 1356 4616
rect 1386 4613 1412 4616
rect 1564 4613 1597 4616
rect 1604 4613 1621 4616
rect 1732 4613 1749 4616
rect 1764 4613 1781 4616
rect 1818 4613 1844 4616
rect 1882 4613 1892 4616
rect 1986 4613 1996 4616
rect 2058 4613 2076 4616
rect 2290 4613 2316 4616
rect 2426 4613 2452 4616
rect 2532 4613 2557 4616
rect 2636 4613 2661 4616
rect 2698 4613 2708 4616
rect 2714 4613 2748 4616
rect 2842 4613 2852 4616
rect 3570 4613 3596 4616
rect 3690 4613 3708 4616
rect 3954 4613 3980 4616
rect 4172 4613 4197 4616
rect 4234 4613 4244 4616
rect 4490 4613 4508 4616
rect 4610 4613 4700 4616
rect 298 4605 301 4613
rect 442 4605 445 4613
rect 594 4605 597 4613
rect 874 4605 877 4613
rect 932 4603 941 4606
rect 1042 4605 1045 4613
rect 1058 4603 1084 4606
rect 1322 4605 1325 4613
rect 38 4567 4837 4573
rect 66 4533 92 4536
rect 164 4533 181 4536
rect 178 4526 181 4533
rect 202 4533 276 4536
rect 356 4533 420 4536
rect 466 4533 476 4536
rect 522 4533 532 4536
rect 570 4533 588 4536
rect 620 4533 637 4536
rect 682 4533 724 4536
rect 778 4533 804 4536
rect 834 4533 868 4536
rect 938 4533 972 4536
rect 1004 4533 1013 4536
rect 1156 4533 1165 4536
rect 1178 4533 1188 4536
rect 1236 4533 1253 4536
rect 1450 4533 1460 4536
rect 1772 4533 1789 4536
rect 1794 4533 1804 4536
rect 1978 4533 2004 4536
rect 2092 4533 2101 4536
rect 2106 4533 2116 4536
rect 2138 4533 2148 4536
rect 2260 4533 2388 4536
rect 202 4526 205 4533
rect 1162 4526 1165 4533
rect 2410 4526 2413 4536
rect 2506 4533 2516 4536
rect 2564 4533 2581 4536
rect 2604 4533 2621 4536
rect 2668 4533 2684 4536
rect 2706 4533 2748 4536
rect 2762 4533 2836 4536
rect 100 4523 140 4526
rect 178 4523 213 4526
rect 306 4523 332 4526
rect 444 4523 461 4526
rect 500 4523 533 4526
rect 578 4523 596 4526
rect 668 4523 725 4526
rect 996 4523 1060 4526
rect 1090 4523 1132 4526
rect 1162 4523 1196 4526
rect 1714 4523 1748 4526
rect 1780 4523 1796 4526
rect 1978 4523 1996 4526
rect 2044 4523 2061 4526
rect 2066 4523 2084 4526
rect 2140 4523 2149 4526
rect 2156 4523 2165 4526
rect 2170 4523 2236 4526
rect 2370 4523 2380 4526
rect 2410 4525 2445 4526
rect 2412 4523 2445 4525
rect 2450 4523 2524 4526
rect 2626 4523 2644 4526
rect 2708 4523 2733 4526
rect 2756 4523 2797 4526
rect 2858 4525 2861 4536
rect 2866 4533 2940 4536
rect 2962 4533 2988 4536
rect 3108 4533 3117 4536
rect 3164 4533 3197 4536
rect 3282 4533 3316 4536
rect 3346 4533 3380 4536
rect 3404 4533 3413 4536
rect 3436 4533 3460 4536
rect 3492 4533 3540 4536
rect 2874 4523 2932 4526
rect 2970 4523 2996 4526
rect 3106 4523 3116 4526
rect 3162 4523 3196 4526
rect 3228 4523 3245 4526
rect 3290 4523 3308 4526
rect 3346 4523 3349 4533
rect 3402 4523 3412 4526
rect 3514 4523 3532 4526
rect 3562 4525 3565 4536
rect 4162 4533 4172 4536
rect 4188 4533 4197 4536
rect 4226 4533 4244 4536
rect 4266 4533 4276 4536
rect 4386 4533 4420 4536
rect 4442 4533 4468 4536
rect 3570 4523 3588 4526
rect 3602 4523 3628 4526
rect 3722 4523 3772 4526
rect 3818 4523 3828 4526
rect 3956 4523 3981 4526
rect 4012 4523 4021 4526
rect 4138 4523 4156 4526
rect 4212 4523 4229 4526
rect 4274 4523 4284 4526
rect 4324 4523 4349 4526
rect 4394 4523 4412 4526
rect 4450 4523 4476 4526
rect 4482 4523 4508 4526
rect 4554 4523 4564 4526
rect 4698 4523 4708 4526
rect 4754 4523 4764 4526
rect 828 4513 861 4516
rect 14 4467 4861 4473
rect 788 4423 821 4426
rect 852 4423 884 4426
rect 220 4413 245 4416
rect 276 4413 285 4416
rect 292 4413 301 4416
rect 340 4413 365 4416
rect 396 4413 421 4416
rect 428 4413 460 4416
rect 498 4413 516 4416
rect 586 4413 620 4416
rect 650 4413 684 4416
rect 722 4413 732 4416
rect 900 4413 941 4416
rect 1004 4413 1060 4416
rect 1090 4413 1132 4416
rect 1162 4413 1236 4416
rect 1266 4413 1292 4416
rect 1322 4413 1348 4416
rect 1394 4413 1428 4416
rect 1564 4413 1581 4416
rect 1636 4413 1661 4416
rect 1756 4413 1765 4416
rect 1906 4413 1940 4416
rect 282 4405 285 4413
rect 418 4405 421 4413
rect 522 4403 540 4406
rect 578 4403 612 4406
rect 650 4403 676 4406
rect 714 4403 724 4406
rect 794 4403 828 4406
rect 852 4403 877 4406
rect 922 4403 948 4406
rect 1090 4403 1124 4406
rect 1212 4403 1221 4406
rect 1396 4403 1413 4406
rect 1708 4403 1725 4406
rect 1748 4403 1773 4406
rect 1868 4403 1893 4406
rect 1908 4403 1941 4406
rect 1970 4403 1973 4414
rect 2012 4413 2037 4416
rect 2068 4413 2077 4416
rect 2172 4413 2197 4416
rect 2234 4413 2260 4416
rect 2364 4413 2381 4416
rect 2452 4413 2477 4416
rect 2514 4413 2540 4416
rect 2716 4413 2725 4416
rect 2866 4413 2900 4416
rect 2994 4413 3020 4416
rect 3090 4413 3116 4416
rect 3162 4413 3204 4416
rect 3282 4413 3292 4416
rect 3298 4413 3332 4416
rect 3386 4413 3396 4416
rect 3426 4413 3452 4416
rect 3626 4413 3652 4416
rect 3770 4413 3796 4416
rect 3834 4413 3860 4416
rect 2074 4406 2077 4413
rect 2074 4403 2092 4406
rect 2378 4405 2381 4413
rect 3386 4406 3389 4413
rect 2682 4403 2692 4406
rect 2708 4403 2757 4406
rect 2930 4403 2948 4406
rect 3186 4403 3196 4406
rect 3228 4403 3237 4406
rect 3242 4403 3252 4406
rect 3274 4403 3284 4406
rect 3314 4403 3340 4406
rect 3356 4403 3389 4406
rect 3498 4403 3532 4406
rect 3554 4403 3580 4406
rect 3698 4403 3724 4406
rect 3834 4403 3868 4406
rect 3890 4403 3893 4414
rect 3898 4413 3932 4416
rect 3962 4403 3965 4414
rect 3978 4413 4020 4416
rect 4026 4413 4084 4416
rect 4116 4414 4133 4416
rect 4114 4413 4133 4414
rect 4138 4413 4148 4416
rect 4186 4413 4196 4416
rect 4226 4413 4252 4416
rect 4346 4413 4364 4416
rect 4394 4413 4412 4416
rect 4028 4403 4037 4406
rect 4042 4403 4092 4406
rect 4114 4403 4117 4413
rect 4186 4406 4189 4413
rect 4146 4403 4156 4406
rect 4172 4403 4189 4406
rect 4372 4403 4413 4406
rect 4442 4403 4445 4414
rect 4540 4413 4557 4416
rect 4674 4413 4700 4416
rect 4482 4403 4532 4406
rect 4546 4403 4572 4406
rect 4594 4403 4628 4406
rect 38 4367 4837 4373
rect 1114 4343 1157 4346
rect 1114 4336 1117 4343
rect 3738 4336 3741 4346
rect 4570 4336 4573 4346
rect 204 4333 221 4336
rect 322 4326 325 4335
rect 388 4333 397 4336
rect 402 4333 420 4336
rect 442 4333 460 4336
rect 602 4333 612 4336
rect 650 4333 668 4336
rect 706 4333 764 4336
rect 794 4333 828 4336
rect 858 4333 892 4336
rect 988 4333 1013 4336
rect 1108 4333 1117 4336
rect 1122 4333 1180 4336
rect 1210 4333 1284 4336
rect 1322 4333 1348 4336
rect 1748 4333 1765 4336
rect 1820 4333 1829 4336
rect 1964 4333 1989 4336
rect 2012 4333 2028 4336
rect 2154 4333 2164 4336
rect 2196 4333 2221 4336
rect 2226 4333 2244 4336
rect 2260 4333 2277 4336
rect 2316 4333 2373 4336
rect 394 4326 397 4333
rect 442 4326 445 4333
rect 2402 4326 2405 4336
rect 2522 4333 2540 4336
rect 2668 4333 2677 4336
rect 2682 4333 2692 4336
rect 2714 4333 2732 4336
rect 2804 4333 2821 4336
rect 2866 4333 2876 4336
rect 2898 4333 2924 4336
rect 3186 4326 3189 4335
rect 3474 4333 3508 4336
rect 3530 4333 3540 4336
rect 3658 4333 3692 4336
rect 3708 4333 3764 4336
rect 3946 4333 3988 4336
rect 4018 4333 4036 4336
rect 4068 4333 4077 4336
rect 4188 4333 4245 4336
rect 4338 4333 4348 4336
rect 4380 4333 4405 4336
rect 4570 4333 4580 4336
rect 66 4323 76 4326
rect 260 4323 285 4326
rect 316 4323 325 4326
rect 332 4323 364 4326
rect 394 4323 445 4326
rect 484 4323 501 4326
rect 538 4323 564 4326
rect 890 4323 900 4326
rect 1010 4323 1028 4326
rect 1074 4323 1084 4326
rect 1114 4323 1245 4326
rect 1372 4323 1389 4326
rect 1556 4323 1613 4326
rect 1620 4323 1637 4326
rect 1676 4323 1701 4326
rect 1746 4323 1780 4326
rect 1842 4323 1860 4326
rect 1970 4323 1988 4326
rect 2026 4323 2036 4326
rect 2202 4323 2236 4326
rect 2268 4323 2285 4326
rect 2362 4323 2372 4326
rect 2402 4325 2421 4326
rect 2404 4323 2421 4325
rect 2516 4323 2525 4326
rect 2612 4323 2621 4326
rect 2900 4323 2917 4326
rect 2932 4323 2941 4326
rect 2978 4323 3004 4326
rect 3042 4323 3076 4326
rect 3108 4323 3117 4326
rect 3186 4323 3212 4326
rect 3314 4323 3332 4326
rect 3362 4323 3380 4326
rect 3410 4323 3436 4326
rect 3474 4323 3500 4326
rect 3586 4323 3612 4326
rect 3666 4323 3684 4326
rect 3738 4323 3772 4326
rect 3898 4323 3908 4326
rect 4138 4323 4164 4326
rect 4194 4323 4308 4326
rect 4338 4323 4356 4326
rect 4564 4323 4581 4326
rect 4626 4323 4652 4326
rect 4690 4323 4700 4326
rect 4746 4323 4756 4326
rect 788 4313 821 4316
rect 852 4313 869 4316
rect 916 4313 925 4316
rect 14 4267 4861 4273
rect 844 4223 869 4226
rect 916 4223 925 4226
rect 140 4213 172 4216
rect 260 4213 285 4216
rect 316 4213 341 4216
rect 348 4213 364 4216
rect 540 4213 549 4216
rect 626 4213 652 4216
rect 698 4213 724 4216
rect 818 4213 828 4216
rect 890 4213 900 4216
rect 962 4213 972 4216
rect 1010 4213 1036 4216
rect 1274 4213 1324 4216
rect 1354 4213 1372 4216
rect 1386 4213 1420 4216
rect 1426 4213 1436 4216
rect 1466 4213 1492 4216
rect 1628 4213 1653 4216
rect 1780 4213 1789 4216
rect 1828 4213 1837 4216
rect 1900 4213 1925 4216
rect 1964 4213 1973 4216
rect 1994 4213 2004 4216
rect 2026 4213 2052 4216
rect 2202 4213 2244 4216
rect 2324 4213 2349 4216
rect 2402 4213 2412 4216
rect 2564 4213 2573 4216
rect 2714 4213 2732 4216
rect 66 4203 132 4206
rect 196 4203 205 4206
rect 338 4205 341 4213
rect 388 4203 429 4206
rect 546 4205 549 4213
rect 618 4203 644 4206
rect 754 4203 772 4206
rect 802 4203 820 4206
rect 844 4203 853 4206
rect 858 4203 892 4206
rect 916 4203 925 4206
rect 1226 4203 1236 4206
rect 1268 4203 1293 4206
rect 1298 4203 1316 4206
rect 1426 4205 1429 4213
rect 1700 4203 1709 4206
rect 1730 4203 1756 4206
rect 1778 4203 1804 4206
rect 1850 4203 1876 4206
rect 1962 4203 1996 4206
rect 2010 4203 2060 4206
rect 2082 4203 2108 4206
rect 2188 4203 2213 4206
rect 2226 4203 2236 4206
rect 2468 4203 2525 4206
rect 2634 4203 2652 4206
rect 2700 4203 2733 4206
rect 2762 4203 2765 4214
rect 2810 4205 2813 4216
rect 2820 4213 2829 4216
rect 2834 4203 2837 4214
rect 2906 4213 2932 4216
rect 3060 4213 3069 4216
rect 3074 4213 3100 4216
rect 3194 4213 3204 4216
rect 3364 4213 3413 4216
rect 3500 4213 3525 4216
rect 3562 4213 3604 4216
rect 3700 4213 3725 4216
rect 3802 4213 3812 4216
rect 3844 4213 3885 4216
rect 3938 4213 3948 4216
rect 3994 4213 4004 4216
rect 4074 4213 4092 4216
rect 4098 4213 4117 4216
rect 4162 4213 4180 4216
rect 4252 4213 4277 4216
rect 4386 4213 4420 4216
rect 4546 4213 4556 4216
rect 4588 4213 4604 4216
rect 4636 4214 4700 4216
rect 4634 4213 4700 4214
rect 3938 4206 3941 4213
rect 2860 4203 2869 4206
rect 3212 4203 3245 4206
rect 3268 4203 3308 4206
rect 3330 4203 3356 4206
rect 3586 4203 3596 4206
rect 3644 4203 3653 4206
rect 3772 4203 3813 4206
rect 3874 4203 3884 4206
rect 3916 4203 3941 4206
rect 4098 4205 4101 4213
rect 4162 4203 4188 4206
rect 4324 4203 4349 4206
rect 4372 4203 4428 4206
rect 4444 4203 4492 4206
rect 4524 4203 4549 4206
rect 4580 4203 4597 4206
rect 4602 4203 4612 4206
rect 4634 4203 4637 4213
rect 38 4167 4837 4173
rect 186 4133 204 4136
rect 354 4126 357 4135
rect 370 4133 396 4136
rect 428 4133 468 4136
rect 506 4133 540 4136
rect 578 4133 612 4136
rect 650 4133 692 4136
rect 730 4133 764 4136
rect 858 4133 892 4136
rect 916 4133 925 4136
rect 1060 4133 1093 4136
rect 1098 4133 1116 4136
rect 1306 4133 1316 4136
rect 1786 4133 1812 4136
rect 1850 4133 1884 4136
rect 1916 4133 1933 4136
rect 2266 4133 2292 4136
rect 2324 4133 2372 4136
rect 1090 4126 1093 4133
rect 2266 4126 2269 4133
rect 66 4123 76 4126
rect 180 4123 212 4126
rect 292 4123 317 4126
rect 348 4123 357 4126
rect 364 4123 404 4126
rect 492 4123 541 4126
rect 650 4123 700 4126
rect 844 4123 869 4126
rect 890 4123 900 4126
rect 1018 4123 1036 4126
rect 1090 4123 1124 4126
rect 1244 4123 1277 4126
rect 1298 4123 1324 4126
rect 1394 4123 1420 4126
rect 1612 4123 1629 4126
rect 1780 4123 1805 4126
rect 2084 4123 2109 4126
rect 2140 4123 2149 4126
rect 2252 4123 2269 4126
rect 2394 4125 2397 4136
rect 2882 4133 2908 4136
rect 3020 4133 3045 4136
rect 3090 4133 3100 4136
rect 3292 4133 3309 4136
rect 3452 4133 3485 4136
rect 3508 4133 3533 4136
rect 3546 4133 3580 4136
rect 3930 4133 3956 4136
rect 4444 4133 4508 4136
rect 4540 4133 4597 4136
rect 4626 4133 4684 4136
rect 2522 4123 2532 4126
rect 2570 4123 2588 4126
rect 2684 4123 2693 4126
rect 2820 4123 2837 4126
rect 2932 4123 2981 4126
rect 3076 4123 3085 4126
rect 3124 4123 3141 4126
rect 3146 4123 3172 4126
rect 3266 4123 3284 4126
rect 3290 4123 3308 4126
rect 3380 4123 3405 4126
rect 3522 4123 3572 4126
rect 3604 4123 3645 4126
rect 3788 4123 3797 4126
rect 3914 4123 3964 4126
rect 4068 4123 4077 4126
rect 4218 4123 4244 4126
rect 4332 4123 4357 4126
rect 4388 4123 4413 4126
rect 4458 4123 4516 4126
rect 4586 4123 4596 4126
rect 788 4113 805 4116
rect 916 4113 933 4116
rect 4394 4113 4413 4116
rect 14 4067 4861 4073
rect 850 4026 853 4036
rect 242 4023 277 4026
rect 748 4023 797 4026
rect 850 4023 892 4026
rect 1636 4023 1653 4026
rect 2354 4023 2373 4026
rect 2370 4016 2373 4023
rect 3090 4023 3100 4026
rect 3130 4023 3172 4026
rect 180 4013 212 4016
rect 324 4013 349 4016
rect 420 4013 445 4016
rect 476 4013 485 4016
rect 492 4013 541 4016
rect 618 4013 628 4016
rect 658 4013 692 4016
rect 778 4013 844 4016
rect 908 4013 941 4016
rect 978 4013 1013 4016
rect 1066 4013 1092 4016
rect 1348 4013 1357 4016
rect 1364 4013 1389 4016
rect 1634 4013 1684 4016
rect 1714 4013 1732 4016
rect 186 4003 204 4006
rect 482 4005 485 4013
rect 538 4005 541 4013
rect 578 4003 620 4006
rect 716 4003 725 4006
rect 852 4003 892 4006
rect 916 4003 933 4006
rect 972 4003 1005 4006
rect 1010 4005 1013 4013
rect 1778 4006 1781 4016
rect 2106 4013 2148 4016
rect 2162 4013 2196 4016
rect 2228 4013 2237 4016
rect 2348 4013 2365 4016
rect 2370 4013 2380 4016
rect 2452 4013 2461 4016
rect 2538 4013 2564 4016
rect 2596 4013 2605 4016
rect 2666 4013 2692 4016
rect 2740 4013 2749 4016
rect 2796 4013 2821 4016
rect 2852 4013 2861 4016
rect 2938 4013 2964 4016
rect 2994 4013 3036 4016
rect 2362 4006 2365 4013
rect 1050 4003 1084 4006
rect 1692 4003 1733 4006
rect 1778 4003 1812 4006
rect 1844 4003 1941 4006
rect 2156 4003 2197 4006
rect 2362 4003 2388 4006
rect 2458 4003 2508 4006
rect 2858 4005 2861 4013
rect 3090 4006 3093 4023
rect 3202 4016 3205 4026
rect 3468 4023 3477 4026
rect 3482 4023 3516 4026
rect 3116 4013 3141 4016
rect 3202 4014 3244 4016
rect 3202 4013 3245 4014
rect 3276 4013 3293 4016
rect 3362 4013 3388 4016
rect 3660 4013 3685 4016
rect 2890 4003 2956 4006
rect 2980 4003 3021 4006
rect 3052 4003 3093 4006
rect 3124 4003 3149 4006
rect 3196 4003 3205 4006
rect 3242 4003 3245 4013
rect 3698 4006 3701 4014
rect 3732 4013 3781 4016
rect 3892 4013 3917 4016
rect 3954 4013 4020 4016
rect 4042 4013 4068 4016
rect 4114 4013 4124 4016
rect 4194 4013 4228 4016
rect 4386 4013 4412 4016
rect 4442 4013 4460 4016
rect 4474 4013 4508 4016
rect 4602 4013 4628 4016
rect 3274 4003 3316 4006
rect 3434 4003 3444 4006
rect 3468 4003 3509 4006
rect 3540 4003 3549 4006
rect 3666 4003 3701 4006
rect 3724 4003 3741 4006
rect 3804 4003 3837 4006
rect 4028 4003 4037 4006
rect 4172 4003 4213 4006
rect 4338 4003 4348 4006
rect 4380 4003 4397 4006
rect 4436 4003 4461 4006
rect 4468 4003 4485 4006
rect 4610 4003 4620 4006
rect 4036 3993 4061 3996
rect 4180 3993 4205 3996
rect 4444 3993 4453 3996
rect 4476 3993 4501 3996
rect 38 3967 4837 3973
rect 170 3926 173 3935
rect 316 3933 349 3936
rect 394 3933 404 3936
rect 418 3933 452 3936
rect 484 3933 509 3936
rect 522 3933 540 3936
rect 578 3933 612 3936
rect 730 3933 780 3936
rect 860 3933 916 3936
rect 1012 3933 1045 3936
rect 1090 3933 1124 3936
rect 1170 3933 1180 3936
rect 1234 3933 1276 3936
rect 1380 3933 1404 3936
rect 1588 3933 1621 3936
rect 1690 3933 1724 3936
rect 1740 3933 1757 3936
rect 1804 3933 1821 3936
rect 1844 3933 1861 3936
rect 1908 3933 1941 3936
rect 2012 3933 2045 3936
rect 2050 3933 2060 3936
rect 2076 3933 2108 3936
rect 108 3923 133 3926
rect 164 3923 173 3926
rect 220 3923 245 3926
rect 394 3923 412 3926
rect 476 3923 493 3926
rect 666 3923 700 3926
rect 796 3923 837 3926
rect 852 3923 877 3926
rect 932 3923 973 3926
rect 1122 3923 1132 3926
rect 1162 3923 1188 3926
rect 1394 3923 1412 3926
rect 1532 3923 1557 3926
rect 1684 3923 1701 3926
rect 1748 3923 1773 3926
rect 1930 3923 1940 3926
rect 1972 3923 1997 3926
rect 2026 3923 2052 3926
rect 2084 3923 2101 3926
rect 2106 3923 2116 3926
rect 708 3913 765 3916
rect 770 3913 780 3916
rect 810 3913 844 3916
rect 858 3913 916 3916
rect 2250 3903 2253 3956
rect 2338 3933 2356 3936
rect 2372 3933 2405 3936
rect 2450 3933 2484 3936
rect 2770 3926 2773 3935
rect 2818 3933 2828 3936
rect 2860 3933 2869 3936
rect 2874 3933 2916 3936
rect 2940 3933 2949 3936
rect 2954 3933 2988 3936
rect 3012 3933 3053 3936
rect 3084 3933 3109 3936
rect 3252 3933 3285 3936
rect 3308 3933 3364 3936
rect 3386 3933 3428 3936
rect 3618 3933 3636 3936
rect 3740 3933 3821 3936
rect 2284 3923 2293 3926
rect 2380 3923 2397 3926
rect 2410 3923 2420 3926
rect 2452 3923 2469 3926
rect 2708 3923 2733 3926
rect 2764 3923 2773 3926
rect 2780 3923 2789 3926
rect 2802 3923 2836 3926
rect 2866 3913 2869 3933
rect 3850 3926 3853 3936
rect 3858 3933 3924 3936
rect 3946 3926 3949 3936
rect 3954 3933 4004 3936
rect 4026 3933 4060 3936
rect 4194 3933 4220 3936
rect 4242 3933 4284 3936
rect 4442 3933 4476 3936
rect 4498 3933 4533 3936
rect 4442 3926 4445 3933
rect 2938 3923 2996 3926
rect 3026 3923 3068 3926
rect 3210 3923 3244 3926
rect 3436 3923 3453 3926
rect 3490 3923 3516 3926
rect 3602 3923 3628 3926
rect 3660 3923 3685 3926
rect 3738 3923 3820 3926
rect 3850 3925 3861 3926
rect 3852 3923 3861 3925
rect 3866 3923 3916 3926
rect 3946 3925 3996 3926
rect 3948 3923 3996 3925
rect 4068 3923 4117 3926
rect 4194 3923 4212 3926
rect 4282 3923 4292 3926
rect 4364 3923 4389 3926
rect 4420 3923 4445 3926
rect 4498 3925 4501 3933
rect 4506 3923 4540 3926
rect 4586 3923 4596 3926
rect 4634 3923 4684 3926
rect 4722 3923 4740 3926
rect 2940 3913 2981 3916
rect 3442 3913 3453 3916
rect 3450 3903 3453 3913
rect 14 3867 4861 3873
rect 1012 3823 1021 3826
rect 3346 3823 3420 3826
rect 178 3813 212 3816
rect 324 3813 333 3816
rect 444 3813 461 3816
rect 500 3813 525 3816
rect 570 3813 621 3816
rect 674 3813 700 3816
rect 780 3813 821 3816
rect 834 3813 844 3816
rect 916 3813 949 3816
rect 994 3813 1004 3816
rect 1074 3813 1116 3816
rect 1146 3813 1172 3816
rect 1300 3813 1325 3816
rect 1346 3813 1380 3816
rect 1426 3813 1436 3816
rect 1466 3813 1492 3816
rect 1634 3813 1652 3816
rect 1698 3813 1708 3816
rect 1852 3813 1861 3816
rect 2108 3813 2133 3816
rect 2202 3813 2220 3816
rect 2418 3813 2436 3816
rect 2762 3813 2772 3816
rect 2802 3813 2836 3816
rect 2866 3813 2900 3816
rect 2930 3813 2956 3816
rect 2978 3813 3020 3816
rect 3186 3813 3212 3816
rect 194 3803 204 3806
rect 506 3803 532 3806
rect 618 3805 621 3813
rect 658 3803 692 3806
rect 730 3803 764 3806
rect 794 3803 836 3806
rect 860 3803 908 3806
rect 922 3803 948 3806
rect 972 3803 996 3806
rect 1076 3803 1108 3806
rect 1196 3803 1205 3806
rect 1346 3803 1372 3806
rect 1426 3805 1429 3813
rect 2180 3803 2221 3806
rect 2244 3803 2261 3806
rect 2538 3803 2548 3806
rect 2588 3803 2597 3806
rect 2796 3803 2804 3806
rect 2874 3803 2892 3806
rect 2964 3803 2997 3806
rect 3044 3803 3077 3806
rect 3194 3803 3204 3806
rect 3228 3803 3245 3806
rect 3250 3803 3253 3814
rect 3290 3813 3332 3816
rect 3466 3813 3484 3816
rect 3516 3813 3525 3816
rect 3596 3813 3605 3816
rect 3658 3813 3708 3816
rect 3740 3813 3757 3816
rect 3842 3813 3868 3816
rect 3914 3813 3932 3816
rect 3962 3813 3996 3816
rect 4042 3813 4052 3816
rect 4108 3813 4149 3816
rect 4170 3813 4276 3816
rect 4290 3813 4316 3816
rect 4330 3813 4364 3816
rect 4522 3813 4540 3816
rect 4594 3813 4604 3816
rect 4650 3813 4668 3816
rect 3962 3806 3965 3813
rect 3482 3803 3492 3806
rect 3514 3803 3548 3806
rect 3746 3803 3796 3806
rect 3956 3803 3965 3806
rect 4090 3803 4100 3806
rect 4138 3803 4164 3806
rect 4514 3803 4532 3806
rect 4642 3803 4676 3806
rect 2404 3793 2429 3796
rect 4172 3793 4221 3796
rect 4292 3793 4309 3796
rect 4332 3793 4341 3796
rect 38 3767 4837 3773
rect 2332 3743 2341 3746
rect 2628 3743 2637 3746
rect 3148 3743 3181 3746
rect 82 3733 148 3736
rect 244 3733 252 3736
rect 290 3733 316 3736
rect 372 3733 381 3736
rect 514 3726 517 3735
rect 570 3733 604 3736
rect 716 3733 764 3736
rect 802 3733 836 3736
rect 860 3733 892 3736
rect 906 3733 948 3736
rect 972 3733 1004 3736
rect 1084 3733 1124 3736
rect 1186 3726 1189 3735
rect 1402 3726 1405 3735
rect 1546 3733 1572 3736
rect 1586 3733 1596 3736
rect 1602 3733 1612 3736
rect 1780 3733 1829 3736
rect 1858 3733 1885 3736
rect 1914 3733 1964 3736
rect 1994 3733 2028 3736
rect 2034 3733 2068 3736
rect 2114 3733 2124 3736
rect 2178 3733 2204 3736
rect 2210 3733 2244 3736
rect 2274 3733 2324 3736
rect 2330 3733 2356 3736
rect 2380 3733 2405 3736
rect 2410 3733 2420 3736
rect 2444 3733 2453 3736
rect 2562 3733 2580 3736
rect 2986 3733 3004 3736
rect 3028 3733 3061 3736
rect 3106 3733 3140 3736
rect 3404 3733 3461 3736
rect 3468 3733 3501 3736
rect 3668 3733 3717 3736
rect 3740 3733 3757 3736
rect 3898 3733 3932 3736
rect 3954 3733 3988 3736
rect 4002 3733 4060 3736
rect 156 3723 204 3726
rect 242 3723 260 3726
rect 354 3723 364 3726
rect 444 3723 469 3726
rect 500 3723 517 3726
rect 524 3723 540 3726
rect 628 3723 692 3726
rect 834 3723 844 3726
rect 900 3723 917 3726
rect 1012 3723 1045 3726
rect 1082 3723 1132 3726
rect 1162 3723 1180 3726
rect 1186 3723 1220 3726
rect 1250 3723 1276 3726
rect 1314 3723 1356 3726
rect 1386 3723 1396 3726
rect 1402 3723 1436 3726
rect 1466 3723 1492 3726
rect 1604 3723 1613 3726
rect 1628 3723 1637 3726
rect 1802 3723 1828 3726
rect 1858 3725 1861 3733
rect 1916 3723 1925 3726
rect 2034 3725 2037 3733
rect 2562 3726 2565 3733
rect 2084 3723 2109 3726
rect 2372 3723 2421 3726
rect 2500 3723 2525 3726
rect 2556 3723 2565 3726
rect 2828 3723 2837 3726
rect 2980 3723 2997 3726
rect 3026 3723 3045 3726
rect 3084 3723 3093 3726
rect 3098 3723 3132 3726
rect 3146 3723 3188 3726
rect 3410 3723 3460 3726
rect 3474 3723 3516 3726
rect 3554 3723 3572 3726
rect 3642 3723 3652 3726
rect 3666 3723 3716 3726
rect 3762 3723 3804 3726
rect 3834 3723 3860 3726
rect 3898 3723 3924 3726
rect 3996 3723 4045 3726
rect 4082 3725 4085 3736
rect 4140 3733 4165 3736
rect 4274 3733 4309 3736
rect 4324 3733 4349 3736
rect 4362 3733 4380 3736
rect 4090 3723 4132 3726
rect 4154 3723 4172 3726
rect 4202 3723 4228 3726
rect 4274 3723 4316 3726
rect 4330 3723 4372 3726
rect 4402 3725 4405 3736
rect 4410 3733 4436 3736
rect 4530 3733 4556 3736
rect 4578 3733 4588 3736
rect 4658 3733 4676 3736
rect 4698 3733 4732 3736
rect 4746 3733 4764 3736
rect 4418 3723 4444 3726
rect 4474 3723 4500 3726
rect 4530 3723 4548 3726
rect 4580 3723 4589 3726
rect 4618 3723 4668 3726
rect 4740 3723 4749 3726
rect 4762 3723 4772 3726
rect 1020 3713 1029 3716
rect 2050 3713 2068 3716
rect 2098 3713 2124 3716
rect 2234 3713 2244 3716
rect 2346 3713 2356 3716
rect 2410 3713 2420 3716
rect 3026 3715 3029 3723
rect 3034 3713 3068 3716
rect 3282 3713 3380 3716
rect 14 3667 4861 3673
rect 748 3623 772 3626
rect 852 3623 869 3626
rect 1636 3623 1661 3626
rect 1746 3623 1764 3626
rect 1850 3623 1868 3626
rect 2042 3623 2076 3626
rect 2218 3623 2236 3626
rect 2490 3623 2516 3626
rect 2562 3623 2596 3626
rect 2842 3623 2893 3626
rect 2956 3623 2965 3626
rect 3106 3623 3116 3626
rect 3722 3623 3757 3626
rect 2890 3616 2893 3623
rect 108 3613 133 3616
rect 164 3613 173 3616
rect 180 3613 205 3616
rect 212 3613 229 3616
rect 268 3613 293 3616
rect 324 3613 333 3616
rect 340 3613 381 3616
rect 420 3613 445 3616
rect 476 3613 509 3616
rect 514 3613 532 3616
rect 722 3613 740 3616
rect 762 3613 780 3616
rect 844 3613 853 3616
rect 908 3613 957 3616
rect 962 3613 972 3616
rect 986 3613 1012 3616
rect 1058 3613 1084 3616
rect 1122 3613 1164 3616
rect 1194 3613 1244 3616
rect 1386 3613 1396 3616
rect 1426 3613 1468 3616
rect 1474 3613 1492 3616
rect 1522 3613 1548 3616
rect 170 3605 173 3613
rect 330 3605 333 3613
rect 498 3603 524 3606
rect 634 3603 660 3606
rect 698 3603 732 3606
rect 788 3603 797 3606
rect 858 3603 892 3606
rect 916 3603 925 3606
rect 1042 3603 1076 3606
rect 1188 3603 1229 3606
rect 1348 3603 1388 3606
rect 1474 3605 1477 3613
rect 1738 3606 1741 3614
rect 1780 3613 1821 3616
rect 1890 3613 1916 3616
rect 1586 3603 1612 3606
rect 1698 3603 1732 3606
rect 1738 3603 1764 3606
rect 1802 3603 1836 3606
rect 1842 3603 1868 3606
rect 1890 3605 1893 3613
rect 2034 3606 2037 3614
rect 2092 3613 2109 3616
rect 2114 3613 2132 3616
rect 2252 3613 2261 3616
rect 2290 3613 2324 3616
rect 2354 3613 2404 3616
rect 2538 3613 2548 3616
rect 2626 3613 2645 3616
rect 2650 3613 2684 3616
rect 2722 3613 2869 3616
rect 2890 3613 2933 3616
rect 2626 3606 2629 3613
rect 2018 3603 2028 3606
rect 2034 3603 2076 3606
rect 2100 3603 2133 3606
rect 2146 3603 2204 3606
rect 2210 3603 2236 3606
rect 2260 3603 2309 3606
rect 2340 3603 2381 3606
rect 2420 3603 2461 3606
rect 2482 3603 2516 3606
rect 2556 3603 2581 3606
rect 2586 3603 2596 3606
rect 2620 3603 2629 3606
rect 2634 3603 2676 3606
rect 2714 3603 2740 3606
rect 2882 3603 2908 3606
rect 2930 3605 2933 3613
rect 2954 3613 2973 3616
rect 2994 3613 3004 3616
rect 3050 3613 3060 3616
rect 2954 3605 2957 3613
rect 3106 3606 3109 3623
rect 3236 3613 3245 3616
rect 3266 3613 3276 3616
rect 3314 3613 3348 3616
rect 3362 3613 3388 3616
rect 2962 3603 2996 3606
rect 3020 3603 3037 3606
rect 3042 3603 3052 3606
rect 3076 3603 3109 3606
rect 3140 3603 3149 3606
rect 3180 3603 3197 3606
rect 3244 3603 3277 3606
rect 3300 3603 3341 3606
rect 3356 3603 3389 3606
rect 3418 3603 3421 3614
rect 3426 3613 3517 3616
rect 3618 3613 3644 3616
rect 3722 3606 3725 3623
rect 3668 3603 3725 3606
rect 3730 3606 3733 3616
rect 3796 3613 3821 3616
rect 3860 3613 3869 3616
rect 3946 3613 3972 3616
rect 4068 3613 4093 3616
rect 4124 3613 4165 3616
rect 4244 3613 4253 3616
rect 4300 3613 4317 3616
rect 4370 3613 4436 3616
rect 4506 3613 4540 3616
rect 4570 3613 4596 3616
rect 4668 3613 4685 3616
rect 4746 3613 4764 3616
rect 4314 3606 4317 3613
rect 4506 3606 4509 3613
rect 3730 3603 3788 3606
rect 3810 3603 3836 3606
rect 3852 3603 3861 3606
rect 3890 3603 3900 3606
rect 4130 3603 4180 3606
rect 4314 3603 4340 3606
rect 4442 3603 4468 3606
rect 4484 3603 4509 3606
rect 4634 3603 4644 3606
rect 4674 3603 4692 3606
rect 1706 3593 1724 3596
rect 2010 3593 2020 3596
rect 2148 3593 2189 3596
rect 2212 3593 2229 3596
rect 2484 3593 2501 3596
rect 3162 3593 3172 3596
rect 38 3567 4837 3573
rect 330 3533 372 3536
rect 426 3533 468 3536
rect 506 3533 540 3536
rect 586 3526 589 3535
rect 748 3533 765 3536
rect 770 3533 788 3536
rect 818 3533 876 3536
rect 900 3533 916 3536
rect 1018 3533 1052 3536
rect 1362 3533 1380 3536
rect 1594 3533 1612 3536
rect 1642 3533 1660 3536
rect 1684 3533 1693 3536
rect 1714 3533 1724 3536
rect 1794 3533 1804 3536
rect 1828 3533 1861 3536
rect 1900 3533 1933 3536
rect 1972 3533 2021 3536
rect 2052 3533 2085 3536
rect 2090 3533 2100 3536
rect 2124 3533 2165 3536
rect 2196 3533 2237 3536
rect 2242 3533 2252 3536
rect 2276 3533 2309 3536
rect 2314 3533 2324 3536
rect 2348 3533 2381 3536
rect 2404 3533 2437 3536
rect 2242 3526 2245 3533
rect 2314 3526 2317 3533
rect 2770 3526 2773 3535
rect 2786 3533 2820 3536
rect 2852 3533 2877 3536
rect 3010 3533 3052 3536
rect 3076 3533 3085 3536
rect 3090 3533 3116 3536
rect 3140 3533 3181 3536
rect 3210 3526 3213 3535
rect 3354 3533 3364 3536
rect 3434 3533 3444 3536
rect 3458 3533 3500 3536
rect 3516 3533 3572 3536
rect 3588 3533 3644 3536
rect 3668 3533 3709 3536
rect 3748 3533 3781 3536
rect 108 3523 133 3526
rect 260 3523 285 3526
rect 316 3523 325 3526
rect 338 3523 380 3526
rect 492 3523 589 3526
rect 706 3523 740 3526
rect 804 3523 869 3526
rect 1308 3523 1333 3526
rect 1340 3523 1357 3526
rect 1442 3523 1452 3526
rect 1482 3523 1508 3526
rect 1580 3523 1589 3526
rect 1676 3523 1732 3526
rect 1826 3523 1884 3526
rect 1906 3523 1956 3526
rect 1978 3523 2036 3526
rect 2058 3523 2108 3526
rect 2138 3523 2180 3526
rect 2194 3523 2245 3526
rect 2250 3523 2260 3526
rect 2282 3523 2317 3526
rect 2354 3523 2396 3526
rect 2476 3523 2501 3526
rect 2532 3523 2541 3526
rect 2700 3523 2725 3526
rect 2756 3523 2773 3526
rect 2818 3523 2828 3526
rect 2930 3523 2956 3526
rect 3050 3523 3060 3526
rect 3074 3523 3124 3526
rect 3210 3523 3244 3526
rect 3372 3523 3381 3526
rect 3452 3523 3485 3526
rect 3524 3523 3549 3526
rect 3596 3523 3621 3526
rect 3642 3523 3652 3526
rect 3674 3523 3724 3526
rect 3786 3525 3789 3536
rect 3818 3525 3821 3536
rect 3930 3533 3948 3536
rect 3964 3533 4005 3536
rect 4114 3533 4164 3536
rect 4186 3533 4244 3536
rect 4274 3533 4292 3536
rect 4410 3533 4460 3536
rect 4530 3533 4564 3536
rect 4002 3526 4005 3533
rect 3826 3523 3860 3526
rect 3874 3523 3940 3526
rect 4002 3523 4020 3526
rect 4066 3523 4076 3526
rect 4114 3523 4156 3526
rect 4194 3523 4252 3526
rect 4258 3523 4284 3526
rect 4298 3523 4372 3526
rect 4404 3523 4437 3526
rect 4450 3523 4468 3526
rect 4594 3525 4597 3536
rect 4634 3533 4660 3536
rect 4628 3523 4652 3526
rect 4682 3525 4685 3536
rect 4746 3523 4764 3526
rect 650 3513 732 3516
rect 1636 3513 1660 3516
rect 1786 3513 1804 3516
rect 2124 3513 2133 3516
rect 2196 3513 2205 3516
rect 3076 3513 3101 3516
rect 3146 3513 3188 3516
rect 4114 3513 4117 3523
rect 4410 3513 4413 3523
rect 14 3467 4861 3473
rect 650 3423 676 3426
rect 788 3423 805 3426
rect 826 3423 836 3426
rect 898 3423 908 3426
rect 3020 3423 3077 3426
rect 3346 3423 3396 3426
rect 140 3413 172 3416
rect 252 3413 277 3416
rect 308 3413 317 3416
rect 332 3413 341 3416
rect 354 3413 372 3416
rect 402 3413 428 3416
rect 554 3413 620 3416
rect 786 3413 805 3416
rect 818 3413 844 3416
rect 924 3413 1069 3416
rect 1082 3413 1188 3416
rect 1218 3413 1228 3416
rect 1258 3413 1284 3416
rect 1410 3413 1436 3416
rect 1450 3413 1468 3416
rect 1548 3413 1573 3416
rect 1954 3413 2005 3416
rect 2036 3413 2077 3416
rect 2172 3413 2197 3416
rect 2228 3413 2245 3416
rect 2252 3413 2293 3416
rect 2516 3413 2533 3416
rect 2556 3413 2613 3416
rect 2650 3413 2716 3416
rect 2796 3413 2821 3416
rect 2866 3413 2916 3416
rect 2922 3413 2948 3416
rect 2994 3413 3004 3416
rect 3034 3413 3100 3416
rect 3114 3413 3148 3416
rect 3242 3413 3252 3416
rect 3298 3413 3308 3416
rect 3340 3413 3365 3416
rect 3418 3413 3460 3416
rect 3490 3413 3516 3416
rect 3580 3413 3589 3416
rect 3634 3413 3660 3416
rect 3834 3413 3884 3416
rect 3890 3413 3940 3416
rect 3986 3413 4028 3416
rect 4132 3413 4157 3416
rect 4298 3413 4324 3416
rect 4362 3413 4388 3416
rect 4394 3413 4404 3416
rect 4450 3413 4460 3416
rect 4554 3413 4613 3416
rect 4682 3413 4692 3416
rect 4698 3413 4708 3416
rect 4754 3413 4764 3416
rect 402 3406 405 3413
rect 196 3403 213 3406
rect 396 3403 413 3406
rect 586 3403 612 3406
rect 692 3403 701 3406
rect 852 3403 908 3406
rect 1026 3403 1069 3406
rect 1140 3403 1173 3406
rect 1212 3403 1221 3406
rect 1332 3403 1341 3406
rect 1346 3403 1388 3406
rect 1642 3403 1652 3406
rect 1684 3403 1709 3406
rect 1748 3403 1781 3406
rect 1794 3403 1804 3406
rect 2002 3403 2012 3406
rect 2058 3403 2100 3406
rect 2242 3405 2245 3413
rect 2274 3403 2292 3406
rect 2324 3403 2341 3406
rect 2538 3403 2548 3406
rect 2562 3403 2612 3406
rect 2658 3403 2708 3406
rect 2778 3403 2788 3406
rect 2810 3403 2828 3406
rect 2860 3403 2877 3406
rect 2898 3403 2908 3406
rect 2956 3403 2965 3406
rect 2970 3403 2996 3406
rect 3020 3403 3085 3406
rect 3116 3403 3141 3406
rect 3260 3403 3309 3406
rect 3418 3405 3421 3413
rect 3802 3403 3876 3406
rect 3930 3403 3948 3406
rect 3978 3403 4020 3406
rect 4034 3403 4060 3406
rect 4202 3403 4228 3406
rect 4298 3403 4316 3406
rect 4354 3403 4380 3406
rect 4540 3403 4677 3406
rect 38 3367 4837 3373
rect 3740 3343 3749 3346
rect 194 3333 244 3336
rect 314 3333 324 3336
rect 410 3333 420 3336
rect 492 3333 533 3336
rect 538 3333 548 3336
rect 586 3333 620 3336
rect 658 3333 700 3336
rect 738 3333 780 3336
rect 804 3333 844 3336
rect 924 3333 972 3336
rect 1076 3333 1117 3336
rect 1162 3333 1196 3336
rect 538 3326 541 3333
rect 1218 3326 1221 3336
rect 1242 3333 1276 3336
rect 1308 3333 1333 3336
rect 1554 3333 1580 3336
rect 1602 3333 1612 3336
rect 1740 3333 1749 3336
rect 1786 3333 1796 3336
rect 1820 3333 1845 3336
rect 1850 3333 1876 3336
rect 1996 3333 2005 3336
rect 2236 3333 2253 3336
rect 2284 3333 2293 3336
rect 2354 3333 2364 3336
rect 2538 3333 2572 3336
rect 2604 3333 2645 3336
rect 2770 3333 2804 3336
rect 2850 3333 2876 3336
rect 3066 3333 3132 3336
rect 3154 3326 3157 3334
rect 3236 3333 3261 3336
rect 3282 3333 3316 3336
rect 3506 3333 3548 3336
rect 3690 3333 3732 3336
rect 116 3323 141 3326
rect 210 3323 252 3326
rect 332 3323 357 3326
rect 444 3323 549 3326
rect 618 3323 628 3326
rect 658 3323 708 3326
rect 810 3323 852 3326
rect 866 3323 916 3326
rect 988 3323 1037 3326
rect 1082 3323 1132 3326
rect 1218 3323 1236 3326
rect 1266 3323 1284 3326
rect 1338 3323 1348 3326
rect 1378 3323 1404 3326
rect 1588 3323 1613 3326
rect 1650 3323 1684 3326
rect 1714 3323 1732 3326
rect 1812 3323 1829 3326
rect 1874 3323 1884 3326
rect 1946 3323 1972 3326
rect 2002 3323 2053 3326
rect 2058 3323 2068 3326
rect 2098 3323 2124 3326
rect 2162 3323 2212 3326
rect 2242 3323 2285 3326
rect 2306 3323 2372 3326
rect 2476 3323 2501 3326
rect 2708 3323 2733 3326
rect 2764 3323 2781 3326
rect 2842 3323 2884 3326
rect 2962 3323 2972 3326
rect 3010 3323 3028 3326
rect 3090 3323 3140 3326
rect 3154 3323 3165 3326
rect 3228 3323 3253 3326
rect 3276 3323 3301 3326
rect 3340 3323 3381 3326
rect 3386 3323 3396 3326
rect 3426 3323 3452 3326
rect 3572 3323 3605 3326
rect 3618 3323 3628 3326
rect 3674 3323 3724 3326
rect 3786 3325 3789 3336
rect 4106 3333 4132 3336
rect 4282 3333 4300 3336
rect 4282 3326 4285 3333
rect 4042 3323 4076 3326
rect 4108 3323 4133 3326
rect 4140 3323 4149 3326
rect 4196 3323 4213 3326
rect 4252 3323 4285 3326
rect 4322 3325 4325 3336
rect 4402 3333 4420 3336
rect 4482 3333 4500 3336
rect 4522 3333 4548 3336
rect 4706 3333 4740 3336
rect 4380 3323 4397 3326
rect 4444 3323 4492 3326
rect 4524 3323 4549 3326
rect 4708 3323 4717 3326
rect 4748 3323 4757 3326
rect 3162 3316 3165 3323
rect 196 3313 221 3316
rect 938 3313 972 3316
rect 1754 3313 1796 3316
rect 3162 3313 3212 3316
rect 14 3267 4861 3273
rect 4434 3233 4453 3236
rect 204 3223 221 3226
rect 292 3223 317 3226
rect 380 3223 389 3226
rect 420 3223 429 3226
rect 556 3223 573 3226
rect 890 3223 908 3226
rect 938 3223 972 3226
rect 2356 3223 2389 3226
rect 2452 3223 2461 3226
rect 2498 3223 2524 3226
rect 2978 3223 3012 3226
rect 3138 3223 3196 3226
rect 3586 3223 3636 3226
rect 2978 3216 2981 3223
rect 4698 3216 4701 3226
rect 108 3213 117 3216
rect 164 3213 173 3216
rect 196 3213 269 3216
rect 324 3213 364 3216
rect 418 3213 540 3216
rect 554 3213 605 3216
rect 650 3213 692 3216
rect 706 3213 756 3216
rect 820 3213 845 3216
rect 852 3213 869 3216
rect 890 3213 916 3216
rect 988 3213 1045 3216
rect 1082 3213 1140 3216
rect 1170 3213 1204 3216
rect 1218 3213 1244 3216
rect 1282 3213 1324 3216
rect 1524 3213 1533 3216
rect 1588 3213 1613 3216
rect 1778 3213 1804 3216
rect 1898 3213 1908 3216
rect 2050 3213 2092 3216
rect 2146 3213 2156 3216
rect 2354 3213 2396 3216
rect 2402 3213 2444 3216
rect 2492 3213 2525 3216
rect 2540 3213 2589 3216
rect 2594 3213 2629 3216
rect 2668 3213 2693 3216
rect 2724 3213 2733 3216
rect 2812 3213 2821 3216
rect 2868 3213 2909 3216
rect 2916 3213 2949 3216
rect 290 3203 316 3206
rect 338 3203 356 3206
rect 420 3203 445 3206
rect 450 3203 460 3206
rect 482 3203 532 3206
rect 554 3205 557 3213
rect 562 3203 612 3206
rect 700 3203 741 3206
rect 762 3203 804 3206
rect 860 3203 909 3206
rect 924 3203 972 3206
rect 1076 3203 1093 3206
rect 1122 3203 1132 3206
rect 1164 3203 1197 3206
rect 1212 3203 1221 3206
rect 1338 3203 1364 3206
rect 1644 3203 1684 3206
rect 2306 3203 2332 3206
rect 2356 3203 2389 3206
rect 2404 3203 2436 3206
rect 2450 3203 2484 3206
rect 2522 3205 2525 3213
rect 2548 3203 2557 3206
rect 2730 3205 2733 3213
rect 2906 3205 2909 3213
rect 2946 3205 2949 3213
rect 2970 3213 2981 3216
rect 3090 3213 3116 3216
rect 3178 3213 3197 3216
rect 3212 3213 3245 3216
rect 3322 3213 3348 3216
rect 3444 3213 3453 3216
rect 3458 3213 3468 3216
rect 3490 3213 3516 3216
rect 3546 3213 3564 3216
rect 3714 3213 3732 3216
rect 3786 3213 3796 3216
rect 3834 3213 3852 3216
rect 3978 3213 4036 3216
rect 4050 3213 4092 3216
rect 4186 3213 4228 3216
rect 4674 3213 4708 3216
rect 4754 3213 4764 3216
rect 2970 3205 2973 3213
rect 3036 3203 3053 3206
rect 3058 3203 3068 3206
rect 3074 3203 3108 3206
rect 3132 3203 3189 3206
rect 3194 3205 3197 3213
rect 3786 3206 3789 3213
rect 3220 3203 3261 3206
rect 3266 3203 3276 3206
rect 3532 3203 3541 3206
rect 3572 3203 3589 3206
rect 3618 3203 3636 3206
rect 3660 3203 3685 3206
rect 3706 3203 3724 3206
rect 3756 3203 3789 3206
rect 3930 3203 3940 3206
rect 3972 3203 4029 3206
rect 4034 3203 4044 3206
rect 4226 3203 4236 3206
rect 4516 3203 4549 3206
rect 3042 3193 3060 3196
rect 4052 3193 4061 3196
rect 38 3167 4837 3173
rect 650 3143 677 3146
rect 3962 3143 3997 3146
rect 4234 3143 4245 3146
rect 650 3136 653 3143
rect 178 3126 181 3134
rect 268 3133 301 3136
rect 340 3133 349 3136
rect 466 3133 476 3136
rect 508 3133 541 3136
rect 628 3133 653 3136
rect 658 3133 684 3136
rect 708 3133 741 3136
rect 922 3133 932 3136
rect 1012 3133 1037 3136
rect 1042 3133 1052 3136
rect 1084 3133 1093 3136
rect 1418 3133 1444 3136
rect 1738 3126 1741 3134
rect 1828 3133 1876 3136
rect 1914 3133 1940 3136
rect 2332 3133 2389 3136
rect 2538 3126 2541 3134
rect 2554 3133 2604 3136
rect 2642 3133 2708 3136
rect 2754 3133 2804 3136
rect 2962 3126 2965 3134
rect 3034 3126 3037 3134
rect 3164 3133 3181 3136
rect 3186 3133 3276 3136
rect 3396 3133 3405 3136
rect 3450 3133 3500 3136
rect 3634 3133 3660 3136
rect 3778 3133 3804 3136
rect 3852 3133 3861 3136
rect 3884 3133 3917 3136
rect 3962 3133 4012 3136
rect 4028 3133 4116 3136
rect 4170 3133 4196 3136
rect 4212 3133 4237 3136
rect 3914 3126 3917 3133
rect 4242 3126 4245 3143
rect 4324 3133 4349 3136
rect 108 3123 133 3126
rect 164 3123 181 3126
rect 188 3123 197 3126
rect 218 3123 228 3126
rect 260 3123 285 3126
rect 332 3123 364 3126
rect 458 3123 484 3126
rect 490 3123 500 3126
rect 548 3123 612 3126
rect 650 3123 692 3126
rect 722 3123 748 3126
rect 810 3123 820 3126
rect 978 3123 988 3126
rect 1026 3123 1060 3126
rect 1276 3123 1285 3126
rect 218 3116 221 3123
rect 196 3113 221 3116
rect 274 3113 300 3116
rect 514 3113 540 3116
rect 628 3113 637 3116
rect 708 3113 733 3116
rect 1364 3113 1373 3116
rect 1378 3113 1388 3116
rect 1402 3106 1405 3125
rect 1460 3123 1469 3126
rect 1492 3123 1501 3126
rect 1548 3123 1573 3126
rect 1652 3123 1677 3126
rect 1708 3123 1741 3126
rect 1754 3123 1804 3126
rect 1900 3123 1988 3126
rect 2074 3123 2092 3126
rect 2130 3123 2189 3126
rect 2194 3123 2228 3126
rect 2258 3123 2316 3126
rect 2452 3123 2477 3126
rect 2508 3123 2541 3126
rect 2548 3123 2565 3126
rect 2578 3123 2612 3126
rect 2650 3123 2716 3126
rect 2746 3123 2812 3126
rect 2962 3123 3037 3126
rect 3044 3123 3093 3126
rect 3098 3123 3140 3126
rect 3172 3123 3189 3126
rect 3210 3123 3268 3126
rect 3314 3123 3380 3126
rect 3436 3123 3461 3126
rect 3466 3123 3492 3126
rect 3620 3123 3653 3126
rect 3668 3123 3677 3126
rect 3714 3123 3740 3126
rect 3818 3123 3844 3126
rect 3914 3123 3940 3126
rect 4124 3123 4133 3126
rect 4138 3123 4188 3126
rect 4220 3123 4229 3126
rect 4242 3123 4300 3126
rect 4388 3123 4397 3126
rect 4450 3123 4460 3126
rect 4506 3123 4516 3126
rect 4596 3123 4621 3126
rect 4730 3123 4748 3126
rect 2930 3113 2948 3116
rect 3530 3113 3604 3116
rect 1402 3103 1437 3106
rect 14 3067 4861 3073
rect 1274 3033 1325 3036
rect 2314 3033 2349 3036
rect 490 3023 508 3026
rect 522 3023 548 3026
rect 642 3016 645 3026
rect 1122 3023 1133 3026
rect 1130 3016 1133 3023
rect 146 3013 188 3016
rect 218 3013 244 3016
rect 308 3013 317 3016
rect 516 3013 541 3016
rect 556 3013 620 3016
rect 634 3013 645 3016
rect 762 3013 836 3016
rect 866 3013 876 3016
rect 906 3013 956 3016
rect 1036 3013 1069 3016
rect 634 3007 637 3013
rect 906 3006 909 3013
rect 1066 3007 1069 3013
rect 1090 3013 1100 3016
rect 1130 3013 1156 3016
rect 1228 3013 1237 3016
rect 1274 3015 1277 3033
rect 1284 3023 1293 3026
rect 1386 3023 1412 3026
rect 2884 3023 2933 3026
rect 3564 3023 3573 3026
rect 4746 3023 4765 3026
rect 4746 3016 4749 3023
rect 1364 3013 1405 3016
rect 1442 3013 1492 3016
rect 1596 3013 1621 3016
rect 1652 3013 1661 3016
rect 1724 3013 1749 3016
rect 1876 3013 1885 3016
rect 1892 3013 1901 3016
rect 1956 3013 1973 3016
rect 2012 3013 2029 3016
rect 2164 3013 2173 3016
rect 1090 3007 1093 3013
rect 1658 3007 1661 3013
rect 1882 3007 1885 3013
rect 2026 3007 2029 3013
rect 300 3003 325 3006
rect 330 3003 340 3006
rect 468 3003 509 3006
rect 860 3003 869 3006
rect 900 3003 909 3006
rect 970 3003 1012 3006
rect 1170 3003 1204 3006
rect 1322 3003 1340 3006
rect 1356 3003 1405 3006
rect 1442 3003 1500 3006
rect 1516 3003 1557 3006
rect 2354 3005 2357 3016
rect 2380 3013 2397 3016
rect 2402 3013 2452 3016
rect 2548 3013 2557 3016
rect 2604 3013 2621 3016
rect 2780 3013 2789 3016
rect 2794 3013 2804 3016
rect 2394 3006 2397 3013
rect 2394 3003 2445 3006
rect 2476 3003 2493 3006
rect 2618 3005 2621 3013
rect 2810 3005 2813 3016
rect 2882 3013 2949 3016
rect 3084 3013 3093 3016
rect 3140 3013 3237 3016
rect 3282 3013 3316 3016
rect 3338 3013 3356 3016
rect 3452 3013 3461 3016
rect 3508 3013 3541 3016
rect 3578 3013 3684 3016
rect 3722 3013 3764 3016
rect 3810 3013 3820 3016
rect 3916 3013 3940 3016
rect 4172 3013 4181 3016
rect 4186 3013 4204 3016
rect 4242 3013 4268 3016
rect 4290 3013 4316 3016
rect 2818 3003 2860 3006
rect 2882 3005 2885 3013
rect 2898 3003 2948 3006
rect 2972 3003 3045 3006
rect 3234 3005 3237 3013
rect 3260 3003 3301 3006
rect 3538 3005 3541 3013
rect 3564 3003 3597 3006
rect 3612 3003 3621 3006
rect 3626 3003 3692 3006
rect 3874 3003 3900 3006
rect 3956 3003 4077 3006
rect 4276 3003 4301 3006
rect 4306 3003 4324 3006
rect 4378 3003 4381 3014
rect 4412 3013 4421 3016
rect 4554 3013 4572 3016
rect 4682 3013 4700 3016
rect 4732 3013 4749 3016
rect 4754 3013 4780 3016
rect 4410 3003 4500 3006
rect 4596 3003 4605 3006
rect 4610 3003 4636 3006
rect 4658 3003 4708 3006
rect 4730 3003 4772 3006
rect 282 2993 292 2996
rect 4220 2993 4261 2996
rect 4284 2993 4317 2996
rect 4332 2993 4341 2996
rect 38 2967 4837 2973
rect 3394 2953 3421 2956
rect 1778 2936 1781 2946
rect 2898 2943 2917 2946
rect 2898 2936 2901 2943
rect 204 2933 221 2936
rect 290 2933 324 2936
rect 356 2933 397 2936
rect 588 2933 597 2936
rect 858 2933 900 2936
rect 1044 2933 1085 2936
rect 1452 2933 1477 2936
rect 1482 2933 1500 2936
rect 1516 2933 1549 2936
rect 1588 2933 1621 2936
rect 1642 2933 1676 2936
rect 1714 2933 1732 2936
rect 1778 2933 1804 2936
rect 2218 2933 2244 2936
rect 1482 2926 1485 2933
rect 108 2923 125 2926
rect 186 2923 196 2926
rect 202 2923 244 2926
rect 268 2923 317 2926
rect 322 2923 332 2926
rect 636 2923 661 2926
rect 692 2923 709 2926
rect 746 2923 772 2926
rect 930 2923 972 2926
rect 1004 2923 1029 2926
rect 1082 2923 1092 2926
rect 1410 2923 1485 2926
rect 1554 2923 1557 2933
rect 1626 2923 1629 2933
rect 2370 2926 2373 2936
rect 2506 2933 2524 2936
rect 2556 2933 2581 2936
rect 2594 2933 2604 2936
rect 2786 2933 2812 2936
rect 2834 2933 2868 2936
rect 2892 2933 2901 2936
rect 2906 2933 2924 2936
rect 2948 2933 3013 2936
rect 3140 2933 3157 2936
rect 3266 2933 3284 2936
rect 3314 2933 3364 2936
rect 3444 2933 3453 2936
rect 3618 2933 3644 2936
rect 3660 2933 3677 2936
rect 1700 2923 1740 2926
rect 1770 2923 1812 2926
rect 1868 2923 1885 2926
rect 2140 2923 2148 2926
rect 2186 2923 2196 2926
rect 2266 2923 2284 2926
rect 2370 2923 2396 2926
rect 2442 2923 2452 2926
rect 2490 2923 2532 2926
rect 2562 2923 2612 2926
rect 2642 2923 2692 2926
rect 2738 2923 2756 2926
rect 2778 2923 2820 2926
rect 2866 2923 2876 2926
rect 3036 2923 3077 2926
rect 3090 2923 3132 2926
rect 3250 2923 3276 2926
rect 3322 2923 3372 2926
rect 3378 2923 3428 2926
rect 3450 2923 3453 2933
rect 3682 2926 3685 2956
rect 3698 2933 3724 2936
rect 4212 2933 4237 2936
rect 4250 2933 4268 2936
rect 4284 2933 4293 2936
rect 4404 2933 4421 2936
rect 4418 2926 4421 2933
rect 4626 2926 4629 2936
rect 4658 2933 4692 2936
rect 3482 2923 3508 2926
rect 3554 2923 3564 2926
rect 3668 2923 3685 2926
rect 3732 2923 3749 2926
rect 3786 2923 3812 2926
rect 3858 2923 3868 2926
rect 3914 2923 3924 2926
rect 3962 2923 3972 2926
rect 4100 2923 4117 2926
rect 4220 2923 4237 2926
rect 4292 2923 4309 2926
rect 4410 2923 4452 2926
rect 4602 2925 4629 2926
rect 4602 2923 4628 2925
rect 4754 2923 4764 2926
rect 1122 2913 1172 2916
rect 1210 2913 1252 2916
rect 1276 2913 1285 2916
rect 2892 2913 2917 2916
rect 3322 2913 3325 2923
rect 4602 2913 4605 2923
rect 1180 2903 1261 2906
rect 14 2867 4861 2873
rect 580 2833 661 2836
rect 2946 2826 2949 2836
rect 522 2823 572 2826
rect 596 2823 653 2826
rect 2924 2823 2949 2826
rect 3170 2823 3204 2826
rect 3362 2823 3404 2826
rect 3594 2823 3644 2826
rect 3906 2823 3925 2826
rect 3922 2816 3925 2823
rect 298 2813 324 2816
rect 394 2813 412 2816
rect 442 2813 492 2816
rect 516 2813 565 2816
rect 690 2813 732 2816
rect 738 2813 772 2816
rect 778 2813 796 2816
rect 108 2803 157 2806
rect 284 2803 317 2806
rect 428 2803 493 2806
rect 508 2803 533 2806
rect 658 2803 676 2806
rect 740 2803 749 2806
rect 780 2803 797 2806
rect 826 2803 829 2814
rect 842 2813 852 2816
rect 906 2806 909 2816
rect 914 2813 932 2816
rect 964 2813 981 2816
rect 1092 2813 1101 2816
rect 1132 2813 1141 2816
rect 1196 2813 1221 2816
rect 1252 2813 1261 2816
rect 1268 2813 1301 2816
rect 1338 2813 1388 2816
rect 1564 2813 1573 2816
rect 1620 2813 1629 2816
rect 1730 2813 1748 2816
rect 1978 2813 1996 2816
rect 2100 2813 2109 2816
rect 2204 2813 2221 2816
rect 2298 2813 2316 2816
rect 2386 2813 2397 2816
rect 2404 2813 2421 2816
rect 2466 2813 2476 2816
rect 2538 2813 2548 2816
rect 2594 2813 2604 2816
rect 2642 2813 2692 2816
rect 2722 2813 2813 2816
rect 2898 2813 2908 2816
rect 2930 2813 2996 2816
rect 3026 2813 3052 2816
rect 3058 2813 3068 2816
rect 3098 2813 3124 2816
rect 1258 2807 1261 2813
rect 2106 2806 2109 2813
rect 2386 2807 2389 2813
rect 3058 2807 3061 2813
rect 3202 2807 3205 2816
rect 3226 2813 3268 2816
rect 3554 2813 3588 2816
rect 3666 2813 3716 2816
rect 3828 2813 3837 2816
rect 3884 2813 3917 2816
rect 3922 2813 3980 2816
rect 4012 2813 4021 2816
rect 4026 2813 4052 2816
rect 4074 2813 4124 2816
rect 4202 2813 4228 2816
rect 4298 2813 4316 2816
rect 4330 2813 4404 2816
rect 4436 2813 4477 2816
rect 4530 2813 4556 2816
rect 4666 2813 4708 2816
rect 4802 2813 4869 2816
rect 3226 2807 3229 2813
rect 4666 2806 4669 2813
rect 906 2803 940 2806
rect 962 2803 988 2806
rect 1282 2803 1300 2806
rect 1332 2803 1373 2806
rect 1658 2803 1684 2806
rect 1716 2803 1725 2806
rect 1916 2803 1925 2806
rect 1930 2803 1948 2806
rect 2004 2803 2037 2806
rect 2106 2803 2124 2806
rect 2210 2803 2228 2806
rect 2332 2803 2341 2806
rect 2410 2803 2428 2806
rect 2460 2803 2469 2806
rect 2658 2803 2684 2806
rect 2882 2803 2900 2806
rect 2924 2803 2941 2806
rect 2946 2803 2988 2806
rect 3012 2803 3045 2806
rect 3362 2803 3389 2806
rect 3394 2803 3404 2806
rect 3428 2803 3485 2806
rect 3506 2803 3580 2806
rect 3634 2803 3644 2806
rect 3668 2803 3677 2806
rect 3724 2803 3749 2806
rect 3762 2803 3797 2806
rect 3826 2803 3876 2806
rect 3890 2803 3988 2806
rect 4034 2803 4044 2806
rect 4058 2803 4132 2806
rect 4148 2803 4181 2806
rect 4186 2803 4236 2806
rect 4252 2803 4269 2806
rect 4290 2803 4324 2806
rect 4434 2803 4500 2806
rect 4580 2803 4629 2806
rect 4652 2803 4669 2806
rect 116 2793 125 2796
rect 154 2793 157 2803
rect 2938 2796 2941 2803
rect 4186 2796 4189 2803
rect 204 2793 245 2796
rect 442 2793 492 2796
rect 2938 2793 2973 2796
rect 4162 2793 4189 2796
rect 4332 2793 4397 2796
rect 38 2767 4837 2773
rect 170 2743 204 2746
rect 938 2736 941 2746
rect 1386 2743 1413 2746
rect 2090 2736 2093 2756
rect 3402 2753 3429 2756
rect 4178 2736 4181 2746
rect 212 2733 237 2736
rect 458 2733 468 2736
rect 580 2733 597 2736
rect 602 2733 612 2736
rect 724 2733 741 2736
rect 802 2733 820 2736
rect 932 2733 941 2736
rect 1314 2733 1340 2736
rect 1770 2733 1788 2736
rect 1802 2733 1852 2736
rect 1922 2733 1940 2736
rect 1956 2733 1973 2736
rect 2036 2733 2045 2736
rect 2084 2733 2093 2736
rect 2322 2733 2340 2736
rect 2378 2733 2396 2736
rect 2418 2733 2436 2736
rect 2468 2733 2493 2736
rect 2610 2733 2620 2736
rect 2852 2733 2877 2736
rect 2882 2733 2892 2736
rect 2930 2733 2988 2736
rect 3012 2733 3093 2736
rect 450 2726 453 2733
rect 1290 2726 1293 2733
rect 1730 2726 1733 2733
rect 1970 2726 1973 2733
rect 3106 2726 3109 2734
rect 3434 2733 3500 2736
rect 3516 2733 3620 2736
rect 3636 2733 3653 2736
rect 3802 2733 3836 2736
rect 3858 2733 3868 2736
rect 4114 2733 4148 2736
rect 4170 2733 4181 2736
rect 4290 2733 4316 2736
rect 4610 2733 4676 2736
rect 4698 2733 4732 2736
rect 4754 2733 4780 2736
rect 3650 2726 3653 2733
rect 4114 2726 4117 2733
rect 100 2723 133 2726
rect 130 2706 133 2723
rect 146 2706 149 2725
rect 220 2723 333 2726
rect 450 2723 461 2726
rect 716 2723 765 2726
rect 1114 2723 1157 2726
rect 1204 2723 1229 2726
rect 1260 2723 1293 2726
rect 1300 2723 1341 2726
rect 1660 2723 1685 2726
rect 1716 2723 1733 2726
rect 1740 2723 1749 2726
rect 1796 2723 1845 2726
rect 1882 2723 1932 2726
rect 1970 2723 2037 2726
rect 2082 2723 2100 2726
rect 2130 2723 2156 2726
rect 2236 2723 2253 2726
rect 2348 2723 2357 2726
rect 2404 2723 2413 2726
rect 2548 2723 2557 2726
rect 2588 2723 2621 2726
rect 2818 2723 2828 2726
rect 2866 2723 2900 2726
rect 2986 2723 2996 2726
rect 3098 2723 3109 2726
rect 3116 2723 3157 2726
rect 3202 2723 3220 2726
rect 3524 2723 3573 2726
rect 3650 2723 3692 2726
rect 3722 2723 3748 2726
rect 3786 2723 3828 2726
rect 3972 2723 3981 2726
rect 4052 2723 4061 2726
rect 4108 2723 4117 2726
rect 4170 2725 4173 2733
rect 4220 2723 4245 2726
rect 4290 2723 4324 2726
rect 4378 2723 4388 2726
rect 4426 2723 4436 2726
rect 4442 2723 4492 2726
rect 4548 2723 4557 2726
rect 4610 2723 4668 2726
rect 4700 2723 4709 2726
rect 4740 2723 4757 2726
rect 4762 2723 4788 2726
rect 164 2713 173 2716
rect 130 2703 149 2706
rect 458 2703 461 2723
rect 730 2713 772 2716
rect 796 2713 813 2716
rect 938 2713 964 2716
rect 978 2713 988 2716
rect 972 2703 1061 2706
rect 14 2667 4861 2673
rect 354 2616 357 2636
rect 410 2633 452 2636
rect 1642 2633 1661 2636
rect 1708 2633 1765 2636
rect 468 2623 493 2626
rect 604 2623 613 2626
rect 882 2623 924 2626
rect 1066 2623 1076 2626
rect 98 2613 108 2616
rect 132 2613 189 2616
rect 186 2607 189 2613
rect 346 2613 357 2616
rect 370 2613 380 2616
rect 404 2613 445 2616
rect 506 2613 524 2616
rect 548 2613 565 2616
rect 634 2613 684 2616
rect 716 2613 765 2616
rect 796 2613 821 2616
rect 826 2613 844 2616
rect 876 2613 917 2616
rect 954 2613 988 2616
rect 1026 2613 1084 2616
rect 1090 2613 1156 2616
rect 1258 2613 1276 2616
rect 1444 2613 1461 2616
rect 346 2607 349 2613
rect 1090 2607 1093 2613
rect 1458 2607 1461 2613
rect 1482 2613 1516 2616
rect 1546 2613 1572 2616
rect 1642 2615 1645 2633
rect 1658 2626 1661 2633
rect 1658 2623 1700 2626
rect 3004 2623 3013 2626
rect 1804 2613 1845 2616
rect 1884 2613 1941 2616
rect 2324 2613 2349 2616
rect 2404 2613 2437 2616
rect 2442 2613 2468 2616
rect 2548 2613 2573 2616
rect 2604 2613 2613 2616
rect 2756 2613 2773 2616
rect 2970 2613 2988 2616
rect 3026 2613 3084 2616
rect 3116 2613 3133 2616
rect 3220 2613 3245 2616
rect 3282 2613 3356 2616
rect 3434 2613 3444 2616
rect 3490 2613 3516 2616
rect 3548 2613 3621 2616
rect 1482 2607 1485 2613
rect 2434 2606 2437 2613
rect 82 2603 116 2606
rect 634 2603 692 2606
rect 794 2603 852 2606
rect 954 2603 996 2606
rect 1114 2603 1132 2606
rect 1180 2603 1197 2606
rect 1300 2603 1309 2606
rect 1746 2603 1780 2606
rect 1876 2603 1909 2606
rect 1914 2603 2020 2606
rect 2052 2603 2069 2606
rect 2434 2603 2461 2606
rect 2476 2603 2509 2606
rect 2644 2603 2653 2606
rect 2770 2605 2773 2613
rect 2786 2603 2980 2606
rect 3004 2603 3077 2606
rect 3108 2603 3148 2606
rect 3172 2603 3181 2606
rect 3314 2603 3348 2606
rect 3452 2603 3517 2606
rect 3540 2603 3557 2606
rect 3618 2596 3621 2613
rect 3626 2606 3629 2616
rect 3692 2613 3717 2616
rect 3836 2613 3853 2616
rect 3858 2613 3908 2616
rect 3940 2613 3949 2616
rect 4020 2613 4045 2616
rect 4058 2613 4076 2616
rect 4204 2613 4229 2616
rect 4234 2613 4276 2616
rect 4330 2606 4333 2616
rect 4338 2613 4372 2616
rect 4410 2613 4460 2616
rect 4554 2613 4564 2616
rect 4578 2613 4596 2616
rect 4628 2613 4677 2616
rect 3626 2603 3684 2606
rect 3732 2603 3765 2606
rect 3828 2603 3893 2606
rect 3938 2603 4012 2606
rect 4084 2603 4101 2606
rect 4140 2603 4149 2606
rect 4196 2603 4205 2606
rect 4300 2603 4380 2606
rect 4396 2603 4445 2606
rect 4450 2603 4468 2606
rect 4572 2603 4589 2606
rect 4620 2603 4637 2606
rect 132 2593 141 2596
rect 482 2593 524 2596
rect 762 2593 772 2596
rect 3618 2593 3661 2596
rect 3740 2593 3797 2596
rect 4476 2593 4493 2596
rect 38 2567 4837 2573
rect 124 2543 157 2546
rect 636 2543 653 2546
rect 874 2536 877 2544
rect 1074 2543 1084 2546
rect 4220 2543 4253 2546
rect 82 2533 108 2536
rect 362 2533 412 2536
rect 434 2533 516 2536
rect 756 2533 765 2536
rect 812 2533 829 2536
rect 874 2533 924 2536
rect 948 2533 957 2536
rect 994 2533 1004 2536
rect 1026 2533 1085 2536
rect 1284 2533 1309 2536
rect 1338 2533 1396 2536
rect 1412 2533 1461 2536
rect 1506 2533 1548 2536
rect 1602 2533 1620 2536
rect 1658 2533 1668 2536
rect 124 2523 165 2526
rect 354 2523 404 2526
rect 458 2523 508 2526
rect 540 2523 612 2526
rect 754 2523 804 2526
rect 810 2523 852 2526
rect 876 2523 925 2526
rect 978 2523 996 2526
rect 1026 2525 1029 2533
rect 1058 2523 1084 2526
rect 1322 2523 1325 2533
rect 1338 2526 1341 2533
rect 1850 2526 1853 2533
rect 2026 2526 2029 2536
rect 2108 2533 2141 2536
rect 2180 2533 2189 2536
rect 2476 2533 2493 2536
rect 2602 2527 2605 2535
rect 1332 2523 1341 2526
rect 1354 2523 1388 2526
rect 1420 2523 1429 2526
rect 1492 2523 1556 2526
rect 1586 2523 1676 2526
rect 1820 2523 1853 2526
rect 1986 2523 2100 2526
rect 2186 2523 2252 2526
rect 2332 2523 2357 2526
rect 2388 2523 2397 2526
rect 2596 2524 2605 2527
rect 2770 2526 2773 2535
rect 2786 2533 2812 2536
rect 2836 2533 2877 2536
rect 2882 2533 2892 2536
rect 2916 2533 3053 2536
rect 3090 2533 3124 2536
rect 3228 2533 3308 2536
rect 2756 2523 2773 2526
rect 2834 2523 2900 2526
rect 3068 2523 3077 2526
rect 3090 2523 3116 2526
rect 3148 2523 3173 2526
rect 3226 2523 3300 2526
rect 3330 2525 3333 2536
rect 3530 2526 3533 2535
rect 3556 2533 3589 2536
rect 3810 2533 3868 2536
rect 3882 2533 3940 2536
rect 3962 2533 4020 2536
rect 4058 2533 4116 2536
rect 4132 2533 4141 2536
rect 4202 2533 4212 2536
rect 4226 2533 4268 2536
rect 4338 2533 4388 2536
rect 4602 2533 4620 2536
rect 4602 2526 4605 2533
rect 3428 2523 3437 2526
rect 3484 2523 3533 2526
rect 3730 2523 3780 2526
rect 3876 2523 3909 2526
rect 3914 2523 3932 2526
rect 4018 2523 4028 2526
rect 4034 2523 4108 2526
rect 4194 2523 4204 2526
rect 4242 2523 4269 2526
rect 4434 2523 4460 2526
rect 4540 2523 4565 2526
rect 4596 2523 4605 2526
rect 4690 2523 4708 2526
rect 298 2513 324 2516
rect 348 2513 397 2516
rect 756 2513 765 2516
rect 882 2513 924 2516
rect 1172 2513 1181 2516
rect 1948 2513 1957 2516
rect 2836 2513 2869 2516
rect 3154 2513 3204 2516
rect 3570 2513 3596 2516
rect 1178 2503 1181 2513
rect 14 2467 4861 2473
rect 1146 2433 1157 2436
rect 1836 2433 1853 2436
rect 1874 2433 1917 2436
rect 2058 2433 2084 2436
rect 386 2423 428 2426
rect 452 2423 501 2426
rect 1138 2423 1148 2426
rect 100 2413 117 2416
rect 148 2413 205 2416
rect 260 2413 301 2416
rect 316 2413 341 2416
rect 372 2413 421 2416
rect 490 2413 516 2416
rect 580 2413 620 2416
rect 692 2413 709 2416
rect 802 2413 828 2416
rect 858 2413 884 2416
rect 932 2413 949 2416
rect 1004 2413 1045 2416
rect 1066 2413 1100 2416
rect 1154 2415 1157 2433
rect 1794 2423 1828 2426
rect 1858 2423 1908 2426
rect 1260 2413 1269 2416
rect 1316 2413 1325 2416
rect 1388 2413 1429 2416
rect 1540 2413 1565 2416
rect 1596 2413 1605 2416
rect 1914 2415 1917 2433
rect 2018 2423 2068 2426
rect 2092 2423 2101 2426
rect 2282 2423 2301 2426
rect 1938 2413 1980 2416
rect 2170 2413 2236 2416
rect 2396 2413 2405 2416
rect 2418 2413 2445 2416
rect 2450 2413 2492 2416
rect 2594 2413 2660 2416
rect 2690 2413 2716 2416
rect 2836 2413 2861 2416
rect 122 2403 140 2406
rect 162 2403 252 2406
rect 266 2403 308 2406
rect 322 2403 348 2406
rect 380 2403 389 2406
rect 636 2403 653 2406
rect 666 2403 684 2406
rect 770 2403 820 2406
rect 898 2403 924 2406
rect 946 2403 988 2406
rect 1034 2403 1044 2406
rect 1068 2403 1077 2406
rect 1178 2403 1213 2406
rect 1338 2403 1364 2406
rect 1380 2403 1421 2406
rect 1602 2405 1605 2413
rect 2004 2403 2061 2406
rect 2162 2403 2228 2406
rect 2402 2405 2405 2413
rect 2442 2406 2445 2413
rect 2442 2403 2484 2406
rect 2858 2405 2861 2413
rect 2930 2406 2933 2426
rect 2996 2423 3013 2426
rect 4442 2416 4445 2426
rect 4754 2416 4757 2436
rect 2970 2413 2980 2416
rect 3132 2413 3165 2416
rect 3202 2413 3228 2416
rect 3322 2413 3364 2416
rect 3444 2413 3469 2416
rect 3506 2413 3540 2416
rect 3554 2413 3580 2416
rect 3612 2413 3637 2416
rect 3682 2413 3732 2416
rect 3762 2413 3796 2416
rect 3834 2413 3860 2416
rect 3906 2413 3916 2416
rect 3954 2413 3964 2416
rect 4154 2413 4180 2416
rect 4202 2413 4228 2416
rect 4340 2413 4357 2416
rect 2924 2403 2933 2406
rect 2946 2403 2972 2406
rect 2996 2403 3037 2406
rect 3162 2405 3165 2413
rect 3188 2403 3213 2406
rect 3372 2403 3381 2406
rect 3548 2403 3573 2406
rect 3578 2403 3588 2406
rect 3604 2403 3613 2406
rect 3698 2403 3724 2406
rect 3820 2403 3845 2406
rect 3850 2403 3853 2413
rect 4236 2403 4301 2406
rect 4332 2403 4397 2406
rect 4402 2405 4405 2416
rect 4442 2413 4484 2416
rect 4594 2413 4605 2416
rect 4644 2413 4661 2416
rect 4674 2413 4693 2416
rect 4706 2413 4716 2416
rect 4748 2413 4757 2416
rect 4762 2413 4788 2416
rect 4436 2403 4445 2406
rect 4508 2403 4549 2406
rect 4594 2405 4597 2413
rect 4626 2403 4636 2406
rect 4642 2403 4676 2406
rect 4706 2403 4724 2406
rect 4754 2403 4780 2406
rect 3380 2393 3397 2396
rect 4602 2393 4628 2396
rect 1650 2383 1677 2386
rect 1858 2383 1901 2386
rect 38 2367 4837 2373
rect 1698 2353 1733 2356
rect 3220 2343 3269 2346
rect 3610 2343 3629 2346
rect 3900 2343 3965 2346
rect 3610 2336 3613 2343
rect 314 2333 324 2336
rect 354 2333 380 2336
rect 492 2333 517 2336
rect 554 2333 580 2336
rect 842 2333 892 2336
rect 1004 2333 1037 2336
rect 1068 2333 1077 2336
rect 1340 2333 1357 2336
rect 2218 2333 2236 2336
rect 2410 2333 2484 2336
rect 2522 2333 2588 2336
rect 2674 2333 2692 2336
rect 2876 2333 2916 2336
rect 2930 2333 2980 2336
rect 3004 2333 3101 2336
rect 3132 2333 3205 2336
rect 3212 2333 3237 2336
rect 3338 2333 3356 2336
rect 3516 2333 3533 2336
rect 3596 2333 3613 2336
rect 3618 2333 3668 2336
rect 306 2326 309 2333
rect 306 2323 325 2326
rect 340 2323 365 2326
rect 490 2323 540 2326
rect 746 2323 773 2326
rect 842 2323 845 2333
rect 1002 2323 1044 2326
rect 1074 2323 1077 2333
rect 1354 2326 1357 2333
rect 1402 2326 1405 2333
rect 2178 2326 2181 2333
rect 1354 2323 1396 2326
rect 1402 2323 1444 2326
rect 1474 2323 1500 2326
rect 1676 2323 1685 2326
rect 2004 2323 2029 2326
rect 2116 2323 2141 2326
rect 2172 2323 2181 2326
rect 2188 2323 2229 2326
rect 2260 2323 2285 2326
rect 2530 2323 2596 2326
rect 2634 2323 2853 2326
rect 2868 2323 2877 2326
rect 2882 2323 2988 2326
rect 2874 2316 2877 2323
rect 3098 2316 3101 2333
rect 3138 2323 3204 2326
rect 3314 2323 3348 2326
rect 3428 2323 3445 2326
rect 3490 2323 3508 2326
rect 3554 2323 3572 2326
rect 3604 2323 3669 2326
rect 3682 2325 3685 2336
rect 3754 2333 3796 2336
rect 3812 2333 3829 2336
rect 3834 2333 3892 2336
rect 3954 2333 3972 2336
rect 4034 2333 4092 2336
rect 4114 2333 4164 2336
rect 4330 2333 4364 2336
rect 4580 2333 4589 2336
rect 4658 2333 4692 2336
rect 3730 2323 3788 2326
rect 3834 2323 3884 2326
rect 4026 2323 4084 2326
rect 4116 2323 4141 2326
rect 4172 2323 4221 2326
rect 4260 2323 4285 2326
rect 4324 2323 4357 2326
rect 4372 2323 4421 2326
rect 4466 2323 4484 2326
rect 4618 2323 4628 2326
rect 4660 2323 4693 2326
rect 4754 2323 4764 2326
rect 90 2313 100 2316
rect 124 2313 141 2316
rect 154 2313 164 2316
rect 1066 2313 1132 2316
rect 1186 2313 1220 2316
rect 1714 2313 1892 2316
rect 1906 2313 1916 2316
rect 2730 2313 2860 2316
rect 2874 2313 2901 2316
rect 3098 2313 3108 2316
rect 108 2303 125 2306
rect 1140 2303 1229 2306
rect 1900 2303 1965 2306
rect 14 2267 4861 2273
rect 122 2233 172 2236
rect 242 2233 268 2236
rect 1066 2233 1085 2236
rect 1140 2233 1309 2236
rect 138 2223 156 2226
rect 202 2223 252 2226
rect 276 2223 301 2226
rect 426 2223 468 2226
rect 1034 2223 1052 2226
rect 362 2213 396 2216
rect 484 2213 493 2216
rect 730 2206 733 2216
rect 980 2213 1013 2216
rect 1066 2215 1069 2233
rect 1082 2226 1085 2233
rect 1082 2223 1132 2226
rect 1156 2223 1197 2226
rect 2130 2223 2172 2226
rect 2196 2223 2229 2226
rect 2900 2223 2949 2226
rect 2988 2223 3005 2226
rect 3074 2223 3132 2226
rect 1274 2213 1316 2216
rect 1386 2213 1444 2216
rect 1474 2213 1516 2216
rect 1570 2207 1573 2216
rect 1610 2213 1636 2216
rect 1642 2213 1685 2216
rect 1722 2213 1740 2216
rect 1794 2213 1804 2216
rect 1834 2213 1876 2216
rect 1882 2213 1908 2216
rect 1938 2213 1964 2216
rect 1642 2207 1645 2213
rect 1882 2207 1885 2213
rect 2050 2207 2053 2216
rect 2060 2213 2085 2216
rect 2274 2206 2277 2214
rect 2282 2213 2324 2216
rect 2354 2213 2372 2216
rect 2410 2213 2420 2216
rect 2484 2213 2501 2216
rect 2540 2213 2549 2216
rect 2562 2213 2572 2216
rect 2620 2213 2629 2216
rect 2700 2213 2709 2216
rect 2748 2213 2757 2216
rect 2762 2213 2788 2216
rect 2906 2213 2965 2216
rect 2986 2213 3052 2216
rect 3148 2213 3157 2216
rect 348 2203 373 2206
rect 412 2203 429 2206
rect 442 2203 468 2206
rect 492 2203 501 2206
rect 730 2203 748 2206
rect 866 2203 884 2206
rect 932 2203 949 2206
rect 962 2203 972 2206
rect 1298 2203 1324 2206
rect 1340 2203 1429 2206
rect 1530 2203 1572 2206
rect 1604 2203 1621 2206
rect 1650 2203 1684 2206
rect 1748 2203 1773 2206
rect 1778 2203 1796 2206
rect 1828 2203 1845 2206
rect 2234 2203 2252 2206
rect 2274 2203 2309 2206
rect 2380 2203 2405 2206
rect 2546 2205 2549 2213
rect 2708 2203 2741 2206
rect 2866 2203 2876 2206
rect 2900 2203 2957 2206
rect 2962 2205 2965 2213
rect 3202 2206 3205 2216
rect 3210 2213 3252 2216
rect 3338 2213 3348 2216
rect 3436 2213 3477 2216
rect 3522 2213 3580 2216
rect 3618 2213 3660 2216
rect 3690 2213 3716 2216
rect 3772 2213 3789 2216
rect 3884 2213 3893 2216
rect 3996 2213 4021 2216
rect 4058 2213 4084 2216
rect 4122 2213 4212 2216
rect 4250 2213 4268 2216
rect 4314 2213 4332 2216
rect 4364 2213 4389 2216
rect 4428 2213 4445 2216
rect 3618 2206 3621 2213
rect 2988 2203 3037 2206
rect 3068 2203 3117 2206
rect 3156 2203 3173 2206
rect 3202 2203 3260 2206
rect 3276 2203 3325 2206
rect 3378 2203 3412 2206
rect 3604 2203 3621 2206
rect 3906 2203 3932 2206
rect 3954 2203 3988 2206
rect 4362 2203 4420 2206
rect 4484 2203 4540 2206
rect 4546 2203 4549 2214
rect 4596 2213 4605 2216
rect 4692 2213 4757 2216
rect 4604 2203 4613 2206
rect 4658 2203 4684 2206
rect 4754 2203 4757 2213
rect 322 2193 332 2196
rect 442 2193 445 2203
rect 1778 2196 1781 2203
rect 1770 2193 1781 2196
rect 4122 2193 4141 2196
rect 38 2167 4837 2173
rect 436 2143 445 2146
rect 1770 2136 1773 2156
rect 3220 2143 3245 2146
rect 244 2133 253 2136
rect 348 2133 372 2136
rect 386 2133 420 2136
rect 594 2133 612 2136
rect 626 2133 684 2136
rect 722 2133 756 2136
rect 778 2133 828 2136
rect 946 2133 972 2136
rect 1066 2133 1124 2136
rect 1650 2133 1676 2136
rect 1708 2133 1717 2136
rect 1770 2133 1780 2136
rect 2124 2133 2157 2136
rect 2162 2133 2180 2136
rect 2218 2133 2276 2136
rect 2292 2133 2341 2136
rect 2444 2133 2453 2136
rect 386 2126 389 2133
rect 2042 2126 2045 2133
rect 2570 2126 2573 2134
rect 2842 2133 2900 2136
rect 2924 2133 2933 2136
rect 3114 2133 3124 2136
rect 3140 2133 3189 2136
rect 3194 2133 3212 2136
rect 3292 2133 3380 2136
rect 3410 2133 3468 2136
rect 3474 2133 3508 2136
rect 3540 2133 3605 2136
rect 3634 2133 3692 2136
rect 3914 2133 3964 2136
rect 3996 2133 4029 2136
rect 4532 2133 4541 2136
rect 4596 2133 4621 2136
rect 4658 2133 4684 2136
rect 178 2123 196 2126
rect 210 2123 236 2126
rect 370 2123 389 2126
rect 586 2123 620 2126
rect 692 2123 717 2126
rect 738 2123 764 2126
rect 826 2123 836 2126
rect 954 2123 980 2126
rect 90 2113 140 2116
rect 284 2113 301 2116
rect 314 2113 324 2116
rect 994 2113 1028 2116
rect 1042 2106 1045 2125
rect 1132 2123 1141 2126
rect 1292 2123 1301 2126
rect 1372 2123 1389 2126
rect 1572 2123 1597 2126
rect 1634 2123 1684 2126
rect 1714 2123 1788 2126
rect 1882 2123 1908 2126
rect 1980 2123 2005 2126
rect 2036 2123 2045 2126
rect 2052 2123 2085 2126
rect 2116 2123 2188 2126
rect 2250 2123 2268 2126
rect 2306 2123 2340 2126
rect 2562 2123 2573 2126
rect 2580 2123 2589 2126
rect 2596 2123 2637 2126
rect 2780 2123 2797 2126
rect 2850 2123 2908 2126
rect 3106 2123 3116 2126
rect 3154 2123 3204 2126
rect 3218 2123 3268 2126
rect 3404 2123 3445 2126
rect 3482 2123 3516 2126
rect 3554 2123 3604 2126
rect 3636 2123 3653 2126
rect 3700 2123 3725 2126
rect 3762 2123 3788 2126
rect 3842 2123 3972 2126
rect 4066 2123 4084 2126
rect 4292 2123 4325 2126
rect 4404 2123 4429 2126
rect 4466 2123 4476 2126
rect 4588 2123 4605 2126
rect 4618 2123 4628 2126
rect 4692 2123 4701 2126
rect 4754 2123 4764 2126
rect 2562 2116 2565 2123
rect 1146 2113 1212 2116
rect 2482 2113 2500 2116
rect 2524 2113 2565 2116
rect 2634 2106 2637 2123
rect 2674 2113 2684 2116
rect 2708 2113 2741 2116
rect 2924 2113 2949 2116
rect 4618 2113 4621 2123
rect 148 2103 157 2106
rect 258 2103 276 2106
rect 1042 2103 1117 2106
rect 1210 2103 1228 2106
rect 2508 2103 2517 2106
rect 2634 2103 2660 2106
rect 2682 2103 2700 2106
rect 14 2067 4861 2073
rect 1842 2043 1861 2046
rect 2028 2033 2069 2036
rect 2354 2033 2373 2036
rect 1530 2023 1556 2026
rect 1580 2023 1597 2026
rect 1746 2023 1773 2026
rect 1978 2023 2020 2026
rect 2044 2023 2053 2026
rect 2058 2023 2076 2026
rect 2234 2023 2284 2026
rect 2354 2023 2364 2026
rect 122 2013 165 2016
rect 196 2013 213 2016
rect 332 2013 341 2016
rect 820 2013 837 2016
rect 1004 2013 1013 2016
rect 1060 2013 1069 2016
rect 1186 2013 1212 2016
rect 1484 2013 1517 2016
rect 1628 2013 1669 2016
rect 1724 2013 1741 2016
rect 1746 2013 1796 2016
rect 162 2006 165 2013
rect 1514 2007 1517 2013
rect 1634 2006 1637 2013
rect 1826 2006 1829 2014
rect 1834 2013 1868 2016
rect 1874 2007 1877 2016
rect 1916 2013 1941 2016
rect 2156 2013 2181 2016
rect 2212 2013 2221 2016
rect 2370 2015 2373 2033
rect 2388 2023 2397 2026
rect 2594 2023 2604 2026
rect 3026 2016 3029 2026
rect 2402 2013 2428 2016
rect 2458 2013 2484 2016
rect 2516 2013 2525 2016
rect 2530 2013 2556 2016
rect 2610 2013 2636 2016
rect 2748 2013 2765 2016
rect 2842 2013 2860 2016
rect 2874 2013 2916 2016
rect 2218 2007 2221 2013
rect 2986 2006 2989 2014
rect 3026 2013 3060 2016
rect 3106 2013 3124 2016
rect 3162 2013 3204 2016
rect 3242 2013 3292 2016
rect 3346 2013 3389 2016
rect 3428 2013 3453 2016
rect 3508 2013 3533 2016
rect 3842 2013 3868 2016
rect 4138 2013 4156 2016
rect 4234 2013 4268 2016
rect 4274 2013 4316 2016
rect 108 2003 157 2006
rect 162 2003 188 2006
rect 684 2003 701 2006
rect 706 2003 716 2006
rect 868 2003 877 2006
rect 1146 2003 1220 2006
rect 1236 2003 1277 2006
rect 1634 2003 1700 2006
rect 1826 2003 1853 2006
rect 2524 2003 2541 2006
rect 2754 2003 2796 2006
rect 2834 2003 2852 2006
rect 2932 2003 2989 2006
rect 3068 2003 3117 2006
rect 3148 2003 3165 2006
rect 3170 2003 3212 2006
rect 3316 2003 3325 2006
rect 3426 2003 3500 2006
rect 3780 2003 3853 2006
rect 3970 2003 3980 2006
rect 4066 2003 4100 2006
rect 4116 2003 4149 2006
rect 4164 2003 4173 2006
rect 4178 2003 4212 2006
rect 4276 2003 4317 2006
rect 4346 2003 4349 2014
rect 4362 2013 4388 2016
rect 4434 2013 4452 2016
rect 4740 2013 4757 2016
rect 4404 2003 4453 2006
rect 4476 2003 4493 2006
rect 4658 2003 4692 2006
rect 3162 1996 3165 2003
rect 26 1993 100 1996
rect 170 1993 180 1996
rect 234 1993 252 1996
rect 3004 1993 3013 1996
rect 3162 1993 3189 1996
rect 26 1936 29 1993
rect 38 1967 4837 1973
rect 1226 1943 1253 1946
rect 26 1933 76 1936
rect 124 1933 141 1936
rect 162 1933 204 1936
rect 228 1933 237 1936
rect 274 1933 308 1936
rect 1018 1933 1068 1936
rect 1100 1933 1141 1936
rect 1146 1933 1196 1936
rect 1212 1933 1253 1936
rect 1354 1933 1412 1936
rect 1506 1933 1524 1936
rect 138 1915 141 1933
rect 1882 1926 1885 1935
rect 1954 1933 1972 1936
rect 2004 1933 2013 1936
rect 2170 1926 2173 1935
rect 2364 1933 2405 1936
rect 2436 1933 2445 1936
rect 2476 1933 2509 1936
rect 2596 1933 2605 1936
rect 2442 1926 2445 1933
rect 2714 1926 2717 1934
rect 2746 1926 2749 1945
rect 3700 1943 3733 1946
rect 3746 1943 3756 1946
rect 3900 1943 3909 1946
rect 346 1923 468 1926
rect 690 1923 716 1926
rect 842 1923 868 1926
rect 1012 1923 1069 1926
rect 1130 1923 1188 1926
rect 1220 1923 1245 1926
rect 1250 1923 1260 1926
rect 1290 1923 1316 1926
rect 1354 1923 1420 1926
rect 1450 1923 1532 1926
rect 1804 1923 1821 1926
rect 1860 1923 1885 1926
rect 1948 1923 1965 1926
rect 2092 1923 2117 1926
rect 2148 1923 2173 1926
rect 2180 1923 2189 1926
rect 2370 1923 2412 1926
rect 2442 1923 2452 1926
rect 2546 1923 2588 1926
rect 2644 1923 2653 1926
rect 2700 1923 2717 1926
rect 2724 1923 2749 1926
rect 2762 1933 2788 1936
rect 2818 1933 2836 1936
rect 2866 1933 2900 1936
rect 3084 1933 3101 1936
rect 3226 1933 3268 1936
rect 3298 1933 3308 1936
rect 3420 1933 3493 1936
rect 3532 1933 3605 1936
rect 3628 1933 3677 1936
rect 3682 1933 3692 1936
rect 3850 1933 3892 1936
rect 3988 1933 3997 1936
rect 4060 1933 4069 1936
rect 4148 1933 4189 1936
rect 4218 1933 4236 1936
rect 4268 1933 4301 1936
rect 4354 1933 4388 1936
rect 4418 1933 4444 1936
rect 4476 1933 4485 1936
rect 4498 1933 4540 1936
rect 4604 1933 4645 1936
rect 4668 1933 4677 1936
rect 2762 1925 2765 1933
rect 2812 1923 2829 1926
rect 2860 1923 2893 1926
rect 2924 1923 2941 1926
rect 2946 1923 2956 1926
rect 3140 1923 3165 1926
rect 3202 1923 3212 1926
rect 3332 1923 3357 1926
rect 3362 1923 3396 1926
rect 3450 1923 3508 1926
rect 3554 1923 3604 1926
rect 3642 1923 3684 1926
rect 3772 1923 3821 1926
rect 3906 1923 3916 1926
rect 3938 1923 3972 1926
rect 4052 1923 4141 1926
rect 4156 1923 4173 1926
rect 4194 1923 4244 1926
rect 4274 1923 4316 1926
rect 4396 1923 4437 1926
rect 4548 1923 4557 1926
rect 4596 1923 4605 1926
rect 4634 1923 4644 1926
rect 4676 1923 4693 1926
rect 4740 1923 4757 1926
rect 234 1913 244 1916
rect 268 1913 285 1916
rect 298 1913 308 1916
rect 1562 1913 1628 1916
rect 1652 1913 1693 1916
rect 1698 1913 1708 1916
rect 2202 1913 2260 1916
rect 2284 1913 2301 1916
rect 1636 1903 1661 1906
rect 2268 1903 2341 1906
rect 2946 1903 2949 1923
rect 14 1867 4861 1873
rect 114 1833 133 1836
rect 114 1815 117 1833
rect 130 1816 133 1833
rect 338 1823 349 1826
rect 3314 1823 3333 1826
rect 346 1816 349 1823
rect 130 1813 148 1816
rect 154 1813 204 1816
rect 218 1813 252 1816
rect 346 1813 356 1816
rect 636 1813 645 1816
rect 650 1813 692 1816
rect 898 1813 908 1816
rect 946 1813 964 1816
rect 1036 1813 1125 1816
rect 1130 1813 1140 1816
rect 1172 1813 1213 1816
rect 1218 1813 1252 1816
rect 1282 1813 1308 1816
rect 1354 1813 1372 1816
rect 1612 1813 1653 1816
rect 1666 1813 1716 1816
rect 1748 1813 1813 1816
rect 1818 1813 1844 1816
rect 1964 1813 2012 1816
rect 2098 1813 2108 1816
rect 2154 1813 2180 1816
rect 2212 1813 2221 1816
rect 2226 1813 2268 1816
rect 2396 1813 2405 1816
rect 2418 1813 2428 1816
rect 2474 1813 2500 1816
rect 2714 1813 2765 1816
rect 2780 1813 2804 1816
rect 2818 1813 2844 1816
rect 2858 1813 2876 1816
rect 1122 1806 1125 1813
rect 212 1803 244 1806
rect 268 1803 301 1806
rect 1018 1803 1028 1806
rect 1122 1803 1148 1806
rect 1164 1803 1237 1806
rect 1316 1803 1325 1806
rect 1330 1803 1364 1806
rect 1650 1805 1653 1813
rect 1714 1803 1724 1806
rect 1868 1803 1877 1806
rect 1890 1803 1940 1806
rect 2074 1803 2100 1806
rect 2138 1803 2188 1806
rect 2204 1803 2229 1806
rect 2242 1803 2260 1806
rect 2402 1805 2405 1813
rect 2714 1803 2740 1806
rect 1122 1793 1125 1803
rect 1210 1793 1229 1796
rect 2762 1795 2765 1813
rect 2772 1803 2805 1806
rect 2812 1803 2837 1806
rect 2882 1805 2885 1816
rect 2924 1813 2941 1816
rect 3004 1813 3013 1816
rect 3154 1813 3164 1816
rect 3186 1813 3212 1816
rect 3244 1813 3253 1816
rect 3330 1813 3356 1816
rect 3506 1813 3556 1816
rect 3588 1813 3637 1816
rect 3660 1813 3685 1816
rect 3730 1813 3740 1816
rect 3868 1813 3877 1816
rect 3946 1813 3972 1816
rect 4066 1813 4076 1816
rect 4146 1813 4172 1816
rect 4244 1813 4253 1816
rect 4516 1813 4533 1816
rect 4578 1813 4588 1816
rect 4610 1813 4636 1816
rect 4668 1813 4693 1816
rect 4740 1813 4749 1816
rect 2890 1803 2900 1806
rect 2930 1803 2940 1806
rect 2970 1803 2980 1806
rect 2996 1803 3053 1806
rect 3180 1803 3213 1806
rect 3242 1803 3300 1806
rect 3322 1803 3364 1806
rect 3546 1803 3564 1806
rect 3586 1803 3652 1806
rect 3714 1803 3732 1806
rect 3890 1803 3916 1806
rect 3938 1803 3980 1806
rect 4018 1803 4028 1806
rect 4602 1803 4644 1806
rect 4674 1803 4692 1806
rect 1682 1783 1709 1786
rect 2930 1783 2933 1803
rect 3372 1793 3397 1796
rect 4036 1793 4061 1796
rect 38 1767 4837 1773
rect 594 1733 628 1736
rect 740 1733 757 1736
rect 1090 1733 1100 1736
rect 1132 1733 1141 1736
rect 1154 1733 1212 1736
rect 1244 1733 1277 1736
rect 1522 1733 1548 1736
rect 1586 1733 1652 1736
rect 2588 1733 2605 1736
rect 2860 1733 2877 1736
rect 3052 1733 3069 1736
rect 3124 1733 3149 1736
rect 3292 1733 3341 1736
rect 92 1723 109 1726
rect 308 1723 333 1726
rect 460 1723 477 1726
rect 572 1723 581 1726
rect 754 1723 757 1733
rect 2082 1726 2085 1733
rect 2210 1726 2213 1733
rect 828 1723 853 1726
rect 884 1723 925 1726
rect 988 1723 1013 1726
rect 1044 1723 1053 1726
rect 1074 1723 1108 1726
rect 1306 1723 1316 1726
rect 1346 1723 1372 1726
rect 1452 1723 1477 1726
rect 1508 1723 1549 1726
rect 1626 1723 1717 1726
rect 1754 1723 1780 1726
rect 1868 1723 1877 1726
rect 1924 1723 1941 1726
rect 2020 1723 2029 1726
rect 2076 1723 2085 1726
rect 2132 1723 2157 1726
rect 2188 1723 2213 1726
rect 2476 1723 2501 1726
rect 2546 1723 2572 1726
rect 2788 1723 2796 1726
rect 2866 1723 2892 1726
rect 2914 1723 2924 1726
rect 2946 1723 2964 1726
rect 3028 1723 3036 1726
rect 3058 1723 3076 1726
rect 3098 1723 3108 1726
rect 3212 1723 3237 1726
rect 3274 1723 3284 1726
rect 3506 1725 3509 1736
rect 3858 1733 3868 1736
rect 3890 1733 3909 1736
rect 4074 1733 4085 1736
rect 4108 1733 4117 1736
rect 4138 1733 4164 1736
rect 4258 1733 4284 1736
rect 4356 1733 4389 1736
rect 4412 1733 4421 1736
rect 4442 1733 4476 1736
rect 4714 1733 4724 1736
rect 3610 1723 3652 1726
rect 3682 1723 3708 1726
rect 3826 1723 3860 1726
rect 3890 1725 3893 1733
rect 3906 1723 3932 1726
rect 3994 1723 4028 1726
rect 106 1716 109 1723
rect 106 1713 132 1716
rect 156 1713 165 1716
rect 2322 1713 2380 1716
rect 4074 1713 4077 1733
rect 4244 1723 4253 1726
rect 4308 1723 4317 1726
rect 4348 1723 4365 1726
rect 4378 1723 4388 1726
rect 4420 1723 4556 1726
rect 4588 1723 4621 1726
rect 4732 1723 4741 1726
rect 2738 1703 2756 1706
rect 14 1667 4861 1673
rect 162 1623 204 1626
rect 1194 1616 1197 1636
rect 2580 1633 2605 1636
rect 2682 1633 2700 1636
rect 2754 1633 2772 1636
rect 2602 1626 2605 1633
rect 2562 1623 2572 1626
rect 2586 1623 2596 1626
rect 2602 1623 2612 1626
rect 2636 1623 2677 1626
rect 2684 1623 2693 1626
rect 2708 1623 2749 1626
rect 2780 1623 2813 1626
rect 4170 1616 4173 1626
rect 292 1613 317 1616
rect 348 1613 357 1616
rect 764 1613 789 1616
rect 898 1613 981 1616
rect 1020 1613 1037 1616
rect 1076 1613 1101 1616
rect 1108 1613 1117 1616
rect 1180 1613 1213 1616
rect 1316 1613 1333 1616
rect 1378 1613 1404 1616
rect 1434 1613 1460 1616
rect 1498 1613 1557 1616
rect 1562 1613 1652 1616
rect 1682 1613 1732 1616
rect 1746 1613 1796 1616
rect 1834 1613 1884 1616
rect 1914 1613 1932 1616
rect 1946 1613 1956 1616
rect 1970 1613 2020 1616
rect 2050 1613 2108 1616
rect 2138 1613 2188 1616
rect 2436 1613 2468 1616
rect 2482 1613 2493 1616
rect 2786 1613 2828 1616
rect 2874 1613 2892 1616
rect 2986 1613 2996 1616
rect 3042 1613 3052 1616
rect 3090 1613 3109 1616
rect 3116 1613 3125 1616
rect 3130 1613 3140 1616
rect 3228 1613 3253 1616
rect 3284 1613 3333 1616
rect 3372 1614 3405 1616
rect 3370 1613 3405 1614
rect 3444 1613 3477 1616
rect 3570 1613 3580 1616
rect 3716 1613 3741 1616
rect 3772 1613 3781 1616
rect 3786 1613 3812 1616
rect 3892 1613 3909 1616
rect 3948 1613 3973 1616
rect 4012 1613 4021 1616
rect 4060 1613 4085 1616
rect 4122 1613 4132 1616
rect 4170 1613 4197 1616
rect 4372 1613 4397 1616
rect 4442 1613 4492 1616
rect 4524 1613 4549 1616
rect 4588 1613 4613 1616
rect 194 1603 204 1606
rect 474 1603 500 1606
rect 612 1603 629 1606
rect 650 1603 660 1606
rect 474 1593 477 1603
rect 898 1583 901 1613
rect 1098 1607 1101 1613
rect 2482 1606 2485 1613
rect 1138 1603 1156 1606
rect 1188 1603 1285 1606
rect 1322 1603 1340 1606
rect 1506 1603 1516 1606
rect 1530 1603 1580 1606
rect 1602 1603 1644 1606
rect 1820 1603 1845 1606
rect 1858 1603 1876 1606
rect 1964 1603 1981 1606
rect 2050 1603 2100 1606
rect 2154 1603 2180 1606
rect 2450 1603 2485 1606
rect 2490 1603 2508 1606
rect 2868 1603 2885 1606
rect 3090 1583 3093 1613
rect 3098 1603 3108 1606
rect 3338 1603 3348 1606
rect 3370 1603 3373 1613
rect 3970 1606 3973 1613
rect 3386 1603 3436 1606
rect 3530 1603 3588 1606
rect 3604 1603 3613 1606
rect 3794 1603 3820 1606
rect 3970 1603 3988 1606
rect 4156 1603 4181 1606
rect 4194 1605 4197 1613
rect 4444 1603 4493 1606
rect 4530 1603 4580 1606
rect 4652 1603 4661 1606
rect 38 1567 4837 1573
rect 90 1543 100 1546
rect 274 1543 316 1546
rect 706 1536 709 1544
rect 3956 1543 4005 1546
rect 4370 1543 4388 1546
rect 108 1533 125 1536
rect 332 1533 357 1536
rect 370 1533 380 1536
rect 522 1533 532 1536
rect 706 1533 717 1536
rect 756 1533 765 1536
rect 770 1533 836 1536
rect 1378 1533 1396 1536
rect 1492 1533 1509 1536
rect 1762 1533 1789 1536
rect 1852 1533 1885 1536
rect 2202 1533 2236 1536
rect 2268 1533 2293 1536
rect 2434 1533 2444 1536
rect 2684 1533 2693 1536
rect 2844 1533 2869 1536
rect 2890 1533 2964 1536
rect 3002 1533 3092 1536
rect 3108 1533 3125 1536
rect 3266 1533 3301 1536
rect 714 1526 717 1533
rect 1554 1526 1557 1533
rect 2178 1526 2181 1533
rect 340 1523 365 1526
rect 498 1523 524 1526
rect 556 1523 581 1526
rect 610 1523 620 1526
rect 658 1523 684 1526
rect 714 1523 748 1526
rect 802 1523 828 1526
rect 866 1523 892 1526
rect 898 1523 908 1526
rect 954 1523 964 1526
rect 1442 1523 1468 1526
rect 1506 1523 1557 1526
rect 1610 1523 1660 1526
rect 1754 1523 1788 1526
rect 1820 1523 1837 1526
rect 1844 1523 1877 1526
rect 2100 1523 2117 1526
rect 2156 1523 2181 1526
rect 2194 1523 2244 1526
rect 2274 1523 2308 1526
rect 2314 1523 2324 1526
rect 2380 1523 2389 1526
rect 2434 1525 2437 1533
rect 3122 1526 3125 1533
rect 3322 1526 3325 1534
rect 3330 1533 3428 1536
rect 3460 1533 3485 1536
rect 3524 1533 3533 1536
rect 3562 1526 3565 1534
rect 3826 1533 3852 1536
rect 3898 1533 3948 1536
rect 4084 1533 4117 1536
rect 4140 1533 4293 1536
rect 4298 1533 4332 1536
rect 4364 1533 4389 1536
rect 4396 1533 4413 1536
rect 4426 1533 4460 1536
rect 4522 1533 4540 1536
rect 4570 1533 4580 1536
rect 4612 1533 4645 1536
rect 4674 1533 4684 1536
rect 2482 1523 2524 1526
rect 2564 1523 2589 1526
rect 2676 1523 2733 1526
rect 2836 1523 2861 1526
rect 2884 1523 2949 1526
rect 3122 1523 3172 1526
rect 3202 1523 3228 1526
rect 3274 1523 3316 1526
rect 3322 1523 3349 1526
rect 3554 1523 3565 1526
rect 3572 1523 3581 1526
rect 3626 1523 3652 1526
rect 3708 1523 3757 1526
rect 3802 1523 3860 1526
rect 3930 1523 3940 1526
rect 4058 1523 4076 1526
rect 4082 1523 4116 1526
rect 4148 1523 4173 1526
rect 4330 1523 4340 1526
rect 4410 1523 4468 1526
rect 4548 1523 4565 1526
rect 4634 1523 4644 1526
rect 2642 1513 2660 1516
rect 2764 1513 2797 1516
rect 4210 1513 4261 1516
rect 2706 1503 2756 1506
rect 14 1467 4861 1473
rect 4618 1453 4677 1456
rect 1106 1423 1133 1426
rect 2954 1423 2989 1426
rect 3402 1423 3445 1426
rect 1106 1416 1109 1423
rect 2954 1416 2957 1423
rect 116 1413 125 1416
rect 186 1413 212 1416
rect 338 1413 356 1416
rect 388 1413 405 1416
rect 412 1413 429 1416
rect 482 1413 492 1416
rect 522 1413 564 1416
rect 636 1413 645 1416
rect 666 1413 692 1416
rect 178 1403 220 1406
rect 242 1403 268 1406
rect 322 1403 364 1406
rect 386 1403 404 1406
rect 426 1396 429 1413
rect 714 1406 717 1414
rect 730 1413 740 1416
rect 810 1413 860 1416
rect 892 1413 917 1416
rect 964 1413 1037 1416
rect 1076 1413 1109 1416
rect 1114 1406 1117 1416
rect 1164 1413 1220 1416
rect 1250 1413 1309 1416
rect 1348 1413 1365 1416
rect 1444 1413 1469 1416
rect 1628 1413 1661 1416
rect 1668 1413 1685 1416
rect 1906 1413 1932 1416
rect 2076 1413 2101 1416
rect 2132 1413 2165 1416
rect 2170 1413 2180 1416
rect 2234 1413 2244 1416
rect 2314 1413 2340 1416
rect 2698 1413 2724 1416
rect 2820 1413 2877 1416
rect 2916 1414 2957 1416
rect 508 1403 533 1406
rect 538 1403 556 1406
rect 570 1403 620 1406
rect 634 1403 700 1406
rect 714 1403 725 1406
rect 748 1403 781 1406
rect 786 1403 796 1406
rect 850 1403 868 1406
rect 898 1403 956 1406
rect 1010 1403 1052 1406
rect 1068 1403 1117 1406
rect 1268 1403 1325 1406
rect 1354 1403 1380 1406
rect 1658 1405 1661 1413
rect 2874 1406 2877 1413
rect 2914 1413 2957 1414
rect 2970 1413 3029 1416
rect 3036 1413 3045 1416
rect 3180 1413 3205 1416
rect 3268 1413 3277 1416
rect 1690 1403 1716 1406
rect 1756 1403 1773 1406
rect 2138 1403 2172 1406
rect 2210 1403 2252 1406
rect 2282 1403 2292 1406
rect 2364 1403 2373 1406
rect 2450 1403 2460 1406
rect 2706 1403 2732 1406
rect 2738 1403 2796 1406
rect 2874 1403 2892 1406
rect 2914 1403 2917 1413
rect 3026 1405 3029 1413
rect 3330 1406 3333 1414
rect 3468 1413 3509 1416
rect 3514 1413 3532 1416
rect 3570 1413 3604 1416
rect 3634 1413 3660 1416
rect 3706 1413 3732 1416
rect 3804 1413 3821 1416
rect 3858 1413 3884 1416
rect 3946 1413 3956 1416
rect 4052 1413 4061 1416
rect 4108 1413 4125 1416
rect 4164 1413 4173 1416
rect 4178 1413 4188 1416
rect 4236 1413 4253 1416
rect 4476 1413 4501 1416
rect 4546 1413 4580 1416
rect 4612 1413 4637 1416
rect 3570 1406 3573 1413
rect 3066 1403 3092 1406
rect 3130 1403 3172 1406
rect 3186 1403 3244 1406
rect 3290 1403 3333 1406
rect 3370 1403 3444 1406
rect 3556 1403 3573 1406
rect 3698 1403 3740 1406
rect 3762 1403 3796 1406
rect 3938 1403 3964 1406
rect 4156 1403 4165 1406
rect 4250 1403 4268 1406
rect 4284 1403 4301 1406
rect 4314 1403 4468 1406
rect 4490 1403 4516 1406
rect 4532 1403 4541 1406
rect 4570 1403 4573 1413
rect 4578 1403 4588 1406
rect 426 1393 436 1396
rect 636 1393 685 1396
rect 2396 1393 2413 1396
rect 2740 1393 2789 1396
rect 38 1367 4837 1373
rect 218 1336 221 1345
rect 2404 1343 2445 1346
rect 3242 1343 3261 1346
rect 3450 1343 3469 1346
rect 3242 1336 3245 1343
rect 3466 1336 3469 1343
rect 114 1333 172 1336
rect 218 1333 228 1336
rect 242 1333 252 1336
rect 114 1325 117 1333
rect 322 1326 325 1334
rect 394 1333 412 1336
rect 506 1333 516 1336
rect 564 1333 581 1336
rect 636 1333 685 1336
rect 322 1323 364 1326
rect 442 1323 476 1326
rect 546 1323 612 1326
rect 690 1323 693 1334
rect 716 1333 725 1336
rect 764 1333 845 1336
rect 868 1333 885 1336
rect 1034 1333 1052 1336
rect 1090 1333 1140 1336
rect 1266 1333 1284 1336
rect 1300 1333 1309 1336
rect 1266 1326 1269 1333
rect 714 1323 756 1326
rect 876 1323 925 1326
rect 1004 1323 1013 1326
rect 1098 1323 1132 1326
rect 1164 1323 1205 1326
rect 1220 1323 1269 1326
rect 1362 1326 1365 1334
rect 1498 1333 1508 1336
rect 1530 1333 1572 1336
rect 1762 1333 1788 1336
rect 1834 1333 1845 1336
rect 1362 1323 1388 1326
rect 1418 1323 1444 1326
rect 1482 1323 1516 1326
rect 1554 1323 1564 1326
rect 1682 1323 1692 1326
rect 1778 1323 1796 1326
rect 682 1313 692 1316
rect 1834 1306 1837 1333
rect 1914 1326 1917 1334
rect 1970 1333 1988 1336
rect 2010 1333 2060 1336
rect 2098 1333 2132 1336
rect 2178 1333 2220 1336
rect 2306 1333 2332 1336
rect 2346 1333 2396 1336
rect 2410 1333 2452 1336
rect 2476 1333 2508 1336
rect 2530 1333 2548 1336
rect 2626 1333 2676 1336
rect 2914 1333 2940 1336
rect 2956 1333 2965 1336
rect 3004 1333 3021 1336
rect 3228 1333 3245 1336
rect 3250 1333 3268 1336
rect 3412 1333 3461 1336
rect 3466 1333 3492 1336
rect 3530 1333 3556 1336
rect 3746 1333 3788 1336
rect 3938 1333 3948 1336
rect 4316 1333 4349 1336
rect 4372 1333 4397 1336
rect 4530 1333 4540 1336
rect 4602 1333 4660 1336
rect 4714 1333 4724 1336
rect 1970 1326 1973 1333
rect 1842 1323 1868 1326
rect 1874 1323 1917 1326
rect 1924 1323 1973 1326
rect 2012 1323 2053 1326
rect 2058 1323 2068 1326
rect 2114 1323 2124 1326
rect 2474 1323 2500 1326
rect 2612 1323 2637 1326
rect 2756 1323 2781 1326
rect 2818 1323 2852 1326
rect 2900 1323 2925 1326
rect 2964 1323 2973 1326
rect 3098 1323 3124 1326
rect 3322 1323 3340 1326
rect 3420 1323 3437 1326
rect 3516 1323 3533 1326
rect 3586 1323 3628 1326
rect 3674 1323 3684 1326
rect 3834 1323 3860 1326
rect 3956 1323 3973 1326
rect 4018 1323 4036 1326
rect 4228 1323 4253 1326
rect 4290 1323 4308 1326
rect 4338 1323 4348 1326
rect 4380 1323 4397 1326
rect 4452 1323 4469 1326
rect 4548 1323 4613 1326
rect 4684 1323 4693 1326
rect 4732 1323 4741 1326
rect 2250 1313 2276 1316
rect 1834 1303 1845 1306
rect 14 1267 4861 1273
rect 516 1223 533 1226
rect 538 1223 548 1226
rect 562 1223 588 1226
rect 602 1223 692 1226
rect 1820 1223 1869 1226
rect 530 1216 533 1223
rect 98 1213 108 1216
rect 228 1213 253 1216
rect 316 1213 341 1216
rect 410 1213 436 1216
rect 474 1213 500 1216
rect 530 1213 556 1216
rect 682 1213 700 1216
rect 74 1203 100 1206
rect 114 1203 124 1206
rect 290 1203 308 1206
rect 330 1203 348 1206
rect 482 1203 492 1206
rect 564 1203 581 1206
rect 604 1203 661 1206
rect 708 1203 725 1206
rect 826 1203 844 1206
rect 890 1205 893 1216
rect 948 1213 973 1216
rect 1028 1213 1069 1216
rect 1164 1213 1189 1216
rect 1226 1213 1260 1216
rect 1290 1213 1340 1216
rect 1420 1213 1445 1216
rect 1476 1213 1509 1216
rect 1516 1213 1533 1216
rect 1618 1213 1660 1216
rect 1010 1203 1020 1206
rect 1058 1203 1068 1206
rect 1290 1203 1332 1206
rect 1506 1205 1509 1213
rect 1530 1203 1533 1213
rect 1634 1203 1652 1206
rect 1730 1203 1733 1214
rect 2020 1213 2061 1216
rect 2156 1213 2173 1216
rect 2212 1213 2237 1216
rect 2274 1213 2284 1216
rect 2442 1213 2452 1216
rect 1756 1203 1773 1206
rect 1970 1203 1996 1206
rect 2034 1203 2037 1213
rect 2292 1203 2309 1206
rect 2442 1203 2460 1206
rect 2482 1203 2485 1214
rect 2490 1213 2500 1216
rect 2666 1213 2684 1216
rect 2780 1213 2813 1216
rect 2852 1213 2861 1216
rect 3026 1213 3060 1216
rect 3346 1213 3396 1216
rect 3442 1213 3452 1216
rect 3524 1213 3549 1216
rect 3588 1213 3653 1216
rect 3660 1213 3677 1216
rect 3682 1213 3724 1216
rect 3820 1213 3861 1216
rect 3924 1213 3957 1216
rect 3994 1213 4020 1216
rect 4100 1213 4133 1216
rect 4186 1213 4212 1216
rect 4252 1213 4261 1216
rect 4298 1213 4324 1216
rect 4396 1213 4421 1216
rect 4474 1213 4484 1216
rect 2810 1206 2813 1213
rect 2708 1203 2756 1206
rect 2810 1203 2828 1206
rect 3084 1203 3237 1206
rect 3530 1203 3564 1206
rect 3594 1203 3652 1206
rect 3666 1203 3732 1206
rect 3748 1203 3796 1206
rect 3834 1203 3884 1206
rect 3906 1203 3916 1206
rect 4106 1203 4148 1206
rect 4164 1203 4181 1206
rect 4468 1203 4485 1206
rect 4514 1203 4517 1214
rect 4610 1213 4636 1216
rect 4730 1213 4756 1216
rect 4522 1203 4540 1206
rect 4674 1203 4684 1206
rect 38 1167 4837 1173
rect 634 1143 653 1146
rect 2524 1143 2565 1146
rect 650 1136 653 1143
rect 290 1133 332 1136
rect 354 1133 405 1136
rect 418 1133 428 1136
rect 452 1133 477 1136
rect 628 1133 645 1136
rect 650 1133 668 1136
rect 1106 1127 1109 1135
rect 1130 1133 1140 1136
rect 1178 1133 1228 1136
rect 1244 1133 1269 1136
rect 1450 1133 1508 1136
rect 1612 1133 1661 1136
rect 1802 1133 1812 1136
rect 172 1123 181 1126
rect 186 1123 196 1126
rect 354 1123 372 1126
rect 394 1123 436 1126
rect 572 1123 581 1126
rect 676 1123 693 1126
rect 780 1123 805 1126
rect 948 1123 973 1126
rect 1044 1123 1069 1126
rect 1100 1124 1109 1127
rect 1978 1126 1981 1135
rect 2018 1133 2084 1136
rect 2114 1133 2196 1136
rect 2210 1133 2244 1136
rect 2434 1133 2516 1136
rect 2580 1133 2629 1136
rect 2652 1133 2677 1136
rect 2844 1133 2885 1136
rect 2018 1126 2021 1133
rect 2914 1126 2917 1136
rect 2986 1133 3004 1136
rect 3036 1133 3061 1136
rect 3066 1133 3076 1136
rect 3210 1133 3220 1136
rect 1116 1123 1133 1126
rect 1164 1123 1189 1126
rect 1210 1123 1220 1126
rect 1252 1123 1285 1126
rect 1380 1123 1405 1126
rect 1442 1123 1516 1126
rect 1578 1123 1588 1126
rect 1620 1123 1637 1126
rect 1692 1123 1756 1126
rect 1786 1123 1820 1126
rect 1892 1123 1917 1126
rect 1948 1123 1981 1126
rect 1988 1123 2021 1126
rect 2050 1123 2076 1126
rect 2252 1123 2269 1126
rect 2498 1123 2508 1126
rect 2554 1123 2572 1126
rect 2602 1123 2628 1126
rect 2660 1123 2685 1126
rect 2740 1123 2765 1126
rect 2802 1123 2836 1126
rect 2842 1123 2884 1126
rect 2914 1125 2949 1126
rect 2916 1123 2949 1125
rect 3148 1123 3173 1126
rect 3242 1125 3245 1136
rect 3380 1133 3421 1136
rect 3436 1133 3469 1136
rect 3508 1133 3533 1136
rect 3250 1123 3292 1126
rect 3306 1123 3356 1126
rect 3428 1123 3445 1126
rect 3458 1123 3484 1126
rect 3514 1123 3532 1126
rect 3562 1125 3565 1136
rect 3706 1133 3724 1136
rect 3746 1133 3796 1136
rect 3900 1133 3956 1136
rect 3978 1133 4020 1136
rect 4066 1133 4076 1136
rect 4092 1133 4148 1136
rect 4234 1133 4252 1136
rect 4290 1133 4316 1136
rect 4458 1133 4532 1136
rect 4610 1133 4644 1136
rect 4666 1133 4684 1136
rect 3626 1123 3652 1126
rect 3690 1123 3716 1126
rect 3804 1123 3837 1126
rect 3906 1123 3948 1126
rect 3986 1123 4028 1126
rect 4042 1123 4068 1126
rect 4146 1123 4156 1126
rect 4218 1123 4244 1126
rect 4282 1123 4324 1126
rect 4380 1123 4389 1126
rect 4436 1123 4493 1126
rect 4498 1123 4540 1126
rect 4570 1123 4636 1126
rect 4738 1123 4756 1126
rect 594 1113 604 1116
rect 690 1115 693 1123
rect 1316 1113 1325 1116
rect 2018 1113 2021 1123
rect 4498 1116 4501 1123
rect 4474 1113 4501 1116
rect 14 1067 4861 1073
rect 3010 1053 3037 1056
rect 242 1023 276 1026
rect 402 1023 428 1026
rect 1602 1023 1628 1026
rect 1794 1023 1828 1026
rect 2066 1023 2092 1026
rect 2116 1023 2125 1026
rect 2258 1023 2284 1026
rect 2906 1023 2925 1026
rect 2906 1016 2909 1023
rect 172 1013 189 1016
rect 194 1013 204 1016
rect 236 1013 269 1016
rect 436 1013 453 1016
rect 914 1013 924 1016
rect 972 1013 997 1016
rect 1044 1013 1069 1016
rect 1100 1013 1109 1016
rect 1116 1013 1157 1016
rect 1210 1013 1252 1016
rect 1282 1013 1316 1016
rect 1372 1013 1421 1016
rect 1436 1013 1461 1016
rect 1732 1013 1757 1016
rect 1788 1013 1805 1016
rect 1866 1013 1900 1016
rect 1930 1013 1989 1016
rect 2122 1013 2148 1016
rect 2322 1013 2357 1016
rect 2418 1013 2428 1016
rect 2466 1013 2484 1016
rect 2530 1013 2564 1016
rect 2748 1013 2797 1016
rect 2836 1013 2861 1016
rect 2892 1013 2909 1016
rect 2914 1013 2940 1016
rect 2996 1013 3156 1016
rect 3188 1013 3228 1016
rect 3260 1013 3277 1016
rect 3292 1013 3309 1016
rect 3354 1013 3380 1016
rect 3426 1013 3436 1016
rect 3586 1013 3596 1016
rect 3634 1013 3668 1016
rect 3762 1013 3804 1016
rect 3834 1013 3860 1016
rect 4036 1013 4061 1016
rect 4098 1013 4108 1016
rect 4114 1013 4164 1016
rect 4202 1013 4228 1016
rect 4458 1013 4468 1016
rect 4546 1013 4572 1016
rect 4610 1013 4636 1016
rect 212 1003 221 1006
rect 228 1003 245 1006
rect 770 1003 796 1006
rect 1106 1005 1109 1013
rect 4202 1006 4205 1013
rect 1130 1003 1164 1006
rect 1234 1003 1244 1006
rect 1298 1003 1308 1006
rect 1322 1003 1364 1006
rect 1442 1003 1468 1006
rect 1506 1003 1556 1006
rect 1964 1003 1973 1006
rect 2002 1003 2012 1006
rect 2044 1003 2053 1006
rect 2156 1003 2181 1006
rect 2266 1003 2284 1006
rect 2308 1003 2436 1006
rect 2452 1003 2477 1006
rect 2668 1003 2709 1006
rect 2756 1003 2805 1006
rect 2828 1003 2868 1006
rect 2900 1003 2909 1006
rect 2948 1003 2965 1006
rect 3066 1003 3164 1006
rect 3180 1003 3229 1006
rect 3258 1003 3284 1006
rect 3418 1003 3428 1006
rect 3572 1003 3589 1006
rect 3620 1003 3653 1006
rect 4188 1003 4205 1006
rect 4396 1003 4469 1006
rect 4492 1003 4564 1006
rect 4596 1003 4637 1006
rect 4660 1003 4701 1006
rect 3042 993 3109 996
rect 3114 993 3117 1003
rect 38 967 4837 973
rect 1498 936 1501 946
rect 204 933 213 936
rect 210 926 213 933
rect 258 926 261 935
rect 290 933 300 936
rect 674 933 708 936
rect 868 933 877 936
rect 882 933 900 936
rect 1410 933 1444 936
rect 1476 933 1501 936
rect 1658 933 1692 936
rect 1780 933 1805 936
rect 1826 933 1852 936
rect 1994 933 2012 936
rect 2044 933 2077 936
rect 2228 933 2269 936
rect 2396 933 2429 936
rect 2524 933 2533 936
rect 2538 933 2548 936
rect 2570 933 2596 936
rect 2618 933 2628 936
rect 2642 933 2700 936
rect 66 923 84 926
rect 122 923 140 926
rect 210 923 221 926
rect 228 923 237 926
rect 252 923 261 926
rect 290 923 317 926
rect 370 923 396 926
rect 466 923 492 926
rect 572 923 597 926
rect 628 923 637 926
rect 706 923 716 926
rect 756 923 781 926
rect 812 923 829 926
rect 860 923 908 926
rect 1044 923 1053 926
rect 1212 923 1237 926
rect 1268 923 1301 926
rect 1306 923 1316 926
rect 1540 923 1565 926
rect 1596 923 1613 926
rect 1690 923 1700 926
rect 1738 923 1756 926
rect 1786 923 1812 926
rect 1868 923 1877 926
rect 2010 923 2020 926
rect 2220 923 2245 926
rect 2258 923 2276 926
rect 2282 923 2292 926
rect 2460 923 2493 926
rect 2578 923 2588 926
rect 2636 923 2661 926
rect 2682 923 2692 926
rect 2722 925 2725 936
rect 2970 933 2988 936
rect 3140 933 3149 936
rect 3266 933 3276 936
rect 3298 933 3324 936
rect 3522 933 3580 936
rect 3610 933 3652 936
rect 3666 933 3716 936
rect 3772 933 3813 936
rect 3842 933 3852 936
rect 3986 933 4004 936
rect 4156 933 4165 936
rect 4436 933 4461 936
rect 2852 923 2861 926
rect 2908 923 2917 926
rect 2964 923 2989 926
rect 2996 923 3021 926
rect 3060 923 3085 926
rect 3122 923 3132 926
rect 3300 923 3309 926
rect 3332 923 3341 926
rect 3386 923 3404 926
rect 3458 923 3508 926
rect 3522 923 3572 926
rect 3604 923 3645 926
rect 3660 923 3717 926
rect 3778 923 3820 926
rect 3922 923 3948 926
rect 3994 923 4012 926
rect 4050 923 4068 926
rect 4228 923 4253 926
rect 4284 923 4293 926
rect 4332 923 4357 926
rect 4394 923 4428 926
rect 4466 925 4469 936
rect 4492 933 4540 936
rect 4572 933 4589 936
rect 4634 933 4652 936
rect 4500 923 4525 926
rect 4594 923 4604 926
rect 4636 923 4653 926
rect 4660 923 4693 926
rect 4730 923 4756 926
rect 290 916 293 923
rect 2258 916 2261 923
rect 276 913 293 916
rect 2234 913 2261 916
rect 2474 913 2500 916
rect 2578 903 2581 923
rect 14 867 4861 873
rect 866 823 876 826
rect 1770 823 1796 826
rect 2562 823 2580 826
rect 74 813 84 816
rect 122 813 140 816
rect 260 813 317 816
rect 324 813 341 816
rect 426 813 468 816
rect 498 813 524 816
rect 242 803 252 806
rect 306 803 316 806
rect 338 795 341 813
rect 348 803 357 806
rect 388 803 397 806
rect 714 803 732 806
rect 770 803 804 806
rect 826 803 829 814
rect 844 813 853 816
rect 906 813 948 816
rect 978 813 996 816
rect 1042 813 1053 816
rect 1090 813 1149 816
rect 1316 813 1325 816
rect 1372 813 1397 816
rect 1428 813 1437 816
rect 1444 813 1493 816
rect 1596 813 1621 816
rect 1652 813 1661 816
rect 1698 813 1748 816
rect 1858 813 1884 816
rect 1956 813 1964 816
rect 2010 813 2028 816
rect 2058 813 2076 816
rect 2298 813 2316 816
rect 2380 813 2428 816
rect 2460 813 2493 816
rect 1042 806 1045 813
rect 972 803 989 806
rect 1004 803 1045 806
rect 1148 803 1157 806
rect 1178 803 1196 806
rect 1434 805 1437 813
rect 2514 806 2517 814
rect 2652 813 2661 816
rect 2772 813 2797 816
rect 2834 813 2844 816
rect 2850 813 2900 816
rect 2932 813 2949 816
rect 3026 813 3052 816
rect 3090 813 3100 816
rect 3164 813 3197 816
rect 3210 813 3220 816
rect 3226 813 3244 816
rect 3538 813 3556 816
rect 3588 813 3605 816
rect 3618 813 3644 816
rect 3826 813 3836 816
rect 3868 813 3909 816
rect 3916 813 3925 816
rect 3972 813 3997 816
rect 4034 813 4052 816
rect 4058 813 4076 816
rect 1458 803 1492 806
rect 1524 803 1541 806
rect 1730 803 1740 806
rect 1922 803 1940 806
rect 2052 803 2061 806
rect 2090 803 2140 806
rect 2250 803 2260 806
rect 2266 803 2276 806
rect 2300 803 2309 806
rect 2324 803 2341 806
rect 2418 803 2436 806
rect 2466 803 2508 806
rect 2514 803 2524 806
rect 2548 803 2573 806
rect 2604 803 2613 806
rect 2852 803 2901 806
rect 3130 803 3140 806
rect 3162 803 3212 806
rect 3498 803 3508 806
rect 3530 803 3564 806
rect 3682 803 3772 806
rect 3788 803 3821 806
rect 3826 803 3844 806
rect 3866 803 3908 806
rect 4060 803 4077 806
rect 4106 803 4109 814
rect 4122 813 4132 816
rect 4226 813 4268 816
rect 4314 813 4324 816
rect 4396 813 4421 816
rect 4466 813 4492 816
rect 4562 813 4572 816
rect 4620 813 4629 816
rect 4692 813 4701 816
rect 4738 813 4764 816
rect 4250 803 4276 806
rect 4468 803 4493 806
rect 4516 803 4564 806
rect 4596 803 4605 806
rect 4626 803 4644 806
rect 4666 803 4684 806
rect 370 793 380 796
rect 38 767 4837 773
rect 594 726 597 735
rect 626 733 644 736
rect 682 733 716 736
rect 738 733 764 736
rect 794 733 836 736
rect 890 733 908 736
rect 970 726 973 736
rect 1018 733 1044 736
rect 1058 733 1092 736
rect 1130 733 1140 736
rect 220 723 237 726
rect 324 723 341 726
rect 380 723 389 726
rect 532 723 557 726
rect 588 723 597 726
rect 604 723 637 726
rect 668 723 685 726
rect 724 723 749 726
rect 802 723 828 726
rect 874 723 900 726
rect 932 725 973 726
rect 932 723 972 725
rect 1004 723 1029 726
rect 1034 723 1100 726
rect 1162 725 1165 736
rect 1276 733 1293 736
rect 1306 733 1316 736
rect 1514 733 1572 736
rect 1714 726 1717 736
rect 1218 723 1252 726
rect 1282 723 1324 726
rect 1388 723 1413 726
rect 1444 723 1493 726
rect 1498 723 1564 726
rect 1596 723 1637 726
rect 1674 725 1717 726
rect 1746 725 1749 736
rect 2218 733 2236 736
rect 2260 733 2285 736
rect 2460 733 2477 736
rect 2492 733 2524 736
rect 2556 733 2589 736
rect 2690 726 2693 735
rect 2780 733 2821 736
rect 2860 733 2901 736
rect 2938 733 2957 736
rect 2986 733 2996 736
rect 3436 733 3453 736
rect 3468 733 3485 736
rect 3524 733 3557 736
rect 3562 733 3572 736
rect 3594 733 3652 736
rect 4060 733 4077 736
rect 4100 733 4148 736
rect 4220 733 4229 736
rect 4258 733 4300 736
rect 4316 733 4372 736
rect 4476 733 4485 736
rect 4508 733 4556 736
rect 4588 733 4597 736
rect 4636 733 4645 736
rect 4650 733 4660 736
rect 1674 723 1716 725
rect 1794 723 1804 726
rect 1834 723 1860 726
rect 1930 723 1940 726
rect 2028 723 2037 726
rect 2202 723 2244 726
rect 2306 723 2324 726
rect 2458 723 2484 726
rect 2538 723 2548 726
rect 2628 723 2637 726
rect 2684 723 2693 726
rect 2786 723 2836 726
rect 2866 723 2900 726
rect 2932 723 2949 726
rect 2954 725 2957 733
rect 2988 723 2997 726
rect 3004 723 3021 726
rect 3058 723 3084 726
rect 3156 723 3165 726
rect 3212 723 3221 726
rect 3330 723 3340 726
rect 3442 723 3460 726
rect 3466 723 3500 726
rect 3596 723 3613 726
rect 3660 723 3685 726
rect 3972 723 3997 726
rect 4034 723 4052 726
rect 4130 723 4140 726
rect 4186 723 4212 726
rect 4218 723 4228 726
rect 4266 723 4292 726
rect 4338 723 4380 726
rect 4458 723 4468 726
rect 4474 723 4484 726
rect 4594 723 4612 726
rect 4682 725 4685 736
rect 4738 723 4764 726
rect 1610 713 1644 716
rect 1668 713 1709 716
rect 14 667 4861 673
rect 1146 633 1181 636
rect 332 623 341 626
rect 1146 623 1172 626
rect 220 613 229 616
rect 276 613 285 616
rect 292 613 316 616
rect 338 613 348 616
rect 372 613 381 616
rect 442 613 468 616
rect 548 613 573 616
rect 684 613 749 616
rect 756 613 813 616
rect 1082 613 1108 616
rect 1178 615 1181 633
rect 2202 626 2205 646
rect 1196 623 1213 626
rect 1258 623 1284 626
rect 2196 623 2205 626
rect 2410 623 2420 626
rect 2530 623 2540 626
rect 1322 613 1356 616
rect 1386 613 1444 616
rect 1474 613 1517 616
rect 1530 613 1564 616
rect 1660 613 1693 616
rect 1698 613 1708 616
rect 1762 613 1772 616
rect 1924 613 1949 616
rect 1980 613 1997 616
rect 2004 613 2021 616
rect 2066 613 2100 616
rect 2202 613 2244 616
rect 2258 613 2300 616
rect 2322 613 2340 616
rect 2436 613 2445 616
rect 2450 613 2484 616
rect 2562 613 2596 616
rect 2618 613 2628 616
rect 2682 613 2692 616
rect 2756 613 2781 616
rect 2866 613 2876 616
rect 2924 613 2940 616
rect 2972 613 2997 616
rect 3162 613 3188 616
rect 3274 613 3308 616
rect 3340 613 3349 616
rect 3618 613 3636 616
rect 3682 613 3692 616
rect 3754 613 3788 616
rect 3924 613 3949 616
rect 3994 613 4044 616
rect 4116 613 4141 616
rect 4178 613 4188 616
rect 4268 613 4293 616
rect 4330 613 4340 616
rect 4346 613 4364 616
rect 4396 613 4413 616
rect 4452 613 4461 616
rect 4570 613 4588 616
rect 4626 613 4644 616
rect 4676 613 4685 616
rect 4730 613 4756 616
rect 282 605 285 613
rect 298 603 308 606
rect 386 603 396 606
rect 412 603 437 606
rect 626 603 660 606
rect 692 603 733 606
rect 810 603 813 613
rect 1244 603 1269 606
rect 1418 603 1436 606
rect 1468 603 1485 606
rect 1490 603 1500 606
rect 1580 603 1597 606
rect 1626 603 1644 606
rect 1666 603 1700 606
rect 1748 603 1757 606
rect 1994 605 1997 613
rect 2018 606 2021 613
rect 3754 606 3757 613
rect 2018 603 2036 606
rect 2154 603 2172 606
rect 2202 603 2236 606
rect 2260 603 2277 606
rect 2316 603 2325 606
rect 2396 603 2413 606
rect 2450 603 2476 606
rect 2514 603 2540 606
rect 2610 603 2620 606
rect 2652 603 2661 606
rect 2852 603 2861 606
rect 2930 603 2948 606
rect 3164 603 3181 606
rect 3196 603 3213 606
rect 3276 603 3293 606
rect 3298 603 3316 606
rect 3338 603 3364 606
rect 3484 603 3525 606
rect 3548 603 3557 606
rect 3570 603 3588 606
rect 3604 603 3629 606
rect 3748 603 3765 606
rect 3812 603 3821 606
rect 3890 603 3900 606
rect 3938 603 3964 606
rect 3996 603 4052 606
rect 4394 603 4413 606
rect 4570 603 4596 606
rect 4674 603 4684 606
rect 2860 593 2869 596
rect 3202 583 3221 586
rect 38 567 4837 573
rect 138 543 164 546
rect 130 533 172 536
rect 268 533 293 536
rect 346 526 349 535
rect 530 533 556 536
rect 636 533 645 536
rect 762 533 788 536
rect 820 533 868 536
rect 900 533 917 536
rect 1050 533 1060 536
rect 1226 526 1229 535
rect 1276 533 1301 536
rect 1404 533 1413 536
rect 1522 533 1580 536
rect 1596 533 1645 536
rect 1740 533 1765 536
rect 1850 533 1868 536
rect 1898 533 1908 536
rect 1980 533 2028 536
rect 1898 526 1901 533
rect 2218 526 2221 535
rect 340 523 349 526
rect 394 523 436 526
rect 466 523 492 526
rect 564 523 589 526
rect 628 523 653 526
rect 692 523 717 526
rect 754 523 796 526
rect 898 523 973 526
rect 1068 523 1101 526
rect 1148 523 1173 526
rect 1204 523 1229 526
rect 1268 523 1277 526
rect 1282 523 1316 526
rect 1604 523 1644 526
rect 1682 523 1781 526
rect 1884 523 1901 526
rect 1924 523 1933 526
rect 1972 523 1997 526
rect 2002 523 2036 526
rect 2066 523 2076 526
rect 2140 523 2165 526
rect 2196 523 2221 526
rect 2266 526 2269 535
rect 2274 533 2316 536
rect 2362 533 2396 536
rect 2644 533 2661 536
rect 2786 526 2789 535
rect 2810 533 2820 536
rect 2860 533 2933 536
rect 2954 533 2988 536
rect 3084 533 3117 536
rect 3162 533 3204 536
rect 2266 523 2285 526
rect 2314 523 2324 526
rect 2498 523 2565 526
rect 2756 523 2789 526
rect 2852 523 2861 526
rect 2996 523 3037 526
rect 3076 523 3109 526
rect 3154 523 3196 526
rect 3226 525 3229 536
rect 3506 533 3524 536
rect 3556 533 3573 536
rect 3602 533 3620 536
rect 3812 533 3861 536
rect 3884 533 3917 536
rect 3986 533 4012 536
rect 4058 533 4100 536
rect 4252 533 4285 536
rect 4290 533 4324 536
rect 4426 533 4460 536
rect 4674 533 4764 536
rect 3276 523 3293 526
rect 3330 523 3356 526
rect 3444 523 3469 526
rect 3514 523 3532 526
rect 3604 523 3613 526
rect 3666 523 3692 526
rect 3786 523 3804 526
rect 3898 523 3932 526
rect 3964 523 3981 526
rect 4090 523 4108 526
rect 4202 523 4236 526
rect 4290 523 4293 533
rect 4332 523 4389 526
rect 4468 523 4509 526
rect 4618 523 4644 526
rect 4676 523 4685 526
rect 4746 523 4772 526
rect 66 513 100 516
rect 124 513 141 516
rect 946 513 988 516
rect 2340 513 2349 516
rect 2890 483 2925 486
rect 14 467 4861 473
rect 834 433 852 436
rect 970 433 996 436
rect 124 423 141 426
rect 154 416 157 425
rect 252 423 260 426
rect 826 423 836 426
rect 860 423 901 426
rect 962 423 980 426
rect 2818 423 2828 426
rect 82 413 108 416
rect 130 413 148 416
rect 154 413 189 416
rect 204 413 229 416
rect 268 413 285 416
rect 330 413 372 416
rect 596 413 629 416
rect 690 413 780 416
rect 178 403 196 406
rect 226 405 229 413
rect 276 403 357 406
rect 570 403 588 406
rect 706 403 772 406
rect 786 403 789 414
rect 866 413 916 416
rect 1010 413 1020 416
rect 1050 413 1108 416
rect 1114 413 1180 416
rect 1284 413 1309 416
rect 1340 413 1357 416
rect 1402 413 1420 416
rect 1452 413 1533 416
rect 1540 413 1557 416
rect 1948 413 1973 416
rect 2004 413 2021 416
rect 2082 413 2092 416
rect 2170 413 2188 416
rect 2282 413 2308 416
rect 2402 413 2420 416
rect 2612 413 2637 416
rect 2668 413 2693 416
rect 2738 413 2748 416
rect 1554 406 1557 413
rect 2082 406 2085 413
rect 1044 403 1077 406
rect 1082 403 1100 406
rect 1204 403 1229 406
rect 1346 403 1364 406
rect 1410 403 1428 406
rect 1522 403 1532 406
rect 1554 403 1572 406
rect 1588 403 1605 406
rect 1660 403 1701 406
rect 1706 403 1716 406
rect 1748 403 1773 406
rect 1778 403 1820 406
rect 1892 403 1901 406
rect 2026 403 2036 406
rect 2052 403 2085 406
rect 2106 403 2124 406
rect 2156 403 2173 406
rect 2690 405 2693 413
rect 2818 406 2821 423
rect 2858 413 2892 416
rect 2978 413 3004 416
rect 3076 413 3101 416
rect 3146 413 3156 416
rect 3188 414 3268 416
rect 3188 413 3269 414
rect 3300 413 3325 416
rect 3362 413 3380 416
rect 3436 413 3445 416
rect 3482 413 3508 416
rect 3610 413 3636 416
rect 3700 413 3725 416
rect 3764 413 3789 416
rect 3876 413 3901 416
rect 3938 413 3964 416
rect 3986 413 4004 416
rect 4130 413 4172 416
rect 4194 413 4220 416
rect 4250 413 4276 416
rect 4308 413 4317 416
rect 4338 413 4364 416
rect 4394 413 4420 416
rect 4466 413 4476 416
rect 4506 413 4532 416
rect 4570 413 4604 416
rect 4666 413 4700 416
rect 4746 413 4756 416
rect 2706 403 2740 406
rect 2796 403 2821 406
rect 2852 403 2900 406
rect 2922 403 2932 406
rect 3148 403 3157 406
rect 3180 403 3221 406
rect 3266 403 3269 413
rect 4338 406 4341 413
rect 3298 403 3388 406
rect 3410 403 3428 406
rect 3946 403 3956 406
rect 3970 403 3996 406
rect 4180 403 4189 406
rect 4194 403 4212 406
rect 4244 403 4277 406
rect 4300 403 4341 406
rect 4586 403 4596 406
rect 4628 403 4645 406
rect 38 367 4837 373
rect 930 336 933 346
rect 3028 343 3077 346
rect 268 333 317 336
rect 380 333 389 336
rect 676 333 692 336
rect 738 333 764 336
rect 882 333 908 336
rect 930 333 956 336
rect 972 333 989 336
rect 1138 333 1148 336
rect 1194 333 1204 336
rect 1290 333 1300 336
rect 1626 333 1644 336
rect 930 326 933 333
rect 1778 326 1781 335
rect 1794 333 1820 336
rect 1852 333 1877 336
rect 1898 333 1916 336
rect 1970 333 1980 336
rect 2170 333 2196 336
rect 2492 333 2501 336
rect 2652 333 2661 336
rect 2674 333 2692 336
rect 2708 333 2725 336
rect 2730 333 2756 336
rect 2780 333 2797 336
rect 2828 333 2868 336
rect 2890 333 2900 336
rect 3020 333 3029 336
rect 3116 333 3164 336
rect 3180 333 3204 336
rect 3226 333 3260 336
rect 3410 333 3452 336
rect 3562 333 3580 336
rect 3596 333 3644 336
rect 3660 333 3677 336
rect 3706 333 3740 336
rect 3788 333 3797 336
rect 3826 333 3852 336
rect 3874 333 3884 336
rect 3898 333 3924 336
rect 3938 333 3948 336
rect 3964 333 3973 336
rect 1898 326 1901 333
rect 130 323 140 326
rect 274 323 356 326
rect 386 323 396 326
rect 460 323 485 326
rect 516 323 533 326
rect 572 323 597 326
rect 730 323 756 326
rect 916 323 933 326
rect 938 323 948 326
rect 1172 323 1212 326
rect 1226 323 1293 326
rect 1324 323 1380 326
rect 1460 323 1485 326
rect 1516 323 1525 326
rect 1564 323 1589 326
rect 1716 323 1733 326
rect 1772 323 1781 326
rect 1850 323 1901 326
rect 1940 323 1965 326
rect 1978 323 1988 326
rect 2164 323 2189 326
rect 2234 323 2244 326
rect 2420 323 2445 326
rect 2556 323 2581 326
rect 2612 323 2621 326
rect 2716 323 2733 326
rect 2738 323 2764 326
rect 2730 316 2733 323
rect 2794 316 2797 333
rect 2826 323 2860 326
rect 2892 323 2901 326
rect 2946 323 2972 326
rect 3138 323 3141 333
rect 3146 323 3156 326
rect 3370 323 3380 326
rect 3412 323 3421 326
rect 3498 323 3524 326
rect 3604 323 3629 326
rect 3730 323 3748 326
rect 3828 323 3837 326
rect 3882 323 3892 326
rect 3898 323 3932 326
rect 4010 325 4013 336
rect 4036 333 4061 336
rect 4170 333 4180 336
rect 4196 333 4220 336
rect 4244 333 4261 336
rect 4284 333 4300 336
rect 4444 333 4453 336
rect 4468 333 4485 336
rect 4522 333 4532 336
rect 4564 333 4573 336
rect 4594 333 4612 336
rect 4634 333 4684 336
rect 4108 323 4133 326
rect 4218 323 4228 326
rect 4442 323 4460 326
rect 4466 323 4484 326
rect 4530 323 4540 326
rect 4578 323 4604 326
rect 794 313 836 316
rect 860 313 893 316
rect 2730 313 2749 316
rect 2794 313 2804 316
rect 3834 293 3837 323
rect 14 267 4861 273
rect 2516 223 2525 226
rect 196 213 221 216
rect 252 213 261 216
rect 348 213 365 216
rect 516 213 541 216
rect 572 213 581 216
rect 588 213 597 216
rect 604 213 637 216
rect 756 213 788 216
rect 826 213 852 216
rect 922 213 940 216
rect 1036 213 1045 216
rect 1090 213 1100 216
rect 1242 213 1252 216
rect 1450 213 1476 216
rect 1636 213 1645 216
rect 1682 213 1748 216
rect 1778 213 1788 216
rect 1828 213 1837 216
rect 1900 213 1917 216
rect 2092 213 2117 216
rect 2148 213 2157 216
rect 2194 213 2204 216
rect 2210 213 2244 216
rect 2274 213 2292 216
rect 2332 213 2357 216
rect 2388 213 2397 216
rect 2404 213 2421 216
rect 258 205 261 213
rect 410 203 468 206
rect 578 205 581 213
rect 826 206 829 213
rect 676 203 709 206
rect 786 203 796 206
rect 812 203 829 206
rect 834 203 844 206
rect 994 203 1012 206
rect 1044 203 1061 206
rect 1522 203 1532 206
rect 1564 203 1589 206
rect 1612 203 1621 206
rect 1676 203 1693 206
rect 1914 203 1924 206
rect 2274 203 2284 206
rect 2394 205 2397 213
rect 2522 206 2525 223
rect 2556 213 2597 216
rect 2690 213 2733 216
rect 2738 213 2748 216
rect 2770 213 2780 216
rect 2858 213 2868 216
rect 2906 213 2932 216
rect 2970 213 2988 216
rect 3084 213 3109 216
rect 3154 213 3188 216
rect 3220 213 3228 216
rect 3594 213 3604 216
rect 3796 213 3805 216
rect 3930 213 3948 216
rect 4116 213 4140 216
rect 4172 213 4181 216
rect 4228 213 4237 216
rect 4298 213 4308 216
rect 4388 213 4413 216
rect 4498 213 4508 216
rect 4578 213 4596 216
rect 4668 213 4677 216
rect 2460 203 2477 206
rect 2482 203 2492 206
rect 2522 203 2540 206
rect 2570 203 2604 206
rect 2642 203 2652 206
rect 2698 203 2708 206
rect 2722 203 2740 206
rect 2796 203 2805 206
rect 2810 203 2820 206
rect 2826 203 2836 206
rect 2860 203 2876 206
rect 2962 203 2980 206
rect 3004 203 3013 206
rect 3156 203 3173 206
rect 3178 203 3196 206
rect 3212 203 3221 206
rect 3258 203 3268 206
rect 3300 203 3309 206
rect 3354 203 3372 206
rect 3394 203 3404 206
rect 3418 203 3428 206
rect 3450 203 3484 206
rect 4076 203 4085 206
rect 4130 203 4148 206
rect 4170 203 4180 206
rect 4290 203 4316 206
rect 4498 203 4516 206
rect 4538 203 4548 206
rect 4586 203 4604 206
rect 4666 203 4692 206
rect 38 167 4837 173
rect 690 133 708 136
rect 762 133 788 136
rect 1034 126 1037 135
rect 1186 126 1189 135
rect 1362 126 1365 135
rect 1506 126 1509 135
rect 2194 126 2197 136
rect 2466 133 2476 136
rect 2626 126 2629 135
rect 2642 133 2660 136
rect 2794 126 2797 135
rect 2954 133 2972 136
rect 354 123 380 126
rect 460 123 485 126
rect 516 123 533 126
rect 572 123 597 126
rect 628 123 645 126
rect 748 123 796 126
rect 866 123 892 126
rect 972 123 997 126
rect 1028 123 1037 126
rect 1108 123 1133 126
rect 1164 123 1189 126
rect 1284 123 1309 126
rect 1340 123 1365 126
rect 1444 123 1469 126
rect 1500 123 1509 126
rect 1516 123 1541 126
rect 1580 123 1605 126
rect 1708 123 1733 126
rect 1764 123 1781 126
rect 1820 123 1845 126
rect 1876 123 1893 126
rect 1932 123 1949 126
rect 2034 123 2044 126
rect 2116 123 2141 126
rect 2172 123 2197 126
rect 2250 123 2268 126
rect 2356 123 2381 126
rect 2412 123 2421 126
rect 2466 123 2501 126
rect 2540 123 2565 126
rect 2596 123 2629 126
rect 2658 123 2668 126
rect 2788 123 2797 126
rect 2890 123 2916 126
rect 3148 123 3173 126
rect 3210 123 3220 126
rect 3370 123 3380 126
rect 3410 123 3436 126
rect 3474 123 3492 126
rect 3522 123 3548 126
rect 3700 123 3717 126
rect 3722 123 3756 126
rect 3802 123 3812 126
rect 3924 123 3933 126
rect 4044 123 4069 126
rect 4100 123 4109 126
rect 4260 123 4285 126
rect 4322 123 4332 126
rect 4396 123 4421 126
rect 4458 123 4476 126
rect 14 67 4861 73
rect 38 37 4837 57
rect 14 13 4861 33
<< metal2 >>
rect 2 883 5 3536
rect 14 13 34 4727
rect 38 37 58 4703
rect 274 4636 277 4740
rect 274 4633 285 4636
rect 66 4533 69 4616
rect 138 4596 141 4616
rect 138 4593 149 4596
rect 130 4533 133 4546
rect 146 4533 149 4593
rect 74 4373 77 4416
rect 114 4333 117 4526
rect 154 4503 157 4526
rect 162 4496 165 4606
rect 202 4593 205 4606
rect 250 4603 253 4616
rect 282 4613 285 4633
rect 186 4533 189 4566
rect 226 4536 229 4566
rect 226 4533 237 4536
rect 274 4533 277 4546
rect 290 4533 293 4606
rect 306 4576 309 4616
rect 298 4573 309 4576
rect 154 4493 165 4496
rect 210 4496 213 4526
rect 210 4493 221 4496
rect 130 4343 133 4416
rect 66 4306 69 4326
rect 130 4313 133 4326
rect 66 4303 77 4306
rect 74 4236 77 4303
rect 154 4276 157 4493
rect 170 4373 173 4406
rect 178 4376 181 4416
rect 194 4393 197 4406
rect 178 4373 189 4376
rect 170 4296 173 4356
rect 178 4323 181 4373
rect 186 4333 189 4346
rect 66 4233 77 4236
rect 146 4273 157 4276
rect 162 4293 173 4296
rect 66 4203 69 4233
rect 146 4186 149 4273
rect 162 4193 165 4293
rect 170 4213 173 4226
rect 178 4203 181 4316
rect 186 4213 189 4246
rect 146 4183 157 4186
rect 66 4123 69 4136
rect 130 4123 133 4146
rect 74 3963 77 4016
rect 130 3993 133 4016
rect 154 3986 157 4183
rect 170 4133 181 4136
rect 186 4116 189 4196
rect 194 4176 197 4326
rect 202 4316 205 4336
rect 218 4333 221 4493
rect 234 4466 237 4533
rect 282 4493 285 4526
rect 298 4523 301 4573
rect 306 4533 309 4566
rect 226 4463 237 4466
rect 226 4353 229 4463
rect 306 4446 309 4526
rect 298 4443 309 4446
rect 242 4413 245 4426
rect 298 4413 301 4443
rect 202 4313 213 4316
rect 210 4226 213 4313
rect 202 4223 213 4226
rect 202 4193 205 4223
rect 234 4203 237 4396
rect 314 4393 317 4596
rect 354 4593 357 4606
rect 402 4603 405 4616
rect 322 4523 325 4536
rect 338 4423 341 4536
rect 346 4416 349 4536
rect 394 4516 397 4536
rect 434 4533 437 4606
rect 394 4513 405 4516
rect 378 4456 381 4506
rect 378 4453 385 4456
rect 338 4413 349 4416
rect 338 4346 341 4413
rect 362 4393 365 4416
rect 382 4346 385 4453
rect 402 4406 405 4513
rect 282 4323 285 4346
rect 330 4343 341 4346
rect 330 4256 333 4343
rect 330 4253 341 4256
rect 338 4236 341 4253
rect 194 4173 201 4176
rect 178 4113 189 4116
rect 178 4026 181 4113
rect 198 4106 201 4173
rect 210 4123 213 4136
rect 218 4133 221 4146
rect 194 4103 201 4106
rect 226 4103 229 4126
rect 194 4036 197 4103
rect 194 4033 201 4036
rect 178 4023 189 4026
rect 154 3983 165 3986
rect 162 3966 165 3983
rect 154 3963 165 3966
rect 170 3963 173 4006
rect 186 3963 189 4023
rect 198 3976 201 4033
rect 210 4013 213 4026
rect 218 3993 221 4006
rect 194 3973 201 3976
rect 82 3826 85 3946
rect 130 3913 133 3926
rect 154 3866 157 3963
rect 154 3863 165 3866
rect 82 3823 93 3826
rect 82 3733 85 3816
rect 90 3766 93 3823
rect 138 3803 141 3816
rect 90 3763 109 3766
rect 106 3656 109 3763
rect 82 3653 109 3656
rect 82 3486 85 3653
rect 130 3613 133 3626
rect 162 3533 165 3863
rect 170 3833 173 3956
rect 194 3953 197 3973
rect 194 3933 197 3946
rect 178 3813 181 3926
rect 186 3776 189 3836
rect 178 3773 189 3776
rect 178 3536 181 3773
rect 194 3646 197 3806
rect 202 3723 205 3736
rect 210 3733 213 3806
rect 218 3803 221 3916
rect 226 3906 229 4036
rect 234 4003 237 4196
rect 242 4023 245 4136
rect 250 3983 253 4126
rect 242 3923 245 3946
rect 258 3936 261 4106
rect 266 3953 269 4216
rect 282 4193 285 4216
rect 314 4123 317 4146
rect 330 4076 333 4236
rect 338 4233 345 4236
rect 326 4073 333 4076
rect 258 3933 265 3936
rect 226 3903 237 3906
rect 234 3846 237 3903
rect 262 3886 265 3933
rect 274 3923 277 4026
rect 298 3993 301 4006
rect 326 3986 329 4073
rect 342 4066 345 4233
rect 354 4136 357 4336
rect 370 4333 373 4346
rect 378 4343 385 4346
rect 394 4403 405 4406
rect 362 4323 373 4326
rect 370 4226 373 4246
rect 378 4233 381 4343
rect 394 4333 397 4403
rect 426 4336 429 4526
rect 402 4313 405 4336
rect 426 4333 437 4336
rect 426 4306 429 4326
rect 418 4303 429 4306
rect 394 4276 397 4296
rect 394 4273 405 4276
rect 370 4223 381 4226
rect 362 4203 365 4216
rect 370 4193 373 4206
rect 378 4183 381 4223
rect 402 4176 405 4273
rect 418 4226 421 4303
rect 434 4236 437 4333
rect 450 4313 453 4536
rect 458 4523 461 4616
rect 466 4533 469 4546
rect 458 4413 469 4416
rect 466 4393 469 4406
rect 474 4353 477 4636
rect 546 4623 549 4740
rect 730 4737 749 4740
rect 482 4463 485 4536
rect 490 4533 493 4606
rect 506 4583 509 4616
rect 530 4603 533 4616
rect 586 4613 589 4626
rect 594 4576 597 4596
rect 506 4533 509 4576
rect 590 4573 597 4576
rect 482 4383 485 4406
rect 474 4333 477 4346
rect 466 4303 469 4326
rect 434 4233 441 4236
rect 418 4223 429 4226
rect 394 4173 405 4176
rect 394 4156 397 4173
rect 386 4153 397 4156
rect 354 4133 373 4136
rect 226 3843 237 3846
rect 258 3883 265 3886
rect 226 3823 229 3843
rect 258 3836 261 3883
rect 282 3836 285 3936
rect 290 3923 293 3986
rect 322 3983 329 3986
rect 338 4063 345 4066
rect 298 3933 301 3946
rect 306 3856 309 3926
rect 322 3896 325 3983
rect 322 3893 333 3896
rect 322 3856 325 3876
rect 306 3853 325 3856
rect 258 3833 269 3836
rect 250 3816 253 3826
rect 226 3813 253 3816
rect 226 3796 229 3806
rect 218 3793 229 3796
rect 218 3723 221 3793
rect 234 3736 237 3806
rect 226 3733 237 3736
rect 242 3733 245 3756
rect 190 3643 197 3646
rect 190 3556 193 3643
rect 202 3613 205 3636
rect 202 3586 205 3606
rect 202 3583 209 3586
rect 190 3553 197 3556
rect 178 3533 189 3536
rect 130 3513 133 3526
rect 82 3483 93 3486
rect 90 3263 93 3483
rect 130 3403 133 3416
rect 162 3413 165 3526
rect 162 3393 165 3406
rect 170 3403 173 3416
rect 178 3403 181 3516
rect 138 3323 141 3346
rect 66 933 69 3036
rect 82 2756 85 3206
rect 114 3036 117 3216
rect 146 3156 149 3286
rect 170 3256 173 3326
rect 162 3253 173 3256
rect 154 3196 157 3246
rect 162 3206 165 3253
rect 178 3243 181 3336
rect 186 3323 189 3533
rect 194 3333 197 3553
rect 206 3426 209 3583
rect 218 3493 221 3626
rect 226 3613 229 3726
rect 234 3723 237 3733
rect 242 3633 245 3726
rect 250 3723 253 3813
rect 266 3756 269 3833
rect 278 3833 285 3836
rect 278 3776 281 3833
rect 298 3793 301 3806
rect 278 3773 285 3776
rect 258 3753 269 3756
rect 282 3756 285 3773
rect 282 3753 293 3756
rect 258 3643 261 3753
rect 266 3623 269 3736
rect 282 3733 285 3746
rect 290 3733 293 3753
rect 322 3736 325 3853
rect 330 3823 333 3893
rect 306 3733 325 3736
rect 330 3733 333 3816
rect 274 3683 277 3726
rect 306 3656 309 3733
rect 322 3713 325 3726
rect 338 3693 341 4063
rect 346 4003 349 4016
rect 306 3653 317 3656
rect 242 3566 245 3606
rect 242 3563 253 3566
rect 250 3546 253 3563
rect 274 3556 277 3646
rect 290 3593 293 3616
rect 314 3556 317 3653
rect 346 3573 349 3936
rect 354 3933 357 3956
rect 362 3933 365 4133
rect 386 4106 389 4153
rect 410 4133 413 4146
rect 426 4133 429 4223
rect 438 4176 441 4233
rect 458 4203 461 4216
rect 438 4173 445 4176
rect 442 4126 445 4173
rect 402 4113 405 4126
rect 386 4103 397 4106
rect 370 3933 373 4006
rect 378 3966 381 4016
rect 394 3993 397 4103
rect 418 4033 421 4126
rect 434 4123 445 4126
rect 378 3963 397 3966
rect 386 3933 389 3946
rect 394 3933 397 3963
rect 362 3913 365 3926
rect 370 3896 373 3926
rect 366 3893 373 3896
rect 366 3726 369 3893
rect 378 3823 381 3926
rect 394 3913 397 3926
rect 402 3836 405 3966
rect 410 3926 413 3996
rect 418 3933 421 3946
rect 410 3923 421 3926
rect 394 3833 405 3836
rect 378 3733 381 3816
rect 394 3786 397 3833
rect 394 3783 405 3786
rect 354 3713 357 3726
rect 366 3723 373 3726
rect 270 3553 277 3556
rect 306 3553 317 3556
rect 234 3533 237 3546
rect 250 3543 261 3546
rect 202 3423 209 3426
rect 170 3223 189 3226
rect 170 3213 173 3223
rect 162 3203 173 3206
rect 178 3203 181 3216
rect 186 3203 189 3223
rect 154 3193 165 3196
rect 162 3176 165 3193
rect 162 3173 173 3176
rect 146 3153 157 3156
rect 114 3033 121 3036
rect 98 2813 101 2896
rect 106 2876 109 3026
rect 118 2966 121 3033
rect 114 2963 121 2966
rect 114 2893 117 2963
rect 106 2873 113 2876
rect 110 2806 113 2873
rect 78 2753 85 2756
rect 106 2803 113 2806
rect 78 2616 81 2753
rect 74 2613 81 2616
rect 74 2563 77 2613
rect 74 2256 77 2556
rect 82 2523 85 2606
rect 90 2583 93 2746
rect 98 2603 101 2616
rect 98 2523 101 2536
rect 82 2496 85 2516
rect 106 2506 109 2803
rect 122 2783 125 2926
rect 130 2743 133 3126
rect 154 3086 157 3153
rect 146 3083 157 3086
rect 146 3013 149 3083
rect 170 3006 173 3173
rect 194 3123 197 3326
rect 202 3283 205 3423
rect 210 3373 213 3406
rect 226 3403 229 3426
rect 210 3203 213 3326
rect 218 3103 221 3386
rect 250 3383 253 3496
rect 258 3423 261 3543
rect 270 3436 273 3553
rect 282 3523 285 3546
rect 266 3433 273 3436
rect 234 3113 237 3136
rect 242 3133 245 3336
rect 258 3333 261 3346
rect 250 3313 253 3326
rect 266 3213 269 3433
rect 306 3426 309 3553
rect 298 3423 309 3426
rect 274 3393 277 3416
rect 274 3333 277 3376
rect 298 3346 301 3423
rect 298 3343 309 3346
rect 306 3323 309 3343
rect 314 3333 317 3416
rect 322 3403 325 3526
rect 330 3523 333 3536
rect 338 3506 341 3526
rect 338 3503 349 3506
rect 346 3436 349 3503
rect 338 3433 349 3436
rect 338 3413 341 3433
rect 354 3323 357 3416
rect 362 3306 365 3416
rect 370 3386 373 3723
rect 394 3706 397 3726
rect 386 3703 397 3706
rect 386 3646 389 3703
rect 402 3656 405 3783
rect 418 3723 421 3923
rect 434 3846 437 4123
rect 442 4003 445 4016
rect 450 3883 453 3936
rect 458 3873 461 4186
rect 482 4133 485 4216
rect 490 4206 493 4336
rect 498 4323 501 4416
rect 506 4323 509 4406
rect 522 4403 525 4536
rect 530 4523 533 4546
rect 538 4483 541 4526
rect 546 4503 549 4536
rect 554 4493 557 4526
rect 546 4413 549 4436
rect 554 4416 557 4446
rect 562 4423 565 4556
rect 570 4416 573 4536
rect 590 4526 593 4573
rect 602 4533 605 4556
rect 618 4533 621 4616
rect 578 4483 581 4526
rect 590 4523 597 4526
rect 554 4413 565 4416
rect 570 4413 581 4416
rect 586 4413 589 4436
rect 554 4383 557 4406
rect 562 4403 573 4406
rect 578 4403 581 4413
rect 594 4396 597 4523
rect 610 4476 613 4526
rect 586 4393 597 4396
rect 606 4473 613 4476
rect 522 4336 525 4356
rect 518 4333 525 4336
rect 518 4276 521 4333
rect 538 4323 541 4346
rect 586 4293 589 4393
rect 606 4356 609 4473
rect 606 4353 613 4356
rect 602 4323 605 4336
rect 610 4313 613 4353
rect 518 4273 525 4276
rect 522 4256 525 4273
rect 522 4253 533 4256
rect 490 4203 501 4206
rect 498 4133 501 4203
rect 530 4196 533 4253
rect 522 4193 533 4196
rect 522 4176 525 4193
rect 518 4173 525 4176
rect 474 4103 477 4126
rect 506 4113 509 4136
rect 518 4106 521 4173
rect 554 4166 557 4216
rect 578 4193 581 4206
rect 538 4163 557 4166
rect 538 4123 541 4163
rect 554 4133 557 4156
rect 514 4103 521 4106
rect 466 3933 469 4006
rect 482 3933 485 3956
rect 490 3923 493 4016
rect 506 3916 509 3936
rect 502 3913 509 3916
rect 434 3843 445 3846
rect 442 3746 445 3843
rect 458 3813 461 3826
rect 490 3776 493 3846
rect 502 3826 505 3913
rect 502 3823 509 3826
rect 486 3773 493 3776
rect 442 3743 453 3746
rect 450 3696 453 3743
rect 466 3723 469 3746
rect 434 3693 453 3696
rect 402 3653 421 3656
rect 386 3643 397 3646
rect 378 3613 381 3626
rect 394 3583 397 3643
rect 386 3533 389 3546
rect 378 3513 381 3526
rect 394 3523 397 3536
rect 378 3393 381 3406
rect 370 3383 377 3386
rect 354 3303 365 3306
rect 374 3306 377 3383
rect 386 3316 389 3446
rect 402 3373 405 3576
rect 410 3333 413 3406
rect 418 3383 421 3653
rect 426 3516 429 3536
rect 434 3533 437 3693
rect 486 3626 489 3773
rect 506 3766 509 3823
rect 498 3763 509 3766
rect 486 3623 493 3626
rect 442 3603 445 3616
rect 466 3533 469 3546
rect 426 3513 437 3516
rect 434 3446 437 3513
rect 474 3483 477 3536
rect 482 3533 485 3606
rect 490 3516 493 3623
rect 486 3513 493 3516
rect 426 3443 437 3446
rect 426 3413 429 3443
rect 434 3403 437 3416
rect 434 3333 437 3396
rect 386 3313 397 3316
rect 374 3303 381 3306
rect 354 3236 357 3303
rect 354 3233 365 3236
rect 274 3193 277 3206
rect 242 3113 245 3126
rect 282 3123 285 3216
rect 314 3213 317 3226
rect 290 3193 293 3206
rect 298 3133 301 3156
rect 306 3123 309 3136
rect 274 3103 277 3116
rect 162 3003 173 3006
rect 146 2816 149 2936
rect 162 2923 165 3003
rect 170 2906 173 2936
rect 178 2923 181 2946
rect 186 2923 189 2936
rect 202 2916 205 2926
rect 142 2813 149 2816
rect 162 2903 173 2906
rect 162 2816 165 2903
rect 162 2813 173 2816
rect 178 2813 181 2916
rect 186 2913 205 2916
rect 142 2736 145 2813
rect 138 2733 145 2736
rect 138 2713 141 2733
rect 154 2703 157 2796
rect 170 2756 173 2813
rect 162 2753 173 2756
rect 162 2686 165 2753
rect 170 2713 173 2746
rect 178 2706 181 2806
rect 154 2683 165 2686
rect 170 2703 181 2706
rect 186 2703 189 2846
rect 202 2796 205 2816
rect 202 2793 209 2796
rect 114 2546 117 2566
rect 114 2543 121 2546
rect 102 2503 109 2506
rect 82 2493 93 2496
rect 90 2426 93 2493
rect 82 2423 93 2426
rect 82 2273 85 2423
rect 102 2406 105 2503
rect 118 2496 121 2543
rect 114 2493 121 2496
rect 114 2413 117 2493
rect 130 2416 133 2676
rect 154 2616 157 2683
rect 170 2626 173 2703
rect 170 2623 181 2626
rect 154 2613 165 2616
rect 138 2543 141 2596
rect 130 2413 137 2416
rect 90 2313 93 2406
rect 102 2403 109 2406
rect 106 2336 109 2403
rect 102 2333 109 2336
rect 74 2253 81 2256
rect 78 2096 81 2253
rect 102 2236 105 2333
rect 102 2233 109 2236
rect 90 2113 93 2206
rect 98 2173 101 2216
rect 106 2213 109 2233
rect 114 2213 117 2326
rect 122 2323 125 2406
rect 134 2336 137 2413
rect 154 2396 157 2546
rect 162 2523 165 2613
rect 178 2566 181 2623
rect 170 2563 181 2566
rect 170 2496 173 2563
rect 194 2553 197 2786
rect 206 2646 209 2793
rect 202 2643 209 2646
rect 202 2623 205 2643
rect 218 2593 221 3016
rect 242 2943 245 2956
rect 266 2943 269 3006
rect 258 2843 261 2936
rect 282 2926 285 3116
rect 314 3106 317 3136
rect 306 3103 317 3106
rect 306 3036 309 3103
rect 306 3033 317 3036
rect 314 2946 317 3033
rect 322 3003 325 3196
rect 330 3153 333 3226
rect 362 3216 365 3233
rect 338 3203 341 3216
rect 362 3213 373 3216
rect 330 3096 333 3116
rect 330 3093 337 3096
rect 334 3026 337 3093
rect 330 3023 337 3026
rect 346 3023 349 3166
rect 354 3133 357 3206
rect 330 2966 333 3023
rect 306 2943 317 2946
rect 322 2963 333 2966
rect 274 2923 285 2926
rect 274 2846 277 2923
rect 274 2843 285 2846
rect 250 2803 253 2816
rect 258 2803 261 2836
rect 274 2813 277 2826
rect 266 2796 269 2806
rect 226 2573 229 2796
rect 242 2793 269 2796
rect 234 2716 237 2736
rect 234 2713 245 2716
rect 242 2646 245 2713
rect 282 2673 285 2843
rect 290 2793 293 2936
rect 298 2813 301 2826
rect 234 2643 245 2646
rect 234 2613 237 2643
rect 306 2633 309 2943
rect 314 2923 317 2936
rect 322 2933 325 2963
rect 338 2933 341 2956
rect 322 2833 325 2926
rect 346 2923 349 3016
rect 354 2983 357 3006
rect 362 2993 365 3206
rect 370 3196 373 3213
rect 378 3203 381 3303
rect 394 3256 397 3313
rect 386 3253 397 3256
rect 426 3253 429 3326
rect 442 3316 445 3386
rect 450 3373 453 3426
rect 474 3393 477 3416
rect 486 3406 489 3513
rect 498 3413 501 3763
rect 514 3683 517 4103
rect 538 3993 541 4006
rect 522 3913 525 3936
rect 546 3873 549 4126
rect 562 4106 565 4166
rect 558 4103 565 4106
rect 558 4036 561 4103
rect 558 4033 565 4036
rect 554 4003 557 4016
rect 554 3933 557 3946
rect 562 3923 565 4033
rect 570 4023 573 4136
rect 578 4113 581 4136
rect 586 4103 589 4286
rect 618 4283 621 4486
rect 634 4466 637 4536
rect 642 4533 645 4546
rect 650 4473 653 4606
rect 666 4603 669 4616
rect 658 4533 661 4586
rect 690 4583 693 4616
rect 746 4613 749 4737
rect 1994 4683 2005 4686
rect 762 4586 765 4616
rect 762 4583 773 4586
rect 674 4533 677 4576
rect 682 4533 685 4566
rect 634 4463 645 4466
rect 626 4403 629 4436
rect 634 4413 637 4446
rect 642 4403 645 4463
rect 666 4426 669 4446
rect 650 4413 653 4426
rect 662 4423 669 4426
rect 650 4393 653 4406
rect 626 4333 629 4356
rect 634 4333 645 4336
rect 594 4203 597 4216
rect 602 4163 605 4246
rect 634 4243 637 4326
rect 650 4323 653 4336
rect 662 4306 665 4423
rect 658 4303 665 4306
rect 658 4236 661 4303
rect 610 4203 613 4226
rect 618 4193 621 4206
rect 626 4186 629 4236
rect 658 4233 669 4236
rect 674 4233 677 4416
rect 690 4403 693 4416
rect 698 4413 701 4446
rect 706 4373 709 4406
rect 714 4403 717 4536
rect 738 4533 741 4546
rect 754 4526 757 4536
rect 770 4533 773 4583
rect 778 4573 781 4606
rect 826 4593 829 4616
rect 778 4533 781 4546
rect 722 4513 725 4526
rect 730 4483 733 4526
rect 746 4493 749 4526
rect 754 4523 765 4526
rect 810 4523 821 4526
rect 762 4456 765 4523
rect 754 4453 765 4456
rect 722 4413 725 4426
rect 746 4413 749 4446
rect 714 4376 717 4396
rect 738 4393 741 4406
rect 754 4403 757 4453
rect 770 4413 773 4426
rect 818 4406 821 4446
rect 762 4393 765 4406
rect 714 4373 725 4376
rect 682 4333 685 4346
rect 690 4333 701 4336
rect 706 4333 709 4346
rect 722 4326 725 4373
rect 618 4183 629 4186
rect 570 3983 573 4006
rect 578 3993 581 4006
rect 570 3903 573 3936
rect 578 3913 581 3936
rect 522 3793 525 3816
rect 538 3813 541 3836
rect 530 3733 533 3806
rect 546 3803 549 3826
rect 554 3763 557 3816
rect 546 3733 549 3746
rect 538 3723 549 3726
rect 554 3693 557 3726
rect 506 3533 509 3616
rect 514 3613 517 3626
rect 522 3576 525 3636
rect 538 3593 541 3606
rect 546 3603 549 3686
rect 562 3676 565 3886
rect 618 3836 621 4183
rect 626 4073 629 4136
rect 634 4076 637 4206
rect 658 4193 661 4206
rect 666 4203 669 4233
rect 674 4203 677 4226
rect 690 4203 693 4326
rect 714 4323 725 4326
rect 642 4123 645 4136
rect 650 4133 653 4146
rect 650 4103 653 4126
rect 682 4116 685 4136
rect 698 4123 701 4216
rect 714 4203 717 4323
rect 730 4203 733 4226
rect 706 4133 709 4176
rect 714 4133 725 4136
rect 706 4123 717 4126
rect 674 4113 685 4116
rect 634 4073 645 4076
rect 634 3983 637 4006
rect 642 3946 645 4073
rect 674 4046 677 4113
rect 674 4043 685 4046
rect 658 4013 661 4026
rect 650 3993 653 4006
rect 682 4003 685 4043
rect 698 4003 701 4116
rect 714 4106 717 4123
rect 710 4103 717 4106
rect 710 4036 713 4103
rect 710 4033 717 4036
rect 706 4003 709 4016
rect 634 3943 645 3946
rect 626 3923 629 3936
rect 634 3876 637 3943
rect 642 3903 645 3936
rect 634 3873 645 3876
rect 570 3813 573 3836
rect 618 3833 629 3836
rect 570 3793 573 3806
rect 570 3703 573 3736
rect 610 3706 613 3746
rect 594 3703 613 3706
rect 554 3673 565 3676
rect 522 3573 533 3576
rect 530 3526 533 3573
rect 554 3543 557 3673
rect 594 3566 597 3703
rect 618 3686 621 3736
rect 610 3683 621 3686
rect 610 3636 613 3683
rect 610 3633 621 3636
rect 618 3613 621 3633
rect 594 3563 613 3566
rect 522 3523 533 3526
rect 486 3403 493 3406
rect 450 3333 453 3356
rect 442 3313 453 3316
rect 386 3233 389 3253
rect 370 3193 381 3196
rect 370 3126 373 3176
rect 378 3133 381 3193
rect 386 3173 389 3226
rect 402 3213 421 3216
rect 386 3133 389 3146
rect 370 3123 381 3126
rect 394 3123 397 3206
rect 426 3173 429 3226
rect 434 3133 437 3266
rect 450 3226 453 3313
rect 490 3226 493 3403
rect 442 3223 453 3226
rect 442 3203 445 3223
rect 474 3213 477 3226
rect 490 3223 509 3226
rect 450 3136 453 3206
rect 450 3133 461 3136
rect 466 3133 469 3166
rect 442 3123 453 3126
rect 378 3113 381 3123
rect 442 3033 445 3123
rect 458 3103 461 3133
rect 314 2803 317 2826
rect 330 2746 333 2816
rect 322 2743 333 2746
rect 322 2693 325 2743
rect 330 2723 333 2736
rect 338 2733 341 2746
rect 346 2726 349 2746
rect 370 2743 373 3016
rect 434 2976 437 2996
rect 426 2973 437 2976
rect 394 2813 397 2936
rect 426 2836 429 2973
rect 450 2836 453 2986
rect 458 2933 461 2996
rect 474 2956 477 3196
rect 482 3133 485 3206
rect 490 3023 493 3216
rect 506 3136 509 3223
rect 522 3193 525 3523
rect 586 3506 589 3526
rect 594 3523 597 3536
rect 602 3533 605 3546
rect 602 3506 605 3526
rect 578 3503 589 3506
rect 598 3503 605 3506
rect 578 3426 581 3503
rect 578 3423 589 3426
rect 530 3333 533 3416
rect 546 3236 549 3326
rect 554 3323 557 3416
rect 586 3403 589 3423
rect 562 3323 565 3336
rect 570 3323 573 3336
rect 578 3313 581 3336
rect 586 3333 589 3346
rect 598 3316 601 3503
rect 598 3313 605 3316
rect 578 3236 581 3306
rect 546 3233 565 3236
rect 578 3233 585 3236
rect 562 3203 565 3233
rect 570 3173 573 3226
rect 582 3166 585 3233
rect 522 3146 525 3166
rect 578 3163 585 3166
rect 522 3143 529 3146
rect 502 3133 509 3136
rect 502 3026 505 3133
rect 514 3103 517 3116
rect 526 3096 529 3143
rect 538 3133 557 3136
rect 498 3023 505 3026
rect 522 3093 529 3096
rect 498 2983 501 3023
rect 506 2993 509 3006
rect 522 3003 525 3093
rect 554 3026 557 3133
rect 538 3013 541 3026
rect 554 3023 565 3026
rect 470 2953 477 2956
rect 562 2953 565 3023
rect 578 3006 581 3163
rect 578 3003 585 3006
rect 470 2906 473 2953
rect 482 2923 485 2946
rect 570 2923 573 2996
rect 582 2946 585 3003
rect 578 2943 585 2946
rect 470 2903 477 2906
rect 426 2833 437 2836
rect 450 2833 461 2836
rect 434 2813 437 2833
rect 442 2813 445 2826
rect 338 2723 349 2726
rect 410 2723 413 2796
rect 442 2783 445 2796
rect 338 2626 341 2723
rect 434 2713 437 2726
rect 354 2633 357 2696
rect 338 2623 357 2626
rect 242 2593 245 2606
rect 178 2533 181 2546
rect 186 2533 189 2546
rect 274 2496 277 2526
rect 170 2493 181 2496
rect 178 2426 181 2493
rect 266 2493 277 2496
rect 170 2423 181 2426
rect 130 2333 137 2336
rect 146 2393 157 2396
rect 106 2203 117 2206
rect 106 2166 109 2203
rect 102 2163 109 2166
rect 102 2106 105 2163
rect 122 2146 125 2306
rect 130 2166 133 2333
rect 138 2303 141 2316
rect 138 2203 141 2226
rect 146 2183 149 2393
rect 154 2313 157 2326
rect 162 2226 165 2406
rect 170 2403 173 2423
rect 202 2413 205 2456
rect 266 2426 269 2493
rect 282 2436 285 2536
rect 290 2533 293 2576
rect 298 2513 301 2586
rect 282 2433 289 2436
rect 266 2423 277 2426
rect 194 2333 197 2346
rect 202 2343 205 2396
rect 266 2393 269 2406
rect 274 2343 277 2423
rect 286 2356 289 2433
rect 298 2413 301 2446
rect 286 2353 301 2356
rect 170 2233 173 2306
rect 178 2293 181 2326
rect 290 2316 293 2326
rect 298 2323 301 2353
rect 162 2223 181 2226
rect 186 2216 189 2316
rect 290 2313 301 2316
rect 162 2213 189 2216
rect 130 2163 141 2166
rect 98 2103 105 2106
rect 78 2093 85 2096
rect 82 1966 85 2093
rect 74 1963 85 1966
rect 74 1896 77 1963
rect 98 1953 101 2103
rect 114 1996 117 2146
rect 122 2143 129 2146
rect 126 2036 129 2143
rect 122 2033 129 2036
rect 122 2013 125 2033
rect 114 1993 125 1996
rect 122 1933 125 1993
rect 138 1946 141 2163
rect 154 2123 173 2126
rect 154 2003 157 2106
rect 130 1943 141 1946
rect 74 1893 81 1896
rect 78 1816 81 1893
rect 90 1836 93 1926
rect 90 1833 109 1836
rect 98 1823 117 1826
rect 122 1823 125 1836
rect 78 1813 85 1816
rect 82 1756 85 1813
rect 78 1753 85 1756
rect 78 1446 81 1753
rect 98 1736 101 1806
rect 90 1733 101 1736
rect 90 1543 93 1733
rect 98 1706 101 1726
rect 98 1703 105 1706
rect 102 1626 105 1703
rect 98 1623 105 1626
rect 98 1593 101 1623
rect 106 1576 109 1606
rect 102 1573 109 1576
rect 74 1443 81 1446
rect 74 1386 77 1443
rect 74 1383 81 1386
rect 78 1226 81 1383
rect 78 1223 85 1226
rect 74 976 77 1206
rect 82 1183 85 1223
rect 74 973 81 976
rect 66 513 69 926
rect 78 836 81 973
rect 74 833 81 836
rect 74 813 77 833
rect 90 733 93 1526
rect 102 1516 105 1573
rect 114 1523 117 1823
rect 130 1806 133 1943
rect 154 1933 157 1956
rect 126 1803 133 1806
rect 126 1616 129 1803
rect 138 1623 141 1836
rect 146 1803 149 1926
rect 162 1846 165 2116
rect 170 2096 173 2123
rect 178 2113 181 2213
rect 186 2133 189 2146
rect 194 2126 197 2226
rect 202 2143 205 2306
rect 298 2303 301 2313
rect 234 2136 237 2156
rect 226 2133 237 2136
rect 242 2136 245 2236
rect 258 2213 261 2296
rect 266 2206 269 2256
rect 298 2223 301 2286
rect 306 2266 309 2616
rect 314 2403 317 2606
rect 330 2543 333 2616
rect 338 2533 341 2616
rect 322 2423 325 2526
rect 314 2286 317 2336
rect 322 2323 325 2406
rect 322 2293 325 2316
rect 314 2283 325 2286
rect 306 2263 313 2266
rect 310 2216 313 2263
rect 258 2203 269 2206
rect 250 2143 253 2156
rect 242 2133 253 2136
rect 186 2123 197 2126
rect 170 2093 177 2096
rect 174 2016 177 2093
rect 170 2013 177 2016
rect 170 1933 173 2013
rect 162 1843 173 1846
rect 154 1813 157 1836
rect 154 1736 157 1806
rect 170 1736 173 1843
rect 146 1733 157 1736
rect 162 1733 173 1736
rect 146 1703 149 1733
rect 162 1623 165 1733
rect 126 1613 133 1616
rect 130 1546 133 1613
rect 130 1543 141 1546
rect 102 1513 109 1516
rect 106 1446 109 1513
rect 106 1443 117 1446
rect 114 1406 117 1443
rect 122 1413 125 1536
rect 138 1466 141 1543
rect 162 1523 165 1536
rect 186 1523 189 2123
rect 210 1916 213 2126
rect 226 2016 229 2133
rect 242 2026 245 2126
rect 250 2106 253 2133
rect 258 2113 261 2203
rect 250 2103 261 2106
rect 242 2023 249 2026
rect 226 2013 237 2016
rect 218 1923 221 1936
rect 234 1933 237 2013
rect 246 1976 249 2023
rect 266 2013 269 2126
rect 282 2046 285 2106
rect 290 2093 293 2216
rect 306 2213 313 2216
rect 298 2113 301 2146
rect 278 2043 285 2046
rect 242 1973 249 1976
rect 210 1913 237 1916
rect 242 1816 245 1973
rect 250 1923 253 1956
rect 258 1903 261 2006
rect 278 1966 281 2043
rect 278 1963 285 1966
rect 274 1933 277 1946
rect 218 1803 221 1816
rect 242 1813 253 1816
rect 242 1793 245 1806
rect 218 1613 221 1626
rect 194 1586 197 1606
rect 226 1603 229 1786
rect 250 1636 253 1813
rect 266 1783 269 1926
rect 282 1913 285 1963
rect 290 1896 293 2036
rect 282 1893 293 1896
rect 282 1826 285 1893
rect 282 1823 293 1826
rect 290 1803 293 1823
rect 298 1803 301 1916
rect 282 1686 285 1736
rect 242 1633 253 1636
rect 266 1683 285 1686
rect 242 1586 245 1633
rect 194 1583 205 1586
rect 242 1583 257 1586
rect 202 1516 205 1583
rect 134 1463 141 1466
rect 194 1513 205 1516
rect 114 1403 121 1406
rect 98 1213 101 1346
rect 106 1333 109 1366
rect 118 1326 121 1403
rect 134 1396 137 1463
rect 194 1423 197 1513
rect 130 1393 137 1396
rect 130 1333 133 1393
rect 118 1323 125 1326
rect 98 1203 117 1206
rect 122 1176 125 1323
rect 154 1316 157 1346
rect 146 1313 157 1316
rect 146 1246 149 1313
rect 146 1243 157 1246
rect 154 1213 157 1243
rect 170 1203 173 1416
rect 178 1343 181 1406
rect 178 1303 181 1326
rect 186 1313 189 1416
rect 194 1323 197 1416
rect 218 1403 221 1436
rect 226 1396 229 1416
rect 234 1403 237 1416
rect 242 1413 245 1526
rect 254 1516 257 1583
rect 266 1523 269 1683
rect 306 1676 309 2213
rect 322 2193 325 2283
rect 330 2213 333 2506
rect 338 2413 341 2526
rect 338 2316 341 2406
rect 346 2403 349 2576
rect 354 2523 357 2623
rect 346 2333 349 2396
rect 354 2346 357 2516
rect 362 2453 365 2706
rect 370 2576 373 2616
rect 378 2593 381 2606
rect 370 2573 377 2576
rect 374 2446 377 2573
rect 386 2496 389 2596
rect 394 2563 397 2606
rect 410 2603 413 2636
rect 434 2573 437 2656
rect 442 2613 445 2776
rect 458 2756 461 2833
rect 474 2773 477 2903
rect 490 2803 509 2806
rect 450 2753 461 2756
rect 450 2733 453 2753
rect 450 2633 453 2726
rect 458 2713 461 2736
rect 474 2726 477 2746
rect 522 2733 525 2826
rect 578 2816 581 2943
rect 562 2813 581 2816
rect 586 2813 589 2826
rect 594 2813 597 3296
rect 602 3213 605 3313
rect 610 3243 613 3563
rect 618 3513 621 3536
rect 626 3533 629 3833
rect 634 3783 637 3806
rect 642 3743 645 3873
rect 634 3716 637 3736
rect 650 3733 653 3806
rect 658 3803 661 3836
rect 666 3786 669 3926
rect 662 3783 669 3786
rect 662 3716 665 3783
rect 634 3713 645 3716
rect 642 3646 645 3713
rect 634 3643 645 3646
rect 658 3713 665 3716
rect 634 3603 637 3643
rect 658 3626 661 3713
rect 650 3623 661 3626
rect 634 3516 637 3586
rect 650 3536 653 3623
rect 674 3616 677 3876
rect 690 3813 693 3936
rect 714 3813 717 4033
rect 722 4003 725 4133
rect 730 4113 733 4136
rect 738 4123 741 4246
rect 746 4203 749 4376
rect 786 4366 789 4406
rect 794 4383 797 4406
rect 814 4403 821 4406
rect 786 4363 805 4366
rect 770 4323 781 4326
rect 754 4193 757 4206
rect 762 4176 765 4256
rect 786 4253 789 4336
rect 794 4333 797 4356
rect 794 4246 797 4316
rect 754 4173 765 4176
rect 770 4243 797 4246
rect 754 4116 757 4173
rect 770 4133 773 4243
rect 778 4183 781 4216
rect 786 4163 789 4236
rect 794 4223 797 4243
rect 802 4233 805 4363
rect 814 4336 817 4403
rect 814 4333 821 4336
rect 770 4123 781 4126
rect 754 4113 765 4116
rect 746 4026 749 4046
rect 746 4023 753 4026
rect 730 3933 733 4006
rect 738 3916 741 4016
rect 750 3956 753 4023
rect 730 3913 741 3916
rect 746 3953 753 3956
rect 730 3836 733 3913
rect 730 3833 741 3836
rect 706 3793 709 3806
rect 714 3803 725 3806
rect 730 3803 733 3816
rect 714 3773 717 3803
rect 738 3786 741 3833
rect 734 3783 741 3786
rect 682 3723 685 3736
rect 698 3733 701 3756
rect 706 3723 709 3746
rect 714 3713 717 3736
rect 666 3613 677 3616
rect 650 3533 661 3536
rect 630 3513 637 3516
rect 630 3436 633 3513
rect 630 3433 637 3436
rect 618 3263 621 3426
rect 626 3393 629 3406
rect 634 3396 637 3433
rect 642 3403 645 3516
rect 650 3423 653 3516
rect 634 3393 645 3396
rect 634 3333 637 3356
rect 642 3326 645 3393
rect 650 3333 653 3406
rect 658 3356 661 3533
rect 666 3423 669 3613
rect 674 3593 677 3606
rect 682 3583 685 3626
rect 690 3603 693 3706
rect 698 3586 701 3606
rect 694 3583 701 3586
rect 658 3353 669 3356
rect 658 3333 661 3346
rect 642 3323 653 3326
rect 618 3213 621 3226
rect 634 3213 637 3246
rect 626 3193 629 3206
rect 642 3203 645 3316
rect 650 3213 653 3323
rect 658 3223 661 3326
rect 602 3133 613 3136
rect 610 3003 613 3133
rect 634 3016 637 3176
rect 658 3133 661 3146
rect 642 3023 645 3046
rect 650 3023 653 3126
rect 666 3066 669 3353
rect 674 3323 677 3536
rect 694 3516 697 3583
rect 706 3523 709 3606
rect 714 3523 717 3646
rect 722 3613 725 3766
rect 734 3656 737 3783
rect 734 3653 741 3656
rect 738 3633 741 3653
rect 746 3643 749 3953
rect 754 3796 757 3936
rect 762 3913 765 4113
rect 786 4106 789 4136
rect 778 4103 789 4106
rect 778 4036 781 4103
rect 778 4033 789 4036
rect 770 3856 773 3916
rect 762 3853 773 3856
rect 762 3813 765 3853
rect 778 3843 781 4016
rect 786 3933 789 4033
rect 794 4023 797 4206
rect 802 4203 805 4216
rect 802 4023 805 4136
rect 802 3933 805 3986
rect 786 3906 789 3926
rect 810 3913 813 4316
rect 818 4313 821 4333
rect 826 4226 829 4536
rect 834 4533 837 4556
rect 850 4453 853 4536
rect 874 4523 877 4586
rect 898 4563 901 4606
rect 906 4553 909 4616
rect 914 4593 917 4606
rect 922 4603 925 4616
rect 938 4603 941 4616
rect 954 4573 957 4626
rect 1002 4593 1005 4616
rect 1058 4563 1061 4606
rect 1090 4596 1093 4616
rect 1106 4613 1109 4636
rect 1082 4593 1093 4596
rect 1098 4593 1101 4606
rect 1114 4593 1117 4616
rect 882 4533 893 4536
rect 858 4513 893 4516
rect 850 4423 853 4446
rect 866 4416 869 4513
rect 834 4393 837 4416
rect 862 4413 869 4416
rect 862 4356 865 4413
rect 862 4353 869 4356
rect 834 4323 837 4336
rect 826 4223 833 4226
rect 818 4203 821 4216
rect 830 4166 833 4223
rect 818 3906 821 4166
rect 786 3903 797 3906
rect 794 3836 797 3903
rect 786 3833 797 3836
rect 810 3903 821 3906
rect 826 4163 833 4166
rect 754 3793 761 3796
rect 758 3716 761 3793
rect 754 3713 761 3716
rect 730 3623 749 3626
rect 694 3513 701 3516
rect 730 3513 733 3623
rect 754 3546 757 3713
rect 762 3613 765 3696
rect 770 3623 773 3826
rect 786 3803 789 3833
rect 794 3793 797 3806
rect 778 3733 781 3746
rect 786 3723 789 3736
rect 794 3723 797 3736
rect 802 3733 805 3746
rect 810 3726 813 3903
rect 818 3813 821 3836
rect 802 3723 813 3726
rect 786 3616 789 3636
rect 782 3613 789 3616
rect 802 3616 805 3723
rect 802 3613 809 3616
rect 746 3543 757 3546
rect 698 3496 701 3513
rect 746 3496 749 3543
rect 782 3536 785 3613
rect 698 3493 709 3496
rect 682 3413 685 3486
rect 706 3416 709 3493
rect 690 3413 709 3416
rect 738 3493 749 3496
rect 690 3313 693 3413
rect 698 3386 701 3406
rect 738 3386 741 3493
rect 762 3476 765 3536
rect 770 3516 773 3536
rect 782 3533 789 3536
rect 770 3513 777 3516
rect 754 3473 765 3476
rect 754 3406 757 3473
rect 774 3466 777 3513
rect 770 3463 777 3466
rect 754 3403 765 3406
rect 770 3403 773 3463
rect 762 3386 765 3403
rect 698 3383 705 3386
rect 738 3383 757 3386
rect 762 3383 769 3386
rect 702 3306 705 3383
rect 714 3333 717 3346
rect 730 3333 733 3366
rect 738 3333 741 3346
rect 698 3303 705 3306
rect 674 3266 677 3286
rect 674 3263 685 3266
rect 682 3166 685 3263
rect 674 3163 685 3166
rect 674 3143 677 3163
rect 698 3106 701 3303
rect 706 3203 709 3216
rect 714 3186 717 3316
rect 722 3243 725 3326
rect 754 3316 757 3383
rect 746 3313 757 3316
rect 746 3246 749 3313
rect 766 3306 769 3383
rect 762 3303 769 3306
rect 746 3243 757 3246
rect 754 3226 757 3243
rect 762 3236 765 3303
rect 778 3246 781 3416
rect 786 3413 789 3533
rect 786 3323 789 3336
rect 778 3243 785 3246
rect 762 3233 773 3236
rect 710 3183 717 3186
rect 710 3126 713 3183
rect 710 3123 717 3126
rect 722 3123 725 3226
rect 754 3223 765 3226
rect 738 3183 741 3206
rect 746 3203 765 3206
rect 738 3133 741 3166
rect 698 3103 705 3106
rect 658 3063 669 3066
rect 634 3013 645 3016
rect 642 2996 645 3013
rect 610 2933 613 2946
rect 634 2876 637 2996
rect 642 2993 649 2996
rect 658 2993 661 3063
rect 702 3036 705 3103
rect 714 3046 717 3123
rect 730 3103 733 3116
rect 714 3043 721 3046
rect 702 3033 709 3036
rect 626 2873 637 2876
rect 626 2826 629 2873
rect 646 2856 649 2993
rect 674 2943 677 3006
rect 698 2966 701 3016
rect 690 2963 701 2966
rect 658 2886 661 2926
rect 690 2916 693 2963
rect 706 2923 709 3033
rect 718 2946 721 3043
rect 754 3026 757 3136
rect 762 3123 765 3176
rect 754 3023 765 3026
rect 746 3013 757 3016
rect 762 3013 765 3023
rect 770 3013 773 3233
rect 782 3176 785 3243
rect 778 3173 785 3176
rect 794 3173 797 3606
rect 806 3566 809 3613
rect 802 3563 809 3566
rect 802 3516 805 3563
rect 810 3533 813 3546
rect 818 3533 821 3596
rect 826 3516 829 4163
rect 834 4023 837 4146
rect 834 3913 837 3926
rect 834 3803 837 3816
rect 834 3723 837 3736
rect 834 3593 837 3606
rect 802 3513 813 3516
rect 810 3446 813 3513
rect 802 3443 813 3446
rect 822 3513 829 3516
rect 822 3446 825 3513
rect 822 3443 829 3446
rect 802 3423 805 3443
rect 826 3423 829 3443
rect 778 3076 781 3173
rect 802 3136 805 3416
rect 810 3303 813 3326
rect 798 3133 805 3136
rect 778 3073 789 3076
rect 786 3006 789 3073
rect 778 3003 789 3006
rect 778 2946 781 3003
rect 798 2986 801 3133
rect 798 2983 805 2986
rect 802 2963 805 2983
rect 714 2943 721 2946
rect 762 2943 781 2946
rect 714 2923 717 2943
rect 690 2913 701 2916
rect 658 2883 669 2886
rect 642 2853 649 2856
rect 626 2823 637 2826
rect 466 2723 477 2726
rect 530 2723 533 2806
rect 458 2653 461 2706
rect 466 2636 469 2723
rect 562 2713 565 2726
rect 570 2706 573 2806
rect 634 2803 637 2823
rect 586 2726 589 2746
rect 538 2686 541 2706
rect 562 2703 573 2706
rect 582 2723 589 2726
rect 458 2633 469 2636
rect 530 2683 541 2686
rect 410 2533 413 2546
rect 418 2516 421 2526
rect 394 2513 421 2516
rect 426 2513 429 2536
rect 434 2533 437 2546
rect 386 2493 397 2496
rect 394 2446 397 2493
rect 370 2443 377 2446
rect 386 2443 397 2446
rect 434 2443 437 2526
rect 458 2523 461 2633
rect 530 2626 533 2683
rect 474 2583 477 2606
rect 482 2593 485 2606
rect 490 2566 493 2626
rect 530 2623 541 2626
rect 506 2596 509 2616
rect 482 2563 493 2566
rect 502 2593 509 2596
rect 362 2423 365 2436
rect 370 2416 373 2443
rect 362 2413 373 2416
rect 362 2393 365 2413
rect 354 2343 365 2346
rect 338 2313 345 2316
rect 342 2206 345 2313
rect 354 2303 357 2336
rect 362 2323 365 2343
rect 338 2203 345 2206
rect 314 2113 317 2136
rect 322 2133 325 2186
rect 338 2136 341 2203
rect 330 2133 341 2136
rect 330 2116 333 2133
rect 326 2113 333 2116
rect 326 2046 329 2113
rect 326 2043 333 2046
rect 322 1973 325 2026
rect 330 2006 333 2043
rect 338 2013 341 2126
rect 346 2103 349 2136
rect 354 2116 357 2216
rect 362 2133 365 2296
rect 370 2223 373 2346
rect 378 2303 381 2426
rect 386 2423 389 2443
rect 482 2436 485 2563
rect 502 2526 505 2593
rect 514 2533 517 2586
rect 538 2563 541 2623
rect 546 2596 549 2686
rect 562 2613 565 2703
rect 570 2596 573 2696
rect 582 2626 585 2723
rect 594 2683 597 2786
rect 602 2713 605 2736
rect 618 2726 621 2746
rect 642 2743 645 2853
rect 650 2823 653 2836
rect 658 2803 661 2836
rect 666 2733 669 2883
rect 682 2803 685 2816
rect 690 2813 693 2836
rect 698 2803 701 2913
rect 738 2813 741 2826
rect 610 2723 621 2726
rect 610 2643 613 2723
rect 706 2713 709 2726
rect 546 2593 557 2596
rect 502 2523 509 2526
rect 434 2423 437 2436
rect 482 2433 493 2436
rect 418 2413 445 2416
rect 386 2343 389 2406
rect 490 2383 493 2433
rect 498 2423 501 2436
rect 506 2416 509 2523
rect 522 2433 525 2526
rect 530 2486 533 2536
rect 538 2503 541 2526
rect 554 2496 557 2593
rect 546 2493 557 2496
rect 566 2593 573 2596
rect 578 2623 585 2626
rect 530 2483 537 2486
rect 498 2413 509 2416
rect 418 2276 421 2296
rect 434 2286 437 2306
rect 474 2303 477 2326
rect 482 2286 485 2336
rect 434 2283 445 2286
rect 410 2273 421 2276
rect 410 2216 413 2273
rect 426 2223 429 2236
rect 442 2216 445 2283
rect 474 2283 485 2286
rect 474 2236 477 2283
rect 474 2233 485 2236
rect 410 2213 421 2216
rect 370 2123 373 2206
rect 354 2113 361 2116
rect 330 2003 341 2006
rect 322 1876 325 1926
rect 330 1923 333 1946
rect 314 1873 325 1876
rect 314 1813 317 1873
rect 338 1823 341 2003
rect 346 1923 349 2096
rect 358 2046 361 2113
rect 354 2043 361 2046
rect 354 2016 357 2043
rect 378 2033 381 2156
rect 418 2143 421 2213
rect 426 2203 429 2216
rect 434 2213 445 2216
rect 482 2213 485 2233
rect 490 2213 493 2326
rect 410 2123 413 2136
rect 418 2113 421 2136
rect 434 2123 437 2213
rect 498 2203 501 2413
rect 506 2283 509 2406
rect 442 2143 445 2196
rect 514 2153 517 2336
rect 522 2306 525 2426
rect 534 2346 537 2483
rect 530 2343 537 2346
rect 530 2323 533 2343
rect 546 2323 549 2493
rect 566 2426 569 2593
rect 566 2423 573 2426
rect 578 2423 581 2623
rect 522 2303 533 2306
rect 530 2166 533 2303
rect 554 2293 557 2336
rect 522 2163 533 2166
rect 450 2116 453 2136
rect 458 2133 461 2146
rect 522 2123 525 2163
rect 446 2113 453 2116
rect 446 2046 449 2113
rect 530 2066 533 2086
rect 446 2043 453 2046
rect 354 2013 365 2016
rect 450 2013 453 2043
rect 458 2013 461 2066
rect 526 2063 533 2066
rect 362 1993 365 2013
rect 466 1976 469 2006
rect 354 1956 357 1976
rect 458 1973 469 1976
rect 354 1953 365 1956
rect 362 1866 365 1953
rect 354 1863 365 1866
rect 314 1786 317 1806
rect 330 1793 333 1816
rect 314 1783 321 1786
rect 298 1673 309 1676
rect 298 1606 301 1673
rect 318 1666 321 1783
rect 338 1766 341 1816
rect 354 1813 357 1863
rect 402 1826 405 1956
rect 458 1866 461 1973
rect 482 1956 485 2006
rect 506 1986 509 2056
rect 474 1953 485 1956
rect 502 1983 509 1986
rect 474 1886 477 1953
rect 474 1883 485 1886
rect 458 1863 469 1866
rect 394 1823 405 1826
rect 394 1776 397 1823
rect 394 1773 405 1776
rect 330 1763 341 1766
rect 330 1723 333 1763
rect 314 1663 321 1666
rect 314 1613 317 1663
rect 338 1606 341 1626
rect 298 1603 309 1606
rect 282 1576 285 1596
rect 282 1573 293 1576
rect 254 1513 261 1516
rect 242 1396 245 1406
rect 226 1393 245 1396
rect 210 1333 213 1346
rect 202 1323 213 1326
rect 122 1173 133 1176
rect 90 626 93 726
rect 114 723 117 1156
rect 130 946 133 1173
rect 178 1123 181 1246
rect 186 1123 189 1256
rect 210 1253 213 1323
rect 218 1243 221 1336
rect 226 1316 229 1376
rect 234 1323 237 1386
rect 242 1333 245 1346
rect 226 1313 237 1316
rect 202 1193 205 1206
rect 194 1166 197 1186
rect 234 1166 237 1313
rect 194 1163 205 1166
rect 186 1096 189 1116
rect 178 1093 189 1096
rect 178 1036 181 1093
rect 202 1086 205 1163
rect 194 1083 205 1086
rect 230 1163 237 1166
rect 178 1033 189 1036
rect 186 1013 189 1033
rect 194 1026 197 1083
rect 230 1036 233 1163
rect 250 1156 253 1426
rect 258 1383 261 1513
rect 274 1413 277 1546
rect 290 1406 293 1573
rect 274 1403 293 1406
rect 258 1323 261 1336
rect 266 1216 269 1316
rect 274 1306 277 1403
rect 306 1373 309 1603
rect 334 1603 341 1606
rect 334 1546 337 1603
rect 334 1543 341 1546
rect 314 1523 333 1526
rect 330 1506 333 1523
rect 322 1503 333 1506
rect 322 1436 325 1503
rect 322 1433 333 1436
rect 322 1403 325 1416
rect 298 1313 301 1326
rect 274 1303 293 1306
rect 266 1213 285 1216
rect 290 1203 293 1303
rect 242 1153 253 1156
rect 230 1033 237 1036
rect 194 1023 213 1026
rect 122 943 133 946
rect 122 923 125 943
rect 122 723 125 816
rect 162 743 165 936
rect 194 923 197 1016
rect 210 996 213 1023
rect 218 1003 221 1016
rect 234 1013 237 1033
rect 242 1013 245 1153
rect 210 993 221 996
rect 210 933 213 946
rect 218 933 221 993
rect 218 923 229 926
rect 234 923 237 946
rect 226 906 229 923
rect 218 903 229 906
rect 218 776 221 903
rect 242 886 245 1006
rect 234 883 245 886
rect 234 826 237 883
rect 250 836 253 1126
rect 274 1033 277 1196
rect 322 1146 325 1226
rect 330 1203 333 1433
rect 338 1413 341 1543
rect 338 1213 341 1236
rect 322 1143 333 1146
rect 290 1113 293 1136
rect 338 1126 341 1206
rect 346 1133 349 1746
rect 354 1613 357 1626
rect 362 1613 365 1726
rect 378 1723 381 1766
rect 402 1723 405 1773
rect 410 1766 413 1816
rect 410 1763 421 1766
rect 434 1763 437 1806
rect 418 1716 421 1763
rect 466 1756 469 1863
rect 482 1856 485 1883
rect 482 1853 493 1856
rect 410 1713 421 1716
rect 458 1753 469 1756
rect 410 1633 413 1713
rect 458 1646 461 1753
rect 490 1733 493 1853
rect 502 1776 505 1983
rect 502 1773 509 1776
rect 506 1743 509 1773
rect 458 1643 469 1646
rect 354 1593 357 1606
rect 354 1363 357 1536
rect 362 1523 365 1536
rect 370 1533 373 1616
rect 386 1556 389 1616
rect 378 1553 389 1556
rect 378 1516 381 1553
rect 386 1523 389 1546
rect 458 1533 461 1596
rect 466 1593 469 1643
rect 474 1616 477 1726
rect 490 1626 493 1726
rect 514 1723 517 2036
rect 526 1986 529 2063
rect 546 2013 549 2126
rect 526 1983 533 1986
rect 530 1963 533 1983
rect 522 1876 525 1926
rect 546 1923 549 1996
rect 554 1953 557 2206
rect 562 2153 565 2406
rect 570 2366 573 2423
rect 570 2363 581 2366
rect 570 2286 573 2346
rect 578 2306 581 2363
rect 586 2323 589 2606
rect 594 2323 597 2626
rect 610 2623 613 2636
rect 602 2496 605 2566
rect 610 2533 613 2616
rect 618 2546 621 2636
rect 626 2623 629 2706
rect 634 2613 637 2646
rect 634 2583 637 2606
rect 690 2603 693 2706
rect 698 2613 701 2636
rect 714 2623 717 2726
rect 730 2713 733 2806
rect 738 2693 741 2796
rect 746 2733 749 2926
rect 754 2703 757 2766
rect 762 2723 765 2943
rect 794 2933 797 2946
rect 778 2716 781 2816
rect 786 2806 789 2876
rect 810 2873 813 3126
rect 818 3076 821 3416
rect 834 3406 837 3516
rect 842 3486 845 4346
rect 850 4313 853 4336
rect 858 4223 861 4336
rect 850 4143 853 4206
rect 858 4173 861 4206
rect 850 4033 853 4136
rect 858 4133 861 4156
rect 866 4123 869 4353
rect 874 4106 877 4406
rect 882 4343 885 4406
rect 890 4336 893 4456
rect 898 4386 901 4536
rect 906 4503 909 4536
rect 914 4523 917 4546
rect 922 4533 933 4536
rect 938 4533 941 4556
rect 922 4513 933 4516
rect 970 4506 973 4536
rect 978 4513 981 4526
rect 986 4523 989 4536
rect 1010 4533 1021 4536
rect 970 4503 981 4506
rect 906 4403 909 4416
rect 922 4403 925 4436
rect 938 4403 941 4416
rect 954 4413 957 4476
rect 970 4423 973 4446
rect 898 4383 905 4386
rect 870 4103 877 4106
rect 882 4333 893 4336
rect 858 3806 861 4026
rect 870 3936 873 4103
rect 882 3966 885 4333
rect 890 4303 893 4326
rect 902 4296 905 4383
rect 898 4293 905 4296
rect 890 4213 893 4226
rect 890 4103 893 4126
rect 898 4086 901 4293
rect 914 4276 917 4336
rect 910 4273 917 4276
rect 910 4166 913 4273
rect 922 4216 925 4316
rect 954 4313 957 4336
rect 922 4213 933 4216
rect 962 4213 965 4366
rect 970 4353 973 4406
rect 978 4403 981 4503
rect 986 4413 989 4436
rect 994 4403 997 4426
rect 1002 4363 1005 4526
rect 1010 4516 1013 4533
rect 1010 4513 1021 4516
rect 1018 4436 1021 4513
rect 1010 4433 1021 4436
rect 1010 4403 1013 4433
rect 970 4333 973 4346
rect 978 4276 981 4326
rect 978 4273 989 4276
rect 986 4226 989 4273
rect 910 4163 917 4166
rect 894 4083 901 4086
rect 894 4006 897 4083
rect 894 4003 901 4006
rect 898 3983 901 4003
rect 906 3966 909 4146
rect 882 3963 893 3966
rect 854 3803 861 3806
rect 866 3933 873 3936
rect 854 3736 857 3803
rect 854 3733 861 3736
rect 858 3623 861 3733
rect 866 3623 869 3933
rect 874 3906 877 3926
rect 874 3903 881 3906
rect 878 3806 881 3903
rect 874 3803 881 3806
rect 850 3576 853 3616
rect 858 3593 861 3606
rect 850 3573 857 3576
rect 854 3506 857 3573
rect 866 3523 869 3546
rect 854 3503 861 3506
rect 842 3483 849 3486
rect 830 3403 837 3406
rect 830 3336 833 3403
rect 846 3396 849 3483
rect 842 3393 849 3396
rect 842 3343 845 3393
rect 858 3366 861 3503
rect 850 3363 861 3366
rect 830 3333 837 3336
rect 826 3193 829 3206
rect 834 3196 837 3333
rect 850 3223 853 3363
rect 858 3313 861 3346
rect 874 3336 877 3803
rect 890 3786 893 3963
rect 902 3963 909 3966
rect 902 3916 905 3963
rect 914 3923 917 4163
rect 922 4143 925 4206
rect 930 4196 933 4213
rect 962 4203 973 4206
rect 978 4203 981 4226
rect 986 4223 997 4226
rect 986 4213 989 4223
rect 930 4193 941 4196
rect 938 4136 941 4193
rect 902 3913 909 3916
rect 882 3783 893 3786
rect 882 3723 885 3783
rect 890 3656 893 3766
rect 906 3763 909 3913
rect 922 3823 925 4136
rect 930 4133 941 4136
rect 962 4133 965 4203
rect 930 4113 933 4133
rect 930 4003 933 4016
rect 938 3993 941 4016
rect 946 4003 949 4076
rect 970 4036 973 4146
rect 978 4123 981 4136
rect 986 4123 989 4136
rect 994 4133 997 4206
rect 970 4033 989 4036
rect 962 4023 973 4026
rect 954 4013 965 4016
rect 922 3783 925 3806
rect 930 3766 933 3986
rect 970 3956 973 4023
rect 962 3953 973 3956
rect 938 3933 941 3946
rect 938 3906 941 3926
rect 938 3903 949 3906
rect 946 3836 949 3903
rect 926 3763 933 3766
rect 938 3833 949 3836
rect 906 3733 909 3756
rect 906 3713 909 3726
rect 882 3653 893 3656
rect 882 3616 885 3653
rect 890 3623 893 3636
rect 882 3613 893 3616
rect 882 3523 885 3576
rect 890 3506 893 3613
rect 898 3606 901 3626
rect 898 3603 905 3606
rect 902 3536 905 3603
rect 886 3503 893 3506
rect 898 3533 905 3536
rect 886 3396 889 3503
rect 898 3403 901 3533
rect 914 3516 917 3726
rect 926 3636 929 3763
rect 926 3633 933 3636
rect 922 3603 925 3616
rect 910 3513 917 3516
rect 910 3436 913 3513
rect 910 3433 917 3436
rect 886 3393 893 3396
rect 874 3333 881 3336
rect 866 3293 869 3326
rect 842 3203 845 3216
rect 834 3193 845 3196
rect 818 3073 829 3076
rect 826 2986 829 3073
rect 842 3036 845 3193
rect 858 3123 861 3246
rect 866 3213 869 3266
rect 878 3246 881 3333
rect 874 3243 881 3246
rect 866 3106 869 3136
rect 822 2983 829 2986
rect 838 3033 845 3036
rect 862 3103 869 3106
rect 862 3036 865 3103
rect 862 3033 869 3036
rect 838 2986 841 3033
rect 838 2983 845 2986
rect 822 2866 825 2983
rect 818 2863 825 2866
rect 786 2803 797 2806
rect 802 2803 805 2826
rect 762 2713 781 2716
rect 618 2543 629 2546
rect 626 2536 629 2543
rect 610 2513 613 2526
rect 602 2493 609 2496
rect 606 2426 609 2493
rect 602 2423 609 2426
rect 602 2333 605 2423
rect 618 2413 621 2536
rect 626 2533 637 2536
rect 634 2523 637 2533
rect 610 2323 613 2406
rect 634 2403 637 2426
rect 650 2403 653 2546
rect 706 2413 709 2606
rect 714 2603 717 2616
rect 762 2613 765 2713
rect 778 2646 781 2706
rect 770 2643 781 2646
rect 770 2613 773 2643
rect 786 2613 789 2726
rect 794 2703 797 2803
rect 802 2713 805 2736
rect 810 2713 813 2816
rect 818 2813 821 2863
rect 818 2763 821 2806
rect 818 2706 821 2756
rect 826 2743 829 2806
rect 834 2743 837 2966
rect 842 2943 845 2983
rect 850 2936 853 3026
rect 866 3013 869 3033
rect 866 2993 869 3006
rect 874 2976 877 3243
rect 870 2973 877 2976
rect 846 2933 853 2936
rect 846 2846 849 2933
rect 842 2843 849 2846
rect 842 2813 845 2843
rect 858 2753 861 2936
rect 870 2906 873 2973
rect 882 2913 885 3226
rect 890 3223 893 3393
rect 906 3313 909 3416
rect 914 3296 917 3433
rect 922 3376 925 3526
rect 930 3513 933 3633
rect 938 3413 941 3833
rect 946 3706 949 3816
rect 954 3793 957 3816
rect 954 3723 957 3746
rect 946 3703 953 3706
rect 950 3636 953 3703
rect 946 3633 953 3636
rect 946 3566 949 3633
rect 954 3593 957 3616
rect 962 3613 965 3953
rect 970 3923 973 3946
rect 978 3933 981 4016
rect 970 3626 973 3826
rect 970 3623 981 3626
rect 962 3583 965 3606
rect 970 3566 973 3616
rect 978 3583 981 3623
rect 946 3563 957 3566
rect 930 3393 933 3406
rect 922 3373 929 3376
rect 906 3293 917 3296
rect 906 3226 909 3293
rect 926 3286 929 3373
rect 922 3283 929 3286
rect 906 3223 917 3226
rect 890 3113 893 3216
rect 906 3193 909 3206
rect 914 3176 917 3223
rect 906 3173 917 3176
rect 906 3026 909 3173
rect 922 3146 925 3283
rect 938 3223 941 3406
rect 954 3246 957 3563
rect 966 3563 973 3566
rect 966 3516 969 3563
rect 978 3523 981 3536
rect 966 3513 973 3516
rect 946 3243 957 3246
rect 946 3213 949 3243
rect 922 3143 933 3146
rect 922 3036 925 3136
rect 930 3116 933 3143
rect 938 3123 941 3136
rect 946 3123 949 3196
rect 930 3113 941 3116
rect 922 3033 929 3036
rect 890 3013 893 3026
rect 906 3023 917 3026
rect 870 2903 877 2906
rect 874 2783 877 2903
rect 890 2723 893 2956
rect 898 2933 901 2946
rect 906 2906 909 3006
rect 902 2903 909 2906
rect 902 2836 905 2903
rect 902 2833 909 2836
rect 906 2813 909 2833
rect 914 2823 917 3023
rect 926 2946 929 3033
rect 922 2943 929 2946
rect 922 2923 925 2943
rect 938 2936 941 3113
rect 954 3016 957 3226
rect 970 3196 973 3513
rect 986 3506 989 4033
rect 1002 4016 1005 4356
rect 1010 4333 1013 4346
rect 1010 4143 1013 4326
rect 1018 4313 1021 4336
rect 1026 4323 1029 4416
rect 1034 4323 1037 4336
rect 1042 4286 1045 4436
rect 1050 4403 1053 4536
rect 1058 4523 1061 4556
rect 1066 4533 1069 4546
rect 1074 4513 1077 4576
rect 1058 4413 1061 4426
rect 1074 4413 1077 4436
rect 1066 4393 1069 4406
rect 1082 4403 1085 4593
rect 1090 4543 1093 4566
rect 1122 4533 1125 4606
rect 1130 4553 1133 4616
rect 1138 4583 1141 4606
rect 1146 4573 1149 4616
rect 1090 4413 1093 4526
rect 1098 4496 1101 4516
rect 1098 4493 1109 4496
rect 1090 4396 1093 4406
rect 1074 4393 1093 4396
rect 1050 4333 1053 4346
rect 1074 4333 1077 4393
rect 1106 4386 1109 4493
rect 1138 4473 1141 4536
rect 1154 4533 1157 4606
rect 1170 4556 1173 4626
rect 1186 4603 1189 4626
rect 1210 4596 1213 4616
rect 1250 4613 1269 4616
rect 1166 4553 1173 4556
rect 1202 4593 1213 4596
rect 1146 4413 1149 4526
rect 1166 4486 1169 4553
rect 1178 4496 1181 4546
rect 1202 4533 1205 4593
rect 1194 4513 1197 4526
rect 1178 4493 1189 4496
rect 1166 4483 1173 4486
rect 1130 4403 1141 4406
rect 1098 4383 1109 4386
rect 1042 4283 1053 4286
rect 1002 4013 1013 4016
rect 1018 4013 1021 4246
rect 1026 4203 1029 4216
rect 1026 4023 1029 4136
rect 1034 4036 1037 4226
rect 1042 4183 1045 4206
rect 1042 4103 1045 4136
rect 1050 4133 1053 4283
rect 1058 4183 1061 4206
rect 1066 4203 1069 4216
rect 1074 4213 1077 4326
rect 1090 4303 1093 4336
rect 1098 4226 1101 4383
rect 1114 4306 1117 4326
rect 1122 4316 1125 4336
rect 1154 4333 1157 4406
rect 1162 4393 1165 4416
rect 1170 4346 1173 4483
rect 1186 4386 1189 4493
rect 1210 4463 1213 4526
rect 1218 4426 1221 4596
rect 1250 4533 1253 4613
rect 1226 4513 1229 4526
rect 1178 4383 1189 4386
rect 1210 4423 1221 4426
rect 1178 4363 1181 4383
rect 1170 4343 1181 4346
rect 1122 4313 1133 4316
rect 1110 4303 1117 4306
rect 1110 4236 1113 4303
rect 1130 4266 1133 4313
rect 1178 4286 1181 4343
rect 1210 4333 1213 4423
rect 1218 4393 1221 4406
rect 1226 4316 1229 4416
rect 1242 4403 1245 4426
rect 1122 4263 1133 4266
rect 1162 4283 1181 4286
rect 1218 4313 1229 4316
rect 1110 4233 1117 4236
rect 1090 4223 1101 4226
rect 1090 4213 1093 4223
rect 1114 4213 1117 4233
rect 1122 4213 1125 4263
rect 1082 4193 1085 4206
rect 1098 4183 1101 4206
rect 1050 4036 1053 4126
rect 1098 4043 1101 4136
rect 1034 4033 1053 4036
rect 1010 4006 1013 4013
rect 1002 3946 1005 4006
rect 1010 4003 1021 4006
rect 1018 3986 1021 4003
rect 1026 3993 1029 4006
rect 1018 3983 1029 3986
rect 1002 3943 1021 3946
rect 994 3913 997 3936
rect 1002 3903 1005 3926
rect 1018 3823 1021 3943
rect 1026 3916 1029 3983
rect 1034 3933 1037 4033
rect 1026 3913 1033 3916
rect 1042 3913 1045 4006
rect 1050 4003 1053 4026
rect 1050 3923 1053 3936
rect 1058 3916 1061 4036
rect 1066 4003 1069 4016
rect 1098 4003 1101 4016
rect 1066 3933 1069 3946
rect 1074 3923 1077 3936
rect 1082 3933 1085 3946
rect 1090 3923 1093 3936
rect 1058 3913 1077 3916
rect 1030 3816 1033 3913
rect 994 3796 997 3816
rect 1026 3813 1033 3816
rect 994 3793 1005 3796
rect 1002 3636 1005 3793
rect 1026 3713 1029 3813
rect 1042 3803 1045 3816
rect 1050 3786 1053 3906
rect 1058 3793 1061 3806
rect 1050 3783 1061 3786
rect 1050 3733 1053 3756
rect 994 3633 1005 3636
rect 994 3583 997 3633
rect 1042 3626 1045 3726
rect 1002 3603 1005 3616
rect 1018 3593 1021 3606
rect 994 3533 997 3546
rect 1002 3523 1005 3536
rect 1010 3533 1013 3546
rect 1018 3523 1021 3536
rect 986 3503 997 3506
rect 994 3376 997 3503
rect 1026 3403 1029 3626
rect 1042 3623 1053 3626
rect 1058 3623 1061 3783
rect 1066 3766 1069 3826
rect 1074 3813 1077 3913
rect 1106 3903 1109 4136
rect 1130 4133 1133 4146
rect 1114 4096 1117 4126
rect 1138 4103 1141 4126
rect 1146 4123 1149 4136
rect 1162 4133 1165 4283
rect 1218 4246 1221 4313
rect 1242 4306 1245 4326
rect 1238 4303 1245 4306
rect 1218 4243 1229 4246
rect 1178 4193 1181 4216
rect 1186 4123 1189 4146
rect 1202 4136 1205 4206
rect 1226 4203 1229 4243
rect 1238 4236 1241 4303
rect 1250 4293 1253 4416
rect 1258 4376 1261 4536
rect 1266 4523 1269 4606
rect 1274 4533 1277 4546
rect 1282 4523 1285 4536
rect 1266 4393 1269 4416
rect 1290 4413 1293 4556
rect 1298 4523 1301 4536
rect 1306 4523 1309 4636
rect 1314 4613 1325 4616
rect 1314 4533 1317 4606
rect 1322 4503 1325 4613
rect 1386 4603 1389 4616
rect 1330 4533 1333 4556
rect 1346 4513 1349 4556
rect 1434 4553 1437 4606
rect 1482 4593 1485 4606
rect 1370 4523 1373 4546
rect 1322 4413 1325 4426
rect 1258 4373 1269 4376
rect 1238 4233 1245 4236
rect 1242 4213 1245 4233
rect 1250 4216 1253 4286
rect 1250 4213 1261 4216
rect 1250 4193 1253 4206
rect 1202 4133 1213 4136
rect 1114 4093 1125 4096
rect 1122 4026 1125 4093
rect 1186 4026 1189 4106
rect 1210 4086 1213 4133
rect 1258 4116 1261 4213
rect 1266 4203 1269 4373
rect 1282 4323 1285 4336
rect 1298 4333 1301 4346
rect 1290 4293 1293 4326
rect 1306 4323 1309 4336
rect 1314 4216 1317 4366
rect 1322 4306 1325 4336
rect 1322 4303 1333 4306
rect 1330 4236 1333 4303
rect 1354 4283 1357 4326
rect 1274 4203 1277 4216
rect 1290 4193 1293 4206
rect 1298 4203 1301 4216
rect 1306 4213 1317 4216
rect 1322 4233 1333 4236
rect 1274 4133 1293 4136
rect 1274 4123 1277 4133
rect 1250 4113 1261 4116
rect 1282 4113 1285 4126
rect 1298 4123 1301 4156
rect 1210 4083 1221 4086
rect 1114 4023 1125 4026
rect 1178 4023 1189 4026
rect 1114 4003 1117 4023
rect 1122 3923 1125 4006
rect 1138 3963 1141 4016
rect 1178 3956 1181 4023
rect 1130 3906 1133 3936
rect 1122 3903 1133 3906
rect 1122 3836 1125 3903
rect 1122 3833 1133 3836
rect 1138 3833 1141 3936
rect 1154 3933 1157 3946
rect 1146 3903 1149 3926
rect 1162 3923 1165 3956
rect 1178 3953 1189 3956
rect 1066 3763 1077 3766
rect 1066 3733 1069 3746
rect 1074 3723 1077 3763
rect 1034 3593 1037 3606
rect 1042 3603 1045 3616
rect 1050 3563 1053 3623
rect 1058 3506 1061 3616
rect 1082 3613 1085 3816
rect 1106 3803 1109 3826
rect 1114 3803 1125 3806
rect 1130 3776 1133 3833
rect 1170 3826 1173 3936
rect 1138 3803 1141 3816
rect 1146 3813 1149 3826
rect 1162 3823 1173 3826
rect 1162 3803 1165 3823
rect 1130 3773 1149 3776
rect 1050 3503 1061 3506
rect 986 3373 997 3376
rect 1050 3376 1053 3503
rect 1066 3413 1069 3536
rect 1074 3523 1077 3606
rect 1090 3573 1093 3606
rect 1098 3603 1101 3616
rect 1122 3613 1125 3736
rect 1130 3733 1141 3736
rect 1146 3706 1149 3773
rect 1154 3733 1157 3756
rect 1142 3703 1149 3706
rect 1106 3593 1109 3606
rect 1106 3566 1109 3586
rect 1082 3533 1085 3546
rect 1082 3413 1085 3526
rect 1050 3373 1061 3376
rect 986 3313 989 3373
rect 994 3333 997 3356
rect 1058 3353 1061 3373
rect 994 3203 997 3326
rect 1034 3323 1037 3346
rect 1042 3323 1045 3336
rect 1050 3333 1061 3336
rect 970 3193 989 3196
rect 962 3113 965 3126
rect 970 3023 973 3136
rect 978 3123 981 3186
rect 986 3116 989 3193
rect 978 3113 989 3116
rect 978 3046 981 3113
rect 1002 3063 1005 3126
rect 1010 3106 1013 3216
rect 1026 3123 1029 3316
rect 1050 3313 1053 3326
rect 1066 3266 1069 3406
rect 1098 3386 1101 3566
rect 1106 3563 1117 3566
rect 1094 3383 1101 3386
rect 1082 3323 1085 3356
rect 1094 3306 1097 3383
rect 1114 3376 1117 3563
rect 1090 3303 1097 3306
rect 1106 3373 1117 3376
rect 1066 3263 1077 3266
rect 1042 3223 1061 3226
rect 1042 3213 1045 3223
rect 1034 3113 1037 3136
rect 1042 3133 1045 3206
rect 1050 3143 1053 3216
rect 1058 3203 1061 3223
rect 1066 3213 1069 3226
rect 1066 3133 1069 3206
rect 1058 3116 1061 3126
rect 1074 3123 1077 3263
rect 1090 3236 1093 3303
rect 1090 3233 1101 3236
rect 1082 3193 1085 3216
rect 1058 3113 1069 3116
rect 1010 3103 1021 3106
rect 1018 3056 1021 3103
rect 1010 3053 1021 3056
rect 978 3043 989 3046
rect 950 3013 957 3016
rect 950 2956 953 3013
rect 950 2953 957 2956
rect 938 2933 945 2936
rect 954 2933 957 2953
rect 914 2803 917 2816
rect 914 2723 917 2796
rect 922 2706 925 2916
rect 930 2813 933 2926
rect 942 2836 945 2933
rect 938 2833 945 2836
rect 938 2743 941 2833
rect 818 2703 829 2706
rect 730 2533 733 2546
rect 762 2533 765 2596
rect 738 2523 757 2526
rect 618 2333 621 2386
rect 578 2303 597 2306
rect 570 2283 581 2286
rect 578 2196 581 2283
rect 570 2193 581 2196
rect 570 2143 573 2193
rect 594 2176 597 2303
rect 578 2173 597 2176
rect 562 2083 565 2136
rect 562 2013 565 2076
rect 578 2033 581 2173
rect 586 2123 589 2156
rect 626 2153 629 2396
rect 666 2393 669 2406
rect 634 2343 645 2346
rect 634 2303 637 2336
rect 690 2256 693 2276
rect 682 2253 693 2256
rect 682 2176 685 2253
rect 682 2173 689 2176
rect 594 2033 597 2136
rect 626 2133 629 2146
rect 674 2136 677 2156
rect 666 2133 677 2136
rect 618 2113 629 2116
rect 666 2046 669 2133
rect 686 2106 689 2173
rect 698 2113 701 2296
rect 714 2123 717 2236
rect 730 2213 733 2326
rect 738 2323 741 2396
rect 746 2333 749 2356
rect 686 2103 693 2106
rect 666 2043 677 2046
rect 570 2003 573 2016
rect 666 2013 669 2026
rect 578 1993 581 2006
rect 626 1986 629 2006
rect 610 1966 613 1986
rect 626 1983 637 1986
rect 522 1873 533 1876
rect 530 1826 533 1873
rect 522 1823 533 1826
rect 522 1786 525 1823
rect 522 1783 533 1786
rect 530 1716 533 1783
rect 562 1723 565 1966
rect 606 1963 613 1966
rect 594 1906 597 1926
rect 586 1903 597 1906
rect 586 1766 589 1903
rect 606 1886 609 1963
rect 634 1936 637 1983
rect 626 1933 637 1936
rect 606 1883 613 1886
rect 586 1763 605 1766
rect 522 1713 533 1716
rect 522 1633 525 1713
rect 578 1633 581 1726
rect 594 1693 597 1736
rect 490 1623 497 1626
rect 474 1613 485 1616
rect 474 1523 477 1596
rect 482 1523 485 1613
rect 494 1556 497 1623
rect 490 1553 497 1556
rect 370 1513 381 1516
rect 370 1456 373 1513
rect 362 1453 373 1456
rect 354 1203 357 1216
rect 362 1186 365 1453
rect 370 1396 373 1416
rect 378 1403 381 1436
rect 386 1396 389 1406
rect 370 1393 389 1396
rect 386 1333 389 1346
rect 394 1326 397 1336
rect 378 1323 397 1326
rect 394 1313 397 1323
rect 402 1303 405 1416
rect 410 1306 413 1356
rect 434 1353 437 1416
rect 458 1413 461 1506
rect 490 1496 493 1553
rect 482 1493 493 1496
rect 482 1426 485 1493
rect 474 1423 485 1426
rect 450 1363 453 1406
rect 410 1303 421 1306
rect 434 1303 437 1326
rect 442 1313 445 1326
rect 370 1223 373 1236
rect 378 1213 381 1226
rect 370 1193 373 1206
rect 410 1193 413 1216
rect 362 1183 373 1186
rect 354 1133 357 1146
rect 338 1123 349 1126
rect 346 1103 349 1123
rect 354 1113 357 1126
rect 370 1056 373 1183
rect 370 1053 377 1056
rect 266 993 269 1016
rect 258 903 261 926
rect 266 923 269 936
rect 274 916 277 1026
rect 266 913 277 916
rect 250 833 257 836
rect 234 823 245 826
rect 242 803 245 823
rect 254 786 257 833
rect 250 783 257 786
rect 218 773 225 776
rect 74 623 93 626
rect 74 603 77 623
rect 82 413 85 616
rect 90 613 93 623
rect 138 543 141 616
rect 146 586 149 616
rect 170 613 173 726
rect 146 583 153 586
rect 106 446 109 526
rect 130 506 133 536
rect 150 516 153 583
rect 170 573 173 606
rect 194 603 197 746
rect 222 716 225 773
rect 250 766 253 783
rect 242 763 253 766
rect 234 723 237 736
rect 222 713 229 716
rect 226 613 229 713
rect 242 656 245 763
rect 266 733 269 913
rect 282 893 285 1016
rect 290 933 293 1006
rect 306 1003 309 1036
rect 330 1013 333 1026
rect 374 996 377 1053
rect 386 1013 389 1146
rect 394 1103 397 1126
rect 402 1116 405 1156
rect 418 1133 421 1303
rect 434 1196 437 1296
rect 458 1293 461 1346
rect 474 1343 477 1423
rect 434 1193 445 1196
rect 458 1193 461 1206
rect 474 1203 477 1216
rect 482 1203 485 1416
rect 490 1393 493 1406
rect 498 1396 501 1526
rect 506 1516 509 1596
rect 506 1513 513 1516
rect 510 1436 513 1513
rect 510 1433 517 1436
rect 522 1433 525 1546
rect 538 1506 541 1526
rect 534 1503 541 1506
rect 514 1413 517 1433
rect 534 1426 537 1503
rect 534 1423 541 1426
rect 522 1403 525 1416
rect 498 1393 517 1396
rect 530 1393 533 1406
rect 538 1403 541 1423
rect 546 1413 549 1536
rect 562 1416 565 1616
rect 578 1523 581 1616
rect 594 1613 597 1626
rect 602 1613 605 1763
rect 610 1613 613 1883
rect 586 1516 589 1566
rect 558 1413 565 1416
rect 578 1513 589 1516
rect 578 1416 581 1513
rect 594 1506 597 1606
rect 610 1563 613 1606
rect 618 1553 621 1826
rect 626 1733 629 1933
rect 650 1923 653 1956
rect 674 1953 677 2043
rect 690 2016 693 2103
rect 722 2066 725 2136
rect 738 2123 741 2306
rect 746 2216 749 2326
rect 754 2293 757 2446
rect 762 2303 765 2516
rect 770 2323 773 2406
rect 778 2396 781 2536
rect 786 2523 789 2606
rect 794 2593 797 2606
rect 802 2413 805 2616
rect 818 2526 821 2616
rect 826 2613 829 2703
rect 834 2606 837 2646
rect 882 2623 885 2706
rect 918 2703 925 2706
rect 918 2636 921 2703
rect 930 2643 933 2736
rect 938 2713 941 2736
rect 918 2633 925 2636
rect 922 2616 925 2633
rect 842 2613 853 2616
rect 810 2523 821 2526
rect 826 2603 837 2606
rect 810 2513 813 2523
rect 826 2403 829 2603
rect 850 2586 853 2613
rect 842 2583 853 2586
rect 842 2466 845 2583
rect 858 2543 861 2616
rect 914 2613 925 2616
rect 866 2563 869 2606
rect 930 2596 933 2636
rect 946 2623 949 2816
rect 954 2763 957 2926
rect 962 2916 965 3006
rect 970 2943 973 3006
rect 986 2956 989 3043
rect 1010 2983 1013 3053
rect 1018 2993 1021 3016
rect 978 2953 989 2956
rect 978 2933 981 2953
rect 962 2913 973 2916
rect 970 2846 973 2913
rect 962 2843 973 2846
rect 962 2813 965 2843
rect 986 2826 989 2926
rect 994 2923 997 2936
rect 1026 2913 1029 2926
rect 1034 2923 1037 3066
rect 1066 3036 1069 3113
rect 1066 3033 1077 3036
rect 1074 3013 1077 3033
rect 1082 3013 1085 3156
rect 1090 3133 1093 3206
rect 1098 3116 1101 3233
rect 1094 3113 1101 3116
rect 1082 2933 1085 2946
rect 1082 2906 1085 2926
rect 1074 2903 1085 2906
rect 1074 2846 1077 2903
rect 1074 2843 1085 2846
rect 970 2823 989 2826
rect 962 2793 965 2806
rect 922 2593 933 2596
rect 842 2463 849 2466
rect 834 2423 837 2446
rect 778 2393 797 2396
rect 794 2256 797 2393
rect 846 2346 849 2463
rect 858 2413 861 2536
rect 922 2523 925 2593
rect 938 2536 941 2616
rect 954 2613 957 2746
rect 962 2696 965 2726
rect 970 2716 973 2823
rect 978 2813 997 2816
rect 1082 2813 1085 2843
rect 1094 2836 1097 3113
rect 1106 3006 1109 3373
rect 1114 3333 1117 3356
rect 1114 3306 1117 3326
rect 1122 3323 1125 3336
rect 1114 3303 1121 3306
rect 1118 3226 1121 3303
rect 1130 3283 1133 3656
rect 1142 3626 1145 3703
rect 1142 3623 1149 3626
rect 1146 3556 1149 3623
rect 1154 3573 1157 3726
rect 1162 3713 1165 3726
rect 1170 3723 1173 3823
rect 1178 3793 1181 3806
rect 1186 3773 1189 3953
rect 1194 3933 1197 4016
rect 1218 3993 1221 4083
rect 1202 3923 1205 3976
rect 1250 3973 1253 4113
rect 1306 4083 1309 4213
rect 1210 3836 1213 3936
rect 1218 3923 1221 3956
rect 1226 3933 1229 3966
rect 1234 3883 1237 3936
rect 1266 3856 1269 4006
rect 1290 3933 1293 4016
rect 1314 4003 1317 4206
rect 1322 4153 1325 4233
rect 1362 4223 1365 4336
rect 1370 4316 1373 4516
rect 1386 4413 1389 4536
rect 1394 4513 1397 4546
rect 1434 4533 1437 4546
rect 1410 4523 1429 4526
rect 1378 4333 1381 4366
rect 1394 4353 1397 4416
rect 1410 4403 1413 4523
rect 1418 4363 1421 4516
rect 1426 4413 1429 4426
rect 1434 4416 1437 4516
rect 1442 4426 1445 4526
rect 1450 4436 1453 4536
rect 1474 4533 1477 4586
rect 1506 4583 1509 4616
rect 1594 4606 1597 4616
rect 1594 4603 1613 4606
rect 1466 4493 1469 4526
rect 1482 4523 1485 4566
rect 1490 4466 1493 4536
rect 1498 4523 1501 4536
rect 1514 4533 1517 4546
rect 1506 4513 1509 4526
rect 1482 4463 1493 4466
rect 1450 4433 1461 4436
rect 1442 4423 1453 4426
rect 1434 4413 1445 4416
rect 1434 4393 1437 4406
rect 1442 4376 1445 4413
rect 1434 4373 1445 4376
rect 1370 4313 1377 4316
rect 1374 4226 1377 4313
rect 1386 4306 1389 4326
rect 1434 4316 1437 4373
rect 1450 4323 1453 4423
rect 1458 4413 1461 4433
rect 1466 4403 1469 4416
rect 1482 4413 1485 4463
rect 1482 4366 1485 4406
rect 1506 4393 1509 4416
rect 1474 4363 1485 4366
rect 1434 4313 1445 4316
rect 1386 4303 1397 4306
rect 1394 4236 1397 4303
rect 1442 4256 1445 4313
rect 1370 4223 1377 4226
rect 1386 4233 1397 4236
rect 1434 4253 1445 4256
rect 1330 4143 1333 4206
rect 1338 4166 1341 4216
rect 1346 4193 1349 4206
rect 1354 4203 1357 4216
rect 1338 4163 1357 4166
rect 1370 4163 1373 4223
rect 1330 4133 1341 4136
rect 1322 4113 1325 4126
rect 1338 4116 1341 4126
rect 1346 4123 1349 4156
rect 1354 4116 1357 4163
rect 1378 4126 1381 4206
rect 1386 4183 1389 4233
rect 1362 4123 1381 4126
rect 1394 4123 1397 4146
rect 1402 4116 1405 4196
rect 1434 4176 1437 4253
rect 1466 4213 1469 4226
rect 1434 4173 1461 4176
rect 1442 4133 1445 4166
rect 1338 4113 1357 4116
rect 1394 4113 1405 4116
rect 1338 4093 1341 4113
rect 1354 4006 1357 4016
rect 1354 4003 1373 4006
rect 1282 3923 1293 3926
rect 1298 3893 1301 3926
rect 1306 3903 1309 3936
rect 1202 3833 1213 3836
rect 1258 3853 1269 3856
rect 1202 3756 1205 3833
rect 1194 3753 1205 3756
rect 1170 3603 1173 3706
rect 1194 3666 1197 3753
rect 1194 3663 1205 3666
rect 1178 3613 1181 3646
rect 1186 3613 1197 3616
rect 1146 3553 1157 3556
rect 1154 3446 1157 3553
rect 1146 3443 1157 3446
rect 1138 3333 1141 3346
rect 1114 3223 1121 3226
rect 1114 3143 1117 3223
rect 1114 3026 1117 3116
rect 1122 3043 1125 3206
rect 1130 3153 1133 3226
rect 1146 3223 1149 3443
rect 1170 3403 1173 3426
rect 1154 3333 1157 3356
rect 1162 3333 1165 3376
rect 1178 3343 1181 3576
rect 1202 3506 1205 3663
rect 1218 3596 1221 3806
rect 1242 3793 1245 3816
rect 1258 3806 1261 3853
rect 1258 3803 1269 3806
rect 1266 3783 1269 3803
rect 1298 3733 1301 3786
rect 1250 3703 1253 3726
rect 1314 3723 1317 3816
rect 1322 3806 1325 3816
rect 1330 3813 1333 3826
rect 1346 3813 1349 3936
rect 1354 3923 1357 3976
rect 1362 3933 1365 3946
rect 1370 3913 1373 3926
rect 1378 3906 1381 3936
rect 1386 3923 1389 4016
rect 1394 4003 1397 4113
rect 1458 4106 1461 4173
rect 1450 4103 1461 4106
rect 1394 3923 1397 3936
rect 1402 3906 1405 4016
rect 1418 4013 1421 4026
rect 1410 3993 1413 4006
rect 1418 3996 1421 4006
rect 1426 3996 1429 4006
rect 1418 3993 1429 3996
rect 1418 3946 1421 3993
rect 1370 3903 1381 3906
rect 1394 3903 1405 3906
rect 1410 3943 1421 3946
rect 1322 3803 1341 3806
rect 1274 3636 1277 3706
rect 1274 3633 1285 3636
rect 1226 3603 1229 3616
rect 1218 3593 1229 3596
rect 1226 3523 1229 3593
rect 1234 3573 1237 3606
rect 1242 3583 1245 3616
rect 1250 3523 1253 3606
rect 1258 3553 1261 3626
rect 1266 3603 1269 3616
rect 1282 3576 1285 3633
rect 1322 3613 1325 3626
rect 1274 3573 1285 3576
rect 1314 3573 1317 3606
rect 1330 3593 1333 3606
rect 1338 3603 1341 3616
rect 1346 3603 1349 3806
rect 1362 3733 1365 3806
rect 1370 3803 1373 3903
rect 1370 3723 1373 3776
rect 1378 3706 1381 3816
rect 1394 3796 1397 3903
rect 1410 3886 1413 3943
rect 1406 3883 1413 3886
rect 1406 3816 1409 3883
rect 1418 3823 1421 3936
rect 1426 3893 1429 3986
rect 1450 3983 1453 4103
rect 1474 4056 1477 4363
rect 1498 4323 1501 4346
rect 1522 4313 1525 4526
rect 1530 4503 1533 4536
rect 1562 4533 1565 4596
rect 1618 4563 1621 4616
rect 1650 4546 1653 4606
rect 1586 4523 1589 4546
rect 1634 4543 1653 4546
rect 1578 4406 1581 4416
rect 1586 4413 1589 4426
rect 1578 4403 1597 4406
rect 1610 4393 1613 4406
rect 1634 4393 1637 4543
rect 1642 4533 1661 4536
rect 1642 4523 1645 4533
rect 1650 4513 1653 4526
rect 1666 4513 1669 4536
rect 1674 4523 1677 4616
rect 1746 4603 1749 4616
rect 1778 4613 1781 4626
rect 1754 4576 1757 4606
rect 1754 4573 1765 4576
rect 1714 4456 1717 4526
rect 1746 4503 1749 4526
rect 1710 4453 1717 4456
rect 1658 4413 1661 4426
rect 1690 4413 1693 4436
rect 1698 4413 1701 4426
rect 1610 4333 1629 4336
rect 1610 4323 1613 4333
rect 1634 4323 1637 4336
rect 1650 4296 1653 4396
rect 1710 4386 1713 4453
rect 1722 4413 1725 4446
rect 1722 4396 1725 4406
rect 1730 4403 1733 4436
rect 1738 4396 1741 4416
rect 1722 4393 1741 4396
rect 1710 4383 1717 4386
rect 1714 4366 1717 4383
rect 1714 4363 1721 4366
rect 1642 4293 1653 4296
rect 1514 4143 1517 4206
rect 1602 4193 1605 4206
rect 1642 4193 1645 4293
rect 1674 4226 1677 4346
rect 1698 4313 1701 4326
rect 1718 4286 1721 4363
rect 1714 4283 1721 4286
rect 1650 4213 1653 4226
rect 1670 4223 1677 4226
rect 1670 4176 1673 4223
rect 1682 4183 1685 4216
rect 1690 4213 1693 4226
rect 1706 4203 1709 4226
rect 1714 4213 1717 4283
rect 1670 4173 1677 4176
rect 1498 4123 1501 4136
rect 1554 4133 1573 4136
rect 1586 4133 1589 4156
rect 1554 4123 1557 4133
rect 1562 4113 1565 4126
rect 1466 4053 1477 4056
rect 1466 3966 1469 4053
rect 1490 3993 1493 4016
rect 1546 4006 1549 4016
rect 1554 4013 1557 4026
rect 1546 4003 1565 4006
rect 1450 3963 1469 3966
rect 1434 3903 1437 3936
rect 1406 3813 1413 3816
rect 1418 3813 1429 3816
rect 1410 3796 1413 3813
rect 1394 3793 1405 3796
rect 1410 3793 1429 3796
rect 1450 3793 1453 3963
rect 1474 3923 1477 3946
rect 1554 3933 1573 3936
rect 1554 3923 1557 3933
rect 1562 3913 1565 3926
rect 1578 3923 1581 3936
rect 1586 3856 1589 4126
rect 1610 4003 1613 4016
rect 1618 4013 1621 4026
rect 1626 4016 1629 4126
rect 1626 4013 1637 4016
rect 1650 4006 1653 4026
rect 1618 3943 1621 4006
rect 1618 3916 1621 3936
rect 1610 3913 1621 3916
rect 1610 3866 1613 3913
rect 1610 3863 1621 3866
rect 1582 3853 1589 3856
rect 1466 3803 1469 3816
rect 1562 3813 1565 3826
rect 1402 3773 1405 3793
rect 1370 3703 1381 3706
rect 1370 3636 1373 3703
rect 1370 3633 1381 3636
rect 1274 3513 1277 3573
rect 1330 3533 1349 3536
rect 1202 3503 1213 3506
rect 1202 3413 1205 3436
rect 1210 3406 1213 3503
rect 1218 3413 1221 3426
rect 1194 3393 1197 3406
rect 1210 3403 1221 3406
rect 1210 3323 1213 3336
rect 1218 3333 1221 3403
rect 1258 3393 1261 3416
rect 1306 3393 1309 3526
rect 1330 3523 1333 3533
rect 1354 3523 1357 3586
rect 1226 3336 1229 3346
rect 1226 3333 1237 3336
rect 1218 3306 1221 3326
rect 1210 3303 1221 3306
rect 1154 3213 1157 3256
rect 1210 3246 1213 3303
rect 1210 3243 1221 3246
rect 1146 3166 1149 3206
rect 1170 3193 1173 3216
rect 1218 3213 1221 3243
rect 1194 3193 1197 3206
rect 1146 3163 1165 3166
rect 1138 3113 1141 3136
rect 1162 3123 1165 3163
rect 1210 3113 1213 3156
rect 1218 3123 1221 3206
rect 1226 3193 1229 3326
rect 1234 3173 1237 3333
rect 1242 3316 1245 3336
rect 1266 3323 1269 3356
rect 1242 3313 1253 3316
rect 1250 3256 1253 3313
rect 1242 3253 1253 3256
rect 1242 3163 1245 3253
rect 1258 3213 1261 3236
rect 1226 3123 1229 3146
rect 1250 3143 1253 3206
rect 1266 3193 1269 3206
rect 1114 3023 1125 3026
rect 1114 3013 1117 3023
rect 1106 3003 1117 3006
rect 1106 2903 1109 2986
rect 1114 2876 1117 3003
rect 1122 2943 1125 3006
rect 1162 3003 1165 3026
rect 1170 2993 1173 3006
rect 1202 3003 1205 3016
rect 1210 3013 1213 3026
rect 1234 3013 1237 3136
rect 1250 3113 1253 3136
rect 1274 3106 1277 3366
rect 1290 3333 1293 3346
rect 1298 3233 1301 3326
rect 1282 3213 1285 3226
rect 1314 3166 1317 3376
rect 1322 3353 1325 3416
rect 1330 3316 1333 3466
rect 1362 3463 1365 3576
rect 1370 3556 1373 3616
rect 1378 3573 1381 3633
rect 1386 3613 1389 3756
rect 1402 3696 1405 3716
rect 1398 3693 1405 3696
rect 1398 3626 1401 3693
rect 1426 3676 1429 3793
rect 1466 3713 1469 3726
rect 1410 3673 1429 3676
rect 1410 3653 1413 3673
rect 1398 3623 1405 3626
rect 1386 3583 1389 3606
rect 1402 3603 1405 3623
rect 1410 3613 1413 3646
rect 1370 3553 1377 3556
rect 1374 3476 1377 3553
rect 1394 3533 1397 3546
rect 1370 3473 1377 3476
rect 1370 3456 1373 3473
rect 1354 3453 1373 3456
rect 1338 3323 1341 3406
rect 1346 3393 1349 3406
rect 1330 3313 1341 3316
rect 1314 3163 1321 3166
rect 1282 3123 1285 3146
rect 1274 3103 1281 3106
rect 1242 2996 1245 3056
rect 1266 3033 1269 3096
rect 1258 3023 1269 3026
rect 1234 2993 1245 2996
rect 1122 2913 1125 2936
rect 1106 2873 1117 2876
rect 1094 2833 1101 2836
rect 994 2793 997 2813
rect 978 2723 989 2726
rect 970 2713 981 2716
rect 994 2706 997 2786
rect 1026 2706 1029 2726
rect 978 2703 997 2706
rect 1018 2703 1029 2706
rect 962 2693 969 2696
rect 954 2593 957 2606
rect 966 2586 969 2693
rect 962 2583 969 2586
rect 938 2533 949 2536
rect 858 2356 861 2406
rect 874 2393 877 2406
rect 858 2353 865 2356
rect 846 2343 853 2346
rect 842 2306 845 2326
rect 778 2253 797 2256
rect 834 2303 845 2306
rect 778 2233 781 2253
rect 834 2246 837 2303
rect 834 2243 845 2246
rect 746 2213 757 2216
rect 842 2213 845 2243
rect 754 2193 757 2213
rect 762 2113 773 2116
rect 770 2083 773 2113
rect 714 2063 725 2066
rect 686 2013 693 2016
rect 686 1966 689 2013
rect 698 1976 701 2006
rect 706 2003 709 2026
rect 714 2016 717 2063
rect 778 2033 781 2136
rect 794 2043 797 2126
rect 802 2033 805 2136
rect 714 2013 725 2016
rect 810 2013 813 2116
rect 818 2013 821 2196
rect 850 2193 853 2343
rect 862 2226 865 2353
rect 882 2346 885 2516
rect 938 2513 941 2526
rect 938 2423 941 2446
rect 946 2413 949 2533
rect 954 2513 957 2536
rect 962 2523 965 2583
rect 978 2523 981 2703
rect 1018 2646 1021 2703
rect 1042 2656 1045 2796
rect 1090 2776 1093 2816
rect 1098 2813 1101 2833
rect 1098 2793 1101 2806
rect 1082 2773 1093 2776
rect 1042 2653 1049 2656
rect 1018 2643 1029 2646
rect 986 2496 989 2616
rect 994 2533 997 2606
rect 1002 2543 1005 2616
rect 1018 2613 1021 2626
rect 1026 2613 1029 2643
rect 1034 2606 1037 2646
rect 1010 2536 1013 2606
rect 1026 2603 1037 2606
rect 1010 2533 1021 2536
rect 970 2493 989 2496
rect 882 2343 889 2346
rect 898 2343 901 2406
rect 946 2343 949 2406
rect 970 2366 973 2493
rect 994 2476 997 2526
rect 1010 2513 1013 2526
rect 1026 2516 1029 2603
rect 1046 2596 1049 2653
rect 1042 2593 1049 2596
rect 1022 2513 1029 2516
rect 986 2473 997 2476
rect 986 2386 989 2473
rect 986 2383 997 2386
rect 970 2363 989 2366
rect 986 2343 989 2363
rect 858 2223 865 2226
rect 826 2023 829 2126
rect 834 2123 837 2186
rect 858 2133 861 2223
rect 722 1993 725 2013
rect 834 2006 837 2016
rect 842 2013 845 2126
rect 866 2123 869 2206
rect 874 2183 877 2336
rect 886 2246 889 2343
rect 986 2316 989 2326
rect 994 2323 997 2383
rect 1002 2333 1005 2506
rect 1022 2426 1025 2513
rect 1010 2406 1013 2426
rect 1022 2423 1029 2426
rect 1010 2403 1017 2406
rect 1014 2326 1017 2403
rect 1002 2316 1005 2326
rect 986 2313 1005 2316
rect 1010 2323 1017 2326
rect 1010 2296 1013 2323
rect 882 2243 889 2246
rect 1002 2293 1013 2296
rect 882 2213 885 2243
rect 1002 2236 1005 2293
rect 906 2213 909 2226
rect 946 2153 949 2236
rect 1002 2233 1013 2236
rect 930 2143 949 2146
rect 938 2113 941 2136
rect 946 2133 949 2143
rect 954 2123 957 2216
rect 962 2203 965 2226
rect 698 1973 709 1976
rect 686 1963 693 1966
rect 674 1923 677 1936
rect 690 1933 693 1963
rect 626 1706 629 1726
rect 634 1723 637 1916
rect 690 1913 693 1926
rect 706 1906 709 1973
rect 698 1903 709 1906
rect 698 1856 701 1903
rect 690 1853 701 1856
rect 642 1723 645 1816
rect 650 1813 653 1826
rect 690 1776 693 1853
rect 746 1813 749 1956
rect 762 1886 765 1926
rect 770 1923 773 2006
rect 794 1923 797 1936
rect 762 1883 773 1886
rect 690 1773 701 1776
rect 674 1723 677 1756
rect 698 1753 701 1773
rect 730 1726 733 1746
rect 770 1743 773 1883
rect 730 1723 741 1726
rect 626 1703 633 1706
rect 630 1626 633 1703
rect 626 1623 633 1626
rect 626 1603 629 1623
rect 642 1596 645 1696
rect 650 1603 653 1626
rect 642 1593 653 1596
rect 642 1533 645 1556
rect 594 1503 605 1506
rect 578 1413 589 1416
rect 498 1333 501 1346
rect 506 1326 509 1336
rect 490 1323 509 1326
rect 506 1313 509 1323
rect 514 1303 517 1393
rect 558 1366 561 1413
rect 570 1393 573 1406
rect 586 1366 589 1413
rect 558 1363 565 1366
rect 562 1346 565 1363
rect 578 1363 589 1366
rect 562 1343 573 1346
rect 538 1303 541 1326
rect 546 1313 549 1326
rect 442 1116 445 1193
rect 458 1116 461 1136
rect 402 1113 413 1116
rect 410 1046 413 1113
rect 402 1043 413 1046
rect 434 1113 445 1116
rect 434 1046 437 1113
rect 434 1043 445 1046
rect 402 1023 405 1043
rect 442 1003 445 1043
rect 450 1013 453 1116
rect 458 1113 465 1116
rect 462 1046 465 1113
rect 474 1083 477 1136
rect 490 1066 493 1196
rect 514 1123 517 1206
rect 538 1153 541 1226
rect 546 1223 565 1226
rect 570 1196 573 1343
rect 578 1316 581 1363
rect 602 1336 605 1503
rect 610 1496 613 1526
rect 610 1493 621 1496
rect 618 1436 621 1493
rect 610 1433 621 1436
rect 610 1413 613 1433
rect 618 1403 637 1406
rect 602 1333 613 1336
rect 578 1313 589 1316
rect 586 1246 589 1313
rect 562 1193 573 1196
rect 578 1243 589 1246
rect 458 1043 465 1046
rect 474 1063 493 1066
rect 374 993 381 996
rect 378 946 381 993
rect 450 986 453 1006
rect 446 983 453 986
rect 458 986 461 1043
rect 474 1003 477 1063
rect 498 1013 501 1086
rect 554 1013 557 1026
rect 562 1003 565 1193
rect 578 1123 581 1243
rect 586 1223 605 1226
rect 594 1113 597 1216
rect 610 1203 613 1333
rect 626 1216 629 1396
rect 642 1376 645 1416
rect 650 1393 653 1593
rect 658 1523 661 1636
rect 738 1633 741 1723
rect 754 1706 757 1726
rect 754 1703 765 1706
rect 762 1636 765 1703
rect 754 1633 765 1636
rect 754 1613 757 1633
rect 786 1613 789 1766
rect 810 1763 813 1926
rect 826 1913 829 2006
rect 834 2003 845 2006
rect 842 1923 845 2003
rect 850 1966 853 2036
rect 858 1983 861 2046
rect 850 1963 857 1966
rect 854 1896 857 1963
rect 850 1893 857 1896
rect 850 1876 853 1893
rect 842 1873 853 1876
rect 842 1746 845 1873
rect 866 1766 869 2006
rect 874 1953 877 2036
rect 890 1923 893 1936
rect 906 1923 917 1926
rect 914 1836 917 1916
rect 914 1833 921 1836
rect 898 1796 901 1816
rect 894 1793 901 1796
rect 866 1763 873 1766
rect 802 1733 805 1746
rect 842 1743 853 1746
rect 850 1723 853 1743
rect 870 1706 873 1763
rect 866 1703 873 1706
rect 866 1686 869 1703
rect 858 1683 869 1686
rect 666 1576 669 1596
rect 666 1573 677 1576
rect 674 1516 677 1573
rect 666 1513 677 1516
rect 666 1413 669 1513
rect 682 1393 685 1406
rect 690 1403 693 1536
rect 706 1506 709 1526
rect 706 1503 717 1506
rect 714 1436 717 1503
rect 706 1433 717 1436
rect 706 1416 709 1433
rect 738 1426 741 1556
rect 770 1553 773 1606
rect 762 1513 765 1536
rect 770 1523 773 1536
rect 802 1523 805 1616
rect 738 1423 757 1426
rect 702 1413 709 1416
rect 642 1373 653 1376
rect 650 1226 653 1373
rect 702 1336 705 1413
rect 682 1323 685 1336
rect 698 1333 705 1336
rect 682 1296 685 1316
rect 674 1293 685 1296
rect 674 1236 677 1293
rect 674 1233 685 1236
rect 690 1233 693 1326
rect 698 1303 701 1333
rect 706 1286 709 1326
rect 714 1323 717 1396
rect 722 1333 725 1406
rect 730 1403 733 1416
rect 754 1326 757 1423
rect 778 1403 781 1426
rect 786 1393 789 1496
rect 802 1413 805 1456
rect 810 1413 813 1436
rect 730 1323 757 1326
rect 702 1283 709 1286
rect 642 1223 653 1226
rect 626 1213 633 1216
rect 578 1003 581 1016
rect 602 1013 605 1136
rect 618 1126 621 1206
rect 630 1166 633 1213
rect 626 1163 633 1166
rect 626 1146 629 1163
rect 626 1143 637 1146
rect 642 1133 645 1223
rect 682 1213 685 1233
rect 618 1123 629 1126
rect 658 1116 661 1206
rect 690 1156 693 1226
rect 682 1153 693 1156
rect 650 1113 661 1116
rect 650 1036 653 1113
rect 650 1033 661 1036
rect 658 1013 661 1033
rect 666 1023 669 1136
rect 682 1113 685 1153
rect 702 1146 705 1283
rect 702 1143 709 1146
rect 690 1066 693 1136
rect 706 1126 709 1143
rect 714 1133 717 1306
rect 730 1266 733 1323
rect 722 1263 733 1266
rect 722 1203 725 1263
rect 762 1213 765 1236
rect 786 1226 789 1246
rect 778 1223 789 1226
rect 738 1136 741 1206
rect 778 1176 781 1223
rect 818 1213 821 1626
rect 858 1613 861 1683
rect 882 1603 885 1746
rect 894 1646 897 1793
rect 894 1643 901 1646
rect 898 1603 901 1643
rect 834 1413 837 1536
rect 842 1513 845 1526
rect 850 1496 853 1546
rect 846 1493 853 1496
rect 846 1426 849 1493
rect 858 1453 861 1526
rect 866 1523 869 1556
rect 898 1533 901 1586
rect 898 1506 901 1526
rect 890 1503 901 1506
rect 890 1446 893 1503
rect 890 1443 901 1446
rect 846 1423 853 1426
rect 842 1333 845 1346
rect 850 1333 853 1423
rect 874 1413 877 1426
rect 842 1316 845 1326
rect 858 1323 861 1346
rect 882 1333 885 1416
rect 898 1403 901 1443
rect 906 1396 909 1826
rect 918 1746 921 1833
rect 914 1743 921 1746
rect 914 1603 917 1743
rect 922 1706 925 1726
rect 922 1703 929 1706
rect 914 1413 917 1596
rect 926 1576 929 1703
rect 922 1573 929 1576
rect 922 1476 925 1573
rect 922 1473 929 1476
rect 926 1406 929 1473
rect 898 1393 909 1396
rect 922 1403 929 1406
rect 842 1313 869 1316
rect 866 1213 869 1313
rect 890 1213 893 1226
rect 778 1173 789 1176
rect 730 1133 741 1136
rect 698 1123 709 1126
rect 690 1063 709 1066
rect 682 1003 685 1016
rect 706 1013 709 1063
rect 458 983 469 986
rect 314 936 317 946
rect 306 933 317 936
rect 370 943 381 946
rect 306 803 309 933
rect 314 896 317 926
rect 322 913 325 926
rect 330 903 333 916
rect 338 906 341 926
rect 370 923 373 943
rect 418 933 421 946
rect 338 903 349 906
rect 314 893 333 896
rect 314 813 317 826
rect 330 823 333 893
rect 346 846 349 903
rect 338 843 349 846
rect 338 773 341 843
rect 354 813 357 826
rect 298 733 301 746
rect 238 653 245 656
rect 238 586 241 653
rect 238 583 245 586
rect 114 503 133 506
rect 98 443 109 446
rect 98 403 101 443
rect 122 403 125 496
rect 138 423 141 516
rect 146 513 153 516
rect 146 493 149 513
rect 82 323 85 336
rect 130 323 133 416
rect 138 333 141 406
rect 162 403 165 546
rect 178 513 181 526
rect 186 413 189 516
rect 194 503 197 526
rect 202 516 205 566
rect 242 563 245 583
rect 226 533 237 536
rect 234 516 237 526
rect 242 523 245 546
rect 250 516 253 536
rect 202 513 213 516
rect 210 436 213 513
rect 202 433 213 436
rect 234 513 253 516
rect 258 513 261 526
rect 274 523 277 726
rect 338 723 341 766
rect 354 763 357 806
rect 370 793 373 916
rect 394 813 397 896
rect 394 793 397 806
rect 362 686 365 776
rect 402 736 405 886
rect 418 803 421 926
rect 402 733 409 736
rect 386 706 389 726
rect 354 683 365 686
rect 378 703 389 706
rect 338 623 341 636
rect 290 533 293 556
rect 298 533 301 606
rect 202 413 205 433
rect 234 413 237 513
rect 306 506 309 526
rect 298 503 309 506
rect 250 423 253 436
rect 178 393 181 406
rect 250 403 277 406
rect 250 346 253 403
rect 242 343 253 346
rect 162 296 165 336
rect 234 323 237 336
rect 242 323 245 343
rect 162 293 173 296
rect 170 203 173 293
rect 218 213 221 226
rect 250 223 253 336
rect 258 323 261 356
rect 266 306 269 326
rect 274 323 277 403
rect 282 353 285 416
rect 298 346 301 503
rect 298 343 309 346
rect 306 323 309 343
rect 314 333 317 616
rect 330 553 333 606
rect 338 593 341 616
rect 322 533 325 546
rect 346 536 349 646
rect 354 603 357 683
rect 378 646 381 703
rect 378 643 389 646
rect 362 603 365 626
rect 322 443 325 516
rect 330 413 333 536
rect 342 533 349 536
rect 362 533 365 546
rect 378 533 381 616
rect 386 613 389 643
rect 342 366 345 533
rect 354 403 357 526
rect 370 506 373 526
rect 386 516 389 606
rect 394 603 397 726
rect 406 666 409 733
rect 426 686 429 816
rect 402 663 409 666
rect 418 683 429 686
rect 402 643 405 663
rect 402 613 405 636
rect 366 503 373 506
rect 378 513 389 516
rect 394 513 397 526
rect 366 376 369 503
rect 378 403 381 513
rect 410 506 413 606
rect 418 586 421 683
rect 434 603 437 926
rect 446 886 449 983
rect 466 923 469 983
rect 446 883 453 886
rect 442 613 445 806
rect 450 723 453 883
rect 474 733 477 946
rect 514 933 517 946
rect 498 793 501 816
rect 506 686 509 886
rect 546 883 549 936
rect 594 923 597 946
rect 634 936 637 956
rect 610 933 637 936
rect 650 933 653 946
rect 610 876 613 933
rect 602 873 613 876
rect 546 803 549 816
rect 554 723 557 746
rect 506 683 525 686
rect 418 583 437 586
rect 402 503 413 506
rect 402 446 405 503
rect 386 413 389 446
rect 394 443 405 446
rect 366 373 373 376
rect 342 363 349 366
rect 266 303 277 306
rect 274 236 277 303
rect 266 233 277 236
rect 266 213 269 233
rect 322 203 325 346
rect 346 343 349 363
rect 346 323 349 336
rect 354 306 357 366
rect 350 303 357 306
rect 350 206 353 303
rect 362 213 365 336
rect 370 323 373 373
rect 386 333 389 406
rect 394 403 397 443
rect 434 426 437 583
rect 482 573 485 606
rect 466 523 469 546
rect 514 533 517 576
rect 522 563 525 683
rect 602 636 605 873
rect 626 826 629 926
rect 634 913 637 926
rect 642 893 645 926
rect 658 903 661 926
rect 666 923 669 936
rect 674 913 677 936
rect 706 903 709 926
rect 666 826 669 896
rect 626 823 633 826
rect 618 773 621 816
rect 630 756 633 823
rect 658 823 669 826
rect 658 766 661 823
rect 674 793 677 816
rect 698 803 701 816
rect 658 763 669 766
rect 626 753 633 756
rect 602 633 613 636
rect 570 593 573 616
rect 586 613 605 616
rect 610 613 613 633
rect 418 423 437 426
rect 378 323 389 326
rect 402 213 405 416
rect 410 403 413 416
rect 418 403 421 423
rect 474 413 477 526
rect 530 523 533 536
rect 586 533 589 613
rect 586 513 589 526
rect 594 523 597 606
rect 626 603 629 753
rect 658 733 661 746
rect 634 723 653 726
rect 666 723 669 763
rect 674 733 677 756
rect 682 733 685 776
rect 682 706 685 726
rect 674 703 685 706
rect 674 636 677 703
rect 674 633 685 636
rect 602 523 605 536
rect 610 513 613 526
rect 530 413 533 426
rect 618 423 621 536
rect 642 483 645 616
rect 658 573 661 606
rect 666 603 669 616
rect 682 613 685 633
rect 674 593 677 606
rect 666 533 669 566
rect 650 503 653 526
rect 626 423 653 426
rect 626 413 629 423
rect 554 366 557 406
rect 546 363 557 366
rect 350 203 357 206
rect 322 123 325 196
rect 354 123 357 203
rect 410 193 413 206
rect 402 133 405 146
rect 434 133 437 336
rect 482 323 485 356
rect 530 323 533 336
rect 546 256 549 363
rect 570 333 573 406
rect 594 323 597 346
rect 626 323 629 406
rect 634 333 637 416
rect 650 413 653 423
rect 642 306 645 406
rect 650 346 653 366
rect 658 353 661 406
rect 650 343 661 346
rect 658 333 661 343
rect 634 303 645 306
rect 650 323 661 326
rect 546 253 557 256
rect 474 213 477 236
rect 490 163 493 206
rect 538 193 541 216
rect 554 176 557 253
rect 634 236 637 303
rect 634 233 645 236
rect 650 233 653 323
rect 594 213 597 226
rect 546 173 557 176
rect 482 123 485 156
rect 530 123 533 136
rect 546 133 549 173
rect 554 163 557 173
rect 594 133 597 206
rect 634 183 637 216
rect 642 176 645 233
rect 650 213 653 226
rect 658 193 661 206
rect 666 196 669 436
rect 674 403 677 486
rect 682 243 685 496
rect 690 413 693 506
rect 698 493 701 756
rect 714 603 717 1036
rect 730 1013 733 1133
rect 730 813 733 946
rect 754 943 757 1136
rect 762 1013 765 1026
rect 770 953 773 1006
rect 786 1003 789 1173
rect 802 1086 805 1126
rect 802 1083 813 1086
rect 802 966 805 1016
rect 810 1003 813 1083
rect 826 1023 829 1206
rect 874 1156 877 1176
rect 858 1153 877 1156
rect 834 1106 837 1126
rect 834 1103 845 1106
rect 842 1036 845 1103
rect 858 1046 861 1153
rect 858 1043 877 1046
rect 834 1033 845 1036
rect 802 963 809 966
rect 778 923 781 946
rect 738 813 741 836
rect 746 793 749 806
rect 754 776 757 816
rect 762 803 765 886
rect 770 803 773 906
rect 778 836 781 856
rect 778 833 785 836
rect 782 776 785 833
rect 794 806 797 956
rect 806 856 809 963
rect 802 853 809 856
rect 802 833 805 853
rect 810 813 813 826
rect 794 803 805 806
rect 818 803 821 1016
rect 826 976 829 1006
rect 834 1003 837 1033
rect 842 1003 845 1016
rect 858 1013 861 1026
rect 866 1006 869 1016
rect 850 1003 869 1006
rect 826 973 837 976
rect 826 876 829 926
rect 834 883 837 973
rect 850 933 853 946
rect 826 873 837 876
rect 746 773 757 776
rect 778 773 785 776
rect 730 566 733 606
rect 738 603 741 736
rect 746 723 749 773
rect 778 756 781 773
rect 762 753 781 756
rect 754 713 757 726
rect 746 613 757 616
rect 730 563 737 566
rect 690 203 693 406
rect 698 306 701 416
rect 706 403 709 526
rect 714 523 717 546
rect 734 486 737 563
rect 746 523 749 606
rect 754 523 757 613
rect 762 506 765 753
rect 778 733 781 746
rect 770 686 773 726
rect 786 703 789 726
rect 794 723 797 736
rect 802 713 805 803
rect 826 703 829 806
rect 834 803 837 873
rect 842 866 845 926
rect 842 863 853 866
rect 850 733 853 863
rect 858 833 861 926
rect 874 916 877 1043
rect 870 913 877 916
rect 870 846 873 913
rect 882 853 885 1146
rect 898 1056 901 1393
rect 922 1323 925 1403
rect 938 1243 941 1836
rect 946 1813 949 2096
rect 970 2033 973 2156
rect 986 2083 989 2226
rect 1010 2213 1013 2233
rect 1018 2196 1021 2306
rect 1010 2193 1021 2196
rect 1010 2116 1013 2193
rect 994 2063 997 2116
rect 1010 2113 1021 2116
rect 1018 2093 1021 2113
rect 978 1976 981 2006
rect 1002 2003 1005 2086
rect 1026 2056 1029 2423
rect 1034 2403 1037 2546
rect 1042 2503 1045 2593
rect 1058 2523 1061 2706
rect 1082 2646 1085 2773
rect 1106 2736 1109 2873
rect 1138 2813 1141 2916
rect 1122 2766 1125 2786
rect 1122 2763 1133 2766
rect 1098 2733 1109 2736
rect 1098 2666 1101 2733
rect 1098 2663 1109 2666
rect 1082 2643 1093 2646
rect 1066 2443 1069 2626
rect 1042 2413 1045 2436
rect 1058 2423 1069 2426
rect 1050 2413 1069 2416
rect 1074 2403 1077 2546
rect 1090 2536 1093 2643
rect 1106 2623 1109 2663
rect 1082 2533 1093 2536
rect 1082 2506 1085 2526
rect 1082 2503 1089 2506
rect 1086 2396 1089 2503
rect 1098 2413 1101 2536
rect 1106 2523 1109 2536
rect 1114 2516 1117 2726
rect 1130 2646 1133 2763
rect 1154 2723 1157 2906
rect 1186 2903 1189 2926
rect 1170 2776 1173 2806
rect 1194 2783 1197 2916
rect 1170 2773 1181 2776
rect 1178 2733 1181 2773
rect 1186 2666 1189 2686
rect 1110 2513 1117 2516
rect 1122 2643 1133 2646
rect 1182 2663 1189 2666
rect 1110 2426 1113 2513
rect 1106 2423 1113 2426
rect 1082 2393 1089 2396
rect 1034 2333 1045 2336
rect 1066 2333 1069 2346
rect 1042 2256 1045 2333
rect 1058 2303 1061 2326
rect 1066 2313 1069 2326
rect 1042 2253 1049 2256
rect 1034 2223 1037 2246
rect 1034 2103 1037 2206
rect 1046 2136 1049 2253
rect 1058 2213 1061 2236
rect 1074 2233 1077 2326
rect 1042 2133 1049 2136
rect 1042 2083 1045 2133
rect 1066 2116 1069 2136
rect 1022 2053 1029 2056
rect 1010 2013 1013 2026
rect 978 1973 989 1976
rect 962 1923 965 1936
rect 986 1856 989 1973
rect 1022 1956 1025 2053
rect 1022 1953 1029 1956
rect 1002 1923 1005 1936
rect 1018 1906 1021 1936
rect 962 1853 989 1856
rect 1010 1903 1021 1906
rect 1010 1856 1013 1903
rect 1010 1853 1021 1856
rect 946 1676 949 1796
rect 962 1723 965 1853
rect 1018 1833 1021 1853
rect 946 1673 957 1676
rect 954 1556 957 1673
rect 986 1653 989 1806
rect 1018 1763 1021 1806
rect 978 1613 981 1626
rect 994 1556 997 1726
rect 1010 1713 1013 1726
rect 1018 1566 1021 1636
rect 946 1553 957 1556
rect 986 1553 997 1556
rect 1010 1563 1021 1566
rect 946 1386 949 1553
rect 986 1533 989 1553
rect 954 1476 957 1526
rect 954 1473 965 1476
rect 962 1426 965 1473
rect 954 1423 965 1426
rect 954 1403 957 1423
rect 946 1383 965 1386
rect 962 1266 965 1383
rect 954 1263 965 1266
rect 922 1133 925 1206
rect 954 1196 957 1263
rect 986 1256 989 1436
rect 1010 1426 1013 1563
rect 1010 1423 1021 1426
rect 994 1316 997 1336
rect 994 1313 1005 1316
rect 1010 1313 1013 1406
rect 1018 1396 1021 1423
rect 1026 1413 1029 1953
rect 1034 1633 1037 1956
rect 1034 1603 1037 1616
rect 1042 1433 1045 2046
rect 1050 1773 1053 2116
rect 1062 2113 1069 2116
rect 1062 2046 1065 2113
rect 1074 2056 1077 2226
rect 1082 2186 1085 2393
rect 1090 2286 1093 2346
rect 1106 2303 1109 2423
rect 1122 2406 1125 2643
rect 1182 2596 1185 2663
rect 1194 2603 1197 2636
rect 1130 2576 1133 2596
rect 1182 2593 1189 2596
rect 1130 2573 1137 2576
rect 1134 2446 1137 2573
rect 1178 2513 1181 2526
rect 1118 2403 1125 2406
rect 1130 2443 1137 2446
rect 1118 2286 1121 2403
rect 1090 2283 1101 2286
rect 1098 2226 1101 2283
rect 1090 2223 1101 2226
rect 1114 2283 1121 2286
rect 1090 2203 1093 2223
rect 1082 2183 1089 2186
rect 1086 2096 1089 2183
rect 1114 2146 1117 2283
rect 1130 2266 1133 2443
rect 1146 2433 1149 2506
rect 1162 2433 1165 2446
rect 1138 2406 1141 2426
rect 1170 2423 1173 2436
rect 1178 2416 1181 2506
rect 1186 2503 1189 2593
rect 1194 2503 1197 2516
rect 1202 2486 1205 2756
rect 1210 2656 1213 2916
rect 1234 2866 1237 2993
rect 1258 2923 1261 3006
rect 1258 2903 1261 2916
rect 1266 2903 1269 2996
rect 1278 2936 1281 3103
rect 1318 3076 1321 3163
rect 1330 3123 1333 3206
rect 1338 3203 1341 3313
rect 1314 3073 1321 3076
rect 1290 2976 1293 3026
rect 1314 2993 1317 3073
rect 1322 3033 1325 3046
rect 1338 3033 1341 3116
rect 1346 3026 1349 3126
rect 1354 3103 1357 3453
rect 1386 3433 1389 3526
rect 1394 3416 1397 3446
rect 1402 3436 1405 3536
rect 1410 3443 1413 3586
rect 1418 3573 1421 3606
rect 1426 3603 1429 3616
rect 1402 3433 1413 3436
rect 1390 3413 1397 3416
rect 1378 3323 1381 3346
rect 1390 3326 1393 3413
rect 1402 3333 1405 3426
rect 1410 3413 1413 3433
rect 1442 3403 1445 3526
rect 1482 3523 1485 3546
rect 1490 3466 1493 3736
rect 1514 3733 1517 3806
rect 1538 3793 1541 3806
rect 1562 3743 1565 3806
rect 1546 3646 1549 3736
rect 1538 3643 1549 3646
rect 1522 3593 1525 3616
rect 1538 3596 1541 3643
rect 1538 3593 1549 3596
rect 1490 3463 1501 3466
rect 1450 3413 1453 3426
rect 1426 3333 1429 3386
rect 1442 3366 1445 3386
rect 1482 3383 1485 3456
rect 1442 3363 1449 3366
rect 1390 3323 1397 3326
rect 1370 3213 1373 3256
rect 1378 3193 1381 3206
rect 1386 3183 1389 3226
rect 1394 3163 1397 3323
rect 1426 3276 1429 3326
rect 1446 3306 1449 3363
rect 1498 3356 1501 3463
rect 1530 3453 1533 3546
rect 1546 3506 1549 3593
rect 1570 3543 1573 3796
rect 1582 3766 1585 3853
rect 1618 3813 1621 3863
rect 1582 3763 1589 3766
rect 1578 3723 1581 3746
rect 1586 3743 1589 3763
rect 1586 3613 1589 3736
rect 1602 3733 1605 3746
rect 1626 3733 1629 3936
rect 1634 3923 1637 4006
rect 1646 4003 1653 4006
rect 1634 3733 1637 3906
rect 1646 3756 1649 4003
rect 1646 3753 1653 3756
rect 1610 3723 1621 3726
rect 1610 3613 1613 3716
rect 1634 3713 1637 3726
rect 1642 3723 1645 3736
rect 1570 3523 1573 3536
rect 1546 3503 1557 3506
rect 1554 3436 1557 3503
rect 1586 3443 1589 3606
rect 1546 3433 1557 3436
rect 1522 3366 1525 3406
rect 1546 3373 1549 3433
rect 1594 3426 1597 3536
rect 1602 3496 1605 3526
rect 1618 3513 1621 3616
rect 1634 3603 1637 3616
rect 1634 3533 1637 3596
rect 1642 3533 1645 3716
rect 1650 3593 1653 3753
rect 1658 3713 1661 4076
rect 1666 4013 1669 4126
rect 1674 4096 1677 4173
rect 1674 4093 1685 4096
rect 1682 4006 1685 4093
rect 1674 4003 1685 4006
rect 1674 3946 1677 4003
rect 1666 3943 1677 3946
rect 1698 3943 1701 4196
rect 1714 4193 1717 4206
rect 1722 4123 1725 4216
rect 1730 4173 1733 4326
rect 1738 4313 1741 4326
rect 1746 4213 1749 4446
rect 1754 4403 1757 4556
rect 1762 4523 1765 4573
rect 1778 4443 1781 4526
rect 1786 4516 1789 4616
rect 1818 4613 1821 4626
rect 1794 4533 1797 4606
rect 1866 4593 1869 4606
rect 1818 4533 1821 4556
rect 1786 4513 1797 4516
rect 1810 4513 1813 4526
rect 1794 4436 1797 4513
rect 1762 4346 1765 4426
rect 1754 4343 1765 4346
rect 1754 4166 1757 4343
rect 1762 4213 1765 4336
rect 1770 4316 1773 4406
rect 1778 4396 1781 4436
rect 1786 4433 1797 4436
rect 1786 4403 1789 4433
rect 1778 4393 1789 4396
rect 1786 4333 1789 4393
rect 1794 4323 1797 4416
rect 1802 4343 1805 4406
rect 1770 4313 1777 4316
rect 1774 4236 1777 4313
rect 1770 4233 1777 4236
rect 1762 4196 1765 4206
rect 1770 4203 1773 4233
rect 1786 4213 1789 4236
rect 1762 4193 1773 4196
rect 1754 4163 1765 4166
rect 1666 3803 1669 3943
rect 1674 3913 1677 3936
rect 1690 3903 1693 3936
rect 1698 3886 1701 3926
rect 1690 3883 1701 3886
rect 1690 3836 1693 3883
rect 1690 3833 1701 3836
rect 1698 3813 1701 3833
rect 1706 3766 1709 3956
rect 1714 3923 1717 4016
rect 1730 3996 1733 4006
rect 1738 4003 1741 4016
rect 1746 3996 1749 4016
rect 1730 3993 1749 3996
rect 1730 3913 1733 3926
rect 1730 3793 1733 3806
rect 1746 3773 1749 3946
rect 1754 3923 1757 4006
rect 1762 3883 1765 4163
rect 1770 3996 1773 4193
rect 1778 4116 1781 4206
rect 1794 4203 1797 4246
rect 1786 4133 1789 4176
rect 1802 4156 1805 4336
rect 1810 4323 1813 4416
rect 1818 4403 1821 4526
rect 1826 4513 1829 4526
rect 1826 4333 1829 4426
rect 1834 4403 1837 4546
rect 1842 4423 1845 4526
rect 1882 4523 1885 4616
rect 1922 4533 1925 4546
rect 1850 4453 1861 4456
rect 1850 4416 1853 4453
rect 1842 4413 1853 4416
rect 1842 4393 1845 4413
rect 1850 4336 1853 4406
rect 1858 4403 1861 4416
rect 1890 4403 1893 4416
rect 1898 4413 1901 4526
rect 1938 4503 1941 4646
rect 1994 4636 1997 4683
rect 1994 4633 2005 4636
rect 1946 4613 1949 4626
rect 1986 4613 1989 4626
rect 1906 4413 1909 4436
rect 1938 4396 1941 4406
rect 1946 4403 1949 4556
rect 1954 4523 1957 4596
rect 1970 4543 1973 4606
rect 1986 4593 1989 4606
rect 2002 4586 2005 4633
rect 2226 4626 2229 4740
rect 3682 4726 3685 4740
rect 3674 4723 3685 4726
rect 2314 4646 2317 4686
rect 3674 4666 3677 4723
rect 3698 4676 3701 4740
rect 3698 4673 3709 4676
rect 3674 4663 3685 4666
rect 2306 4643 2317 4646
rect 2226 4623 2233 4626
rect 1994 4583 2005 4586
rect 1962 4523 1965 4536
rect 1978 4533 1981 4556
rect 1954 4396 1957 4416
rect 1962 4403 1965 4426
rect 1938 4393 1957 4396
rect 1850 4333 1861 4336
rect 1938 4333 1941 4366
rect 1810 4213 1813 4226
rect 1818 4203 1821 4216
rect 1834 4213 1837 4246
rect 1794 4153 1805 4156
rect 1778 4113 1785 4116
rect 1782 4036 1785 4113
rect 1778 4033 1785 4036
rect 1778 4013 1781 4033
rect 1794 4003 1797 4153
rect 1802 4123 1805 4146
rect 1810 4133 1829 4136
rect 1842 4133 1845 4326
rect 1858 4286 1861 4333
rect 1914 4313 1917 4326
rect 1954 4313 1957 4326
rect 1850 4283 1861 4286
rect 1850 4216 1853 4283
rect 1850 4213 1861 4216
rect 1850 4133 1853 4206
rect 1810 4106 1813 4133
rect 1806 4103 1813 4106
rect 1806 4006 1809 4103
rect 1818 4013 1821 4126
rect 1834 4116 1837 4126
rect 1858 4123 1861 4213
rect 1866 4203 1869 4266
rect 1834 4113 1845 4116
rect 1834 4096 1837 4113
rect 1874 4106 1877 4236
rect 1914 4226 1917 4246
rect 1906 4223 1917 4226
rect 1882 4193 1885 4216
rect 1890 4203 1893 4216
rect 1906 4156 1909 4223
rect 1906 4153 1917 4156
rect 1866 4103 1877 4106
rect 1834 4093 1845 4096
rect 1842 4036 1845 4093
rect 1866 4046 1869 4103
rect 1890 4053 1893 4126
rect 1866 4043 1877 4046
rect 1834 4033 1845 4036
rect 1834 4013 1837 4033
rect 1806 4003 1813 4006
rect 1770 3993 1781 3996
rect 1778 3946 1781 3993
rect 1770 3943 1781 3946
rect 1770 3923 1773 3943
rect 1666 3733 1669 3766
rect 1706 3763 1717 3766
rect 1674 3723 1685 3726
rect 1714 3686 1717 3763
rect 1754 3733 1757 3796
rect 1770 3793 1773 3816
rect 1794 3813 1797 3926
rect 1730 3713 1733 3726
rect 1770 3713 1773 3726
rect 1778 3696 1781 3776
rect 1706 3683 1717 3686
rect 1770 3693 1781 3696
rect 1658 3606 1661 3626
rect 1658 3603 1669 3606
rect 1666 3546 1669 3603
rect 1602 3493 1613 3496
rect 1610 3436 1613 3493
rect 1590 3423 1597 3426
rect 1602 3433 1613 3436
rect 1570 3393 1573 3416
rect 1522 3363 1541 3366
rect 1490 3353 1501 3356
rect 1458 3313 1461 3326
rect 1418 3273 1429 3276
rect 1442 3303 1449 3306
rect 1418 3186 1421 3273
rect 1442 3203 1445 3303
rect 1466 3193 1469 3216
rect 1418 3183 1429 3186
rect 1418 3123 1421 3136
rect 1370 3043 1373 3116
rect 1330 3013 1333 3026
rect 1338 3023 1349 3026
rect 1290 2973 1301 2976
rect 1274 2933 1281 2936
rect 1234 2863 1245 2866
rect 1218 2803 1221 2816
rect 1242 2766 1245 2863
rect 1242 2763 1249 2766
rect 1218 2676 1221 2746
rect 1226 2723 1229 2736
rect 1246 2686 1249 2763
rect 1242 2683 1249 2686
rect 1218 2673 1229 2676
rect 1210 2653 1217 2656
rect 1214 2546 1217 2653
rect 1162 2413 1181 2416
rect 1194 2483 1205 2486
rect 1210 2543 1217 2546
rect 1138 2403 1149 2406
rect 1146 2346 1149 2403
rect 1126 2263 1133 2266
rect 1138 2343 1149 2346
rect 1126 2166 1129 2263
rect 1126 2163 1133 2166
rect 1114 2143 1125 2146
rect 1082 2093 1089 2096
rect 1082 2073 1085 2093
rect 1074 2053 1085 2056
rect 1062 2043 1069 2046
rect 1058 1896 1061 2026
rect 1066 2013 1069 2043
rect 1082 2006 1085 2053
rect 1098 2016 1101 2136
rect 1114 2103 1117 2126
rect 1122 2043 1125 2143
rect 1130 2033 1133 2163
rect 1138 2133 1141 2343
rect 1162 2326 1165 2413
rect 1146 2303 1149 2326
rect 1162 2323 1169 2326
rect 1146 2213 1149 2226
rect 1138 2026 1141 2126
rect 1130 2023 1141 2026
rect 1146 2023 1149 2116
rect 1074 2003 1085 2006
rect 1094 2013 1101 2016
rect 1074 1953 1077 2003
rect 1094 1946 1097 2013
rect 1094 1943 1101 1946
rect 1074 1933 1085 1936
rect 1066 1913 1069 1926
rect 1074 1923 1085 1926
rect 1058 1893 1065 1896
rect 1062 1796 1065 1893
rect 1058 1793 1065 1796
rect 1050 1723 1053 1766
rect 1058 1656 1061 1793
rect 1066 1706 1069 1776
rect 1074 1723 1077 1923
rect 1090 1913 1093 1926
rect 1098 1896 1101 1943
rect 1090 1893 1101 1896
rect 1090 1786 1093 1893
rect 1106 1793 1109 2006
rect 1114 1923 1117 2016
rect 1122 2003 1125 2016
rect 1130 2013 1133 2023
rect 1138 2016 1141 2023
rect 1138 2013 1149 2016
rect 1130 1906 1133 1926
rect 1122 1903 1133 1906
rect 1122 1836 1125 1903
rect 1122 1833 1133 1836
rect 1090 1783 1101 1786
rect 1066 1703 1077 1706
rect 1058 1653 1065 1656
rect 1062 1576 1065 1653
rect 1058 1573 1065 1576
rect 1034 1413 1037 1426
rect 1042 1413 1053 1416
rect 1058 1413 1061 1573
rect 1018 1393 1025 1396
rect 1050 1393 1053 1413
rect 1074 1406 1077 1703
rect 1066 1403 1077 1406
rect 986 1253 993 1256
rect 970 1213 973 1236
rect 946 1193 957 1196
rect 946 1146 949 1193
rect 946 1143 957 1146
rect 954 1096 957 1143
rect 970 1123 973 1136
rect 990 1116 993 1253
rect 1002 1213 1005 1313
rect 1022 1306 1025 1393
rect 1018 1303 1025 1306
rect 1010 1186 1013 1206
rect 1002 1183 1013 1186
rect 1002 1123 1005 1183
rect 1018 1153 1021 1303
rect 1034 1286 1037 1356
rect 1030 1283 1037 1286
rect 1030 1176 1033 1283
rect 1030 1173 1037 1176
rect 1042 1173 1045 1386
rect 1066 1346 1069 1403
rect 1090 1383 1093 1746
rect 1098 1736 1101 1783
rect 1098 1733 1109 1736
rect 1098 1703 1101 1726
rect 1106 1646 1109 1733
rect 1114 1713 1117 1736
rect 1122 1723 1125 1796
rect 1130 1706 1133 1833
rect 1102 1643 1109 1646
rect 1126 1703 1133 1706
rect 1102 1416 1105 1643
rect 1102 1413 1109 1416
rect 1114 1413 1117 1636
rect 1126 1446 1129 1703
rect 1126 1443 1133 1446
rect 1130 1423 1133 1443
rect 1106 1396 1109 1413
rect 1050 1343 1069 1346
rect 1034 1143 1037 1173
rect 990 1113 1005 1116
rect 946 1093 957 1096
rect 898 1053 905 1056
rect 902 976 905 1053
rect 946 1033 949 1093
rect 898 973 905 976
rect 870 843 877 846
rect 770 683 789 686
rect 786 566 789 683
rect 730 483 737 486
rect 754 503 765 506
rect 778 563 789 566
rect 706 333 709 346
rect 714 323 717 336
rect 698 303 705 306
rect 702 226 705 303
rect 722 286 725 406
rect 730 403 733 483
rect 754 356 757 503
rect 778 466 781 563
rect 802 533 805 546
rect 802 506 805 526
rect 810 523 813 616
rect 818 533 821 576
rect 826 523 829 656
rect 842 636 845 726
rect 858 703 861 726
rect 866 653 869 826
rect 874 753 877 843
rect 890 833 893 846
rect 882 813 885 826
rect 898 823 901 973
rect 914 933 917 1016
rect 906 813 909 836
rect 874 713 877 726
rect 838 633 845 636
rect 838 586 841 633
rect 838 583 845 586
rect 770 463 781 466
rect 794 503 805 506
rect 770 413 773 463
rect 794 446 797 503
rect 778 413 781 446
rect 794 443 805 446
rect 754 353 765 356
rect 730 333 741 336
rect 698 223 705 226
rect 714 283 725 286
rect 666 193 677 196
rect 698 193 701 223
rect 714 206 717 283
rect 730 256 733 326
rect 722 253 733 256
rect 722 213 725 253
rect 738 213 741 306
rect 642 173 653 176
rect 594 113 597 126
rect 642 123 645 146
rect 650 133 653 173
rect 658 123 661 186
rect 666 133 669 156
rect 674 123 677 193
rect 682 123 685 136
rect 690 133 693 146
rect 706 143 709 206
rect 714 203 725 206
rect 722 133 725 203
rect 730 126 733 206
rect 746 203 749 226
rect 714 123 733 126
rect 738 113 741 136
rect 746 123 749 196
rect 754 73 757 146
rect 762 103 765 353
rect 770 323 773 396
rect 778 323 781 336
rect 786 213 789 406
rect 794 403 797 426
rect 802 413 805 443
rect 810 403 813 516
rect 794 303 797 316
rect 802 213 805 386
rect 818 213 821 506
rect 826 393 829 426
rect 834 376 837 436
rect 842 413 845 583
rect 858 563 861 606
rect 882 533 885 616
rect 890 613 893 736
rect 906 656 909 806
rect 922 733 925 1026
rect 930 883 933 986
rect 946 976 949 1006
rect 962 1003 973 1006
rect 962 976 965 996
rect 946 973 965 976
rect 970 973 973 1003
rect 962 933 965 973
rect 914 703 917 726
rect 922 723 933 726
rect 938 716 941 856
rect 954 803 957 906
rect 986 903 989 926
rect 962 813 981 816
rect 970 733 973 746
rect 978 733 981 813
rect 986 793 989 886
rect 994 833 997 1016
rect 930 713 941 716
rect 902 653 909 656
rect 902 546 905 653
rect 930 626 933 713
rect 970 696 973 716
rect 926 623 933 626
rect 962 693 973 696
rect 926 576 929 623
rect 914 573 929 576
rect 902 543 909 546
rect 874 513 877 526
rect 890 523 893 536
rect 898 513 901 526
rect 906 506 909 543
rect 898 503 909 506
rect 890 476 893 496
rect 882 473 893 476
rect 866 413 869 436
rect 882 416 885 473
rect 898 423 901 503
rect 914 496 917 573
rect 938 533 941 616
rect 962 546 965 693
rect 986 676 989 726
rect 994 713 997 736
rect 978 673 989 676
rect 978 566 981 673
rect 994 656 997 706
rect 990 653 997 656
rect 990 586 993 653
rect 990 583 997 586
rect 978 563 989 566
rect 962 543 973 546
rect 970 523 973 543
rect 986 526 989 563
rect 978 523 989 526
rect 994 523 997 583
rect 906 493 917 496
rect 882 413 893 416
rect 830 373 837 376
rect 830 316 833 373
rect 842 323 845 406
rect 830 313 837 316
rect 834 223 837 313
rect 850 273 853 306
rect 882 213 885 336
rect 890 313 893 413
rect 906 393 909 493
rect 914 353 917 416
rect 922 213 925 406
rect 930 343 933 416
rect 938 373 941 406
rect 946 383 949 516
rect 978 506 981 523
rect 1002 516 1005 1113
rect 1010 876 1013 986
rect 1018 963 1021 1136
rect 1042 936 1045 1156
rect 1050 983 1053 1343
rect 1058 1303 1061 1326
rect 1058 1106 1061 1256
rect 1066 1233 1069 1336
rect 1074 1313 1077 1326
rect 1066 1213 1069 1226
rect 1074 1213 1077 1306
rect 1082 1293 1085 1336
rect 1090 1213 1093 1336
rect 1098 1323 1101 1396
rect 1106 1393 1113 1396
rect 1138 1393 1141 2006
rect 1146 2003 1149 2013
rect 1146 1913 1149 1936
rect 1146 1716 1149 1856
rect 1154 1823 1157 2316
rect 1166 2056 1169 2323
rect 1162 2053 1169 2056
rect 1162 1816 1165 2053
rect 1170 1853 1173 2036
rect 1178 1876 1181 2406
rect 1194 2336 1197 2483
rect 1210 2403 1213 2543
rect 1226 2526 1229 2673
rect 1242 2593 1245 2683
rect 1226 2523 1237 2526
rect 1218 2386 1221 2426
rect 1234 2393 1237 2523
rect 1250 2466 1253 2556
rect 1258 2523 1261 2856
rect 1274 2846 1277 2933
rect 1282 2903 1285 2916
rect 1298 2876 1301 2973
rect 1270 2843 1277 2846
rect 1290 2873 1301 2876
rect 1270 2706 1273 2843
rect 1282 2716 1285 2836
rect 1290 2806 1293 2873
rect 1298 2813 1301 2826
rect 1306 2813 1309 2856
rect 1322 2813 1325 3006
rect 1338 2993 1341 3023
rect 1346 3003 1349 3016
rect 1354 2986 1357 3036
rect 1378 3013 1381 3116
rect 1394 3063 1397 3106
rect 1410 3053 1413 3116
rect 1426 3033 1429 3183
rect 1474 3133 1477 3336
rect 1490 3333 1493 3353
rect 1514 3323 1517 3346
rect 1538 3236 1541 3363
rect 1590 3346 1593 3423
rect 1602 3413 1605 3433
rect 1650 3406 1653 3546
rect 1658 3543 1669 3546
rect 1658 3513 1661 3543
rect 1674 3513 1677 3526
rect 1690 3516 1693 3536
rect 1686 3513 1693 3516
rect 1658 3413 1661 3446
rect 1590 3343 1597 3346
rect 1554 3313 1557 3336
rect 1594 3323 1597 3343
rect 1602 3306 1605 3366
rect 1626 3333 1629 3346
rect 1610 3313 1613 3326
rect 1522 3233 1541 3236
rect 1594 3303 1605 3306
rect 1338 2983 1357 2986
rect 1338 2876 1341 2983
rect 1330 2873 1341 2876
rect 1290 2803 1301 2806
rect 1306 2803 1317 2806
rect 1282 2713 1289 2716
rect 1270 2703 1277 2706
rect 1274 2683 1277 2703
rect 1286 2666 1289 2713
rect 1282 2663 1289 2666
rect 1282 2643 1285 2663
rect 1290 2613 1293 2626
rect 1266 2563 1269 2606
rect 1282 2603 1293 2606
rect 1298 2586 1301 2803
rect 1294 2583 1301 2586
rect 1250 2463 1261 2466
rect 1258 2406 1261 2463
rect 1266 2413 1269 2536
rect 1274 2523 1285 2526
rect 1282 2513 1285 2523
rect 1294 2466 1297 2583
rect 1306 2533 1309 2726
rect 1314 2693 1317 2736
rect 1322 2686 1325 2766
rect 1318 2683 1325 2686
rect 1318 2546 1321 2683
rect 1330 2593 1333 2873
rect 1338 2813 1341 2856
rect 1346 2806 1349 2846
rect 1362 2816 1365 2986
rect 1338 2803 1349 2806
rect 1358 2813 1365 2816
rect 1338 2733 1341 2803
rect 1358 2756 1361 2813
rect 1358 2753 1365 2756
rect 1346 2733 1357 2736
rect 1362 2726 1365 2753
rect 1338 2713 1341 2726
rect 1346 2703 1349 2726
rect 1354 2723 1365 2726
rect 1370 2723 1373 2806
rect 1378 2753 1381 2866
rect 1354 2713 1357 2723
rect 1314 2543 1321 2546
rect 1294 2463 1301 2466
rect 1258 2403 1269 2406
rect 1194 2333 1201 2336
rect 1186 2086 1189 2316
rect 1198 2246 1201 2333
rect 1198 2243 1205 2246
rect 1194 2093 1197 2226
rect 1202 2086 1205 2243
rect 1210 2236 1213 2386
rect 1218 2383 1229 2386
rect 1226 2323 1229 2383
rect 1226 2283 1229 2306
rect 1234 2303 1237 2376
rect 1250 2363 1253 2396
rect 1266 2346 1269 2403
rect 1254 2343 1269 2346
rect 1242 2303 1245 2316
rect 1254 2296 1257 2343
rect 1250 2293 1257 2296
rect 1218 2256 1221 2276
rect 1218 2253 1229 2256
rect 1210 2233 1217 2236
rect 1214 2166 1217 2233
rect 1210 2163 1217 2166
rect 1210 2103 1213 2163
rect 1226 2146 1229 2253
rect 1218 2143 1229 2146
rect 1218 2123 1221 2143
rect 1234 2113 1237 2126
rect 1186 2083 1197 2086
rect 1202 2083 1213 2086
rect 1194 2026 1197 2083
rect 1194 2023 1201 2026
rect 1186 1893 1189 2016
rect 1198 1976 1201 2023
rect 1194 1973 1201 1976
rect 1194 1926 1197 1973
rect 1210 1956 1213 2083
rect 1226 2013 1229 2096
rect 1250 2026 1253 2293
rect 1274 2213 1277 2396
rect 1298 2366 1301 2463
rect 1290 2363 1301 2366
rect 1290 2236 1293 2363
rect 1306 2346 1309 2506
rect 1302 2343 1309 2346
rect 1302 2256 1305 2343
rect 1302 2253 1309 2256
rect 1290 2233 1301 2236
rect 1306 2233 1309 2253
rect 1298 2216 1301 2233
rect 1314 2226 1317 2543
rect 1322 2413 1325 2526
rect 1330 2513 1333 2526
rect 1338 2403 1341 2626
rect 1346 2583 1349 2696
rect 1378 2686 1381 2746
rect 1386 2743 1389 3026
rect 1402 3013 1413 3016
rect 1418 3013 1421 3026
rect 1434 3023 1437 3106
rect 1466 3103 1469 3126
rect 1498 3073 1501 3126
rect 1506 3066 1509 3176
rect 1522 3103 1525 3233
rect 1594 3226 1597 3303
rect 1530 3206 1533 3216
rect 1538 3213 1541 3226
rect 1594 3223 1605 3226
rect 1530 3203 1549 3206
rect 1546 3146 1549 3186
rect 1578 3163 1581 3206
rect 1602 3176 1605 3223
rect 1610 3213 1613 3226
rect 1618 3213 1621 3326
rect 1634 3313 1637 3326
rect 1634 3213 1637 3226
rect 1594 3173 1605 3176
rect 1546 3143 1557 3146
rect 1554 3096 1557 3143
rect 1570 3123 1573 3146
rect 1498 3063 1509 3066
rect 1546 3093 1557 3096
rect 1442 3013 1445 3036
rect 1402 3003 1413 3006
rect 1442 2983 1445 3006
rect 1410 2816 1413 2926
rect 1474 2903 1477 2936
rect 1490 2926 1493 3016
rect 1482 2923 1493 2926
rect 1482 2886 1485 2923
rect 1498 2916 1501 3063
rect 1506 3013 1509 3026
rect 1514 3013 1525 3016
rect 1506 2923 1509 2996
rect 1402 2813 1413 2816
rect 1466 2883 1485 2886
rect 1490 2913 1501 2916
rect 1394 2733 1397 2806
rect 1410 2793 1413 2806
rect 1466 2786 1469 2883
rect 1466 2783 1485 2786
rect 1482 2763 1485 2783
rect 1362 2683 1381 2686
rect 1362 2603 1365 2683
rect 1410 2656 1413 2746
rect 1426 2733 1429 2746
rect 1450 2723 1453 2736
rect 1402 2653 1413 2656
rect 1386 2603 1389 2616
rect 1354 2506 1357 2526
rect 1350 2503 1357 2506
rect 1350 2436 1353 2503
rect 1350 2433 1357 2436
rect 1322 2323 1325 2336
rect 1330 2273 1333 2326
rect 1314 2223 1325 2226
rect 1282 2116 1285 2136
rect 1274 2113 1285 2116
rect 1274 2036 1277 2113
rect 1274 2033 1285 2036
rect 1250 2023 1261 2026
rect 1202 1953 1213 1956
rect 1202 1933 1205 1953
rect 1226 1926 1229 1946
rect 1194 1923 1205 1926
rect 1210 1923 1221 1926
rect 1226 1923 1233 1926
rect 1242 1923 1245 2016
rect 1258 1966 1261 2023
rect 1282 2013 1285 2033
rect 1274 1993 1277 2006
rect 1290 1983 1293 2216
rect 1298 2213 1309 2216
rect 1306 2206 1309 2213
rect 1298 2113 1301 2206
rect 1306 2203 1317 2206
rect 1306 2106 1309 2146
rect 1298 2103 1309 2106
rect 1250 1963 1261 1966
rect 1250 1943 1253 1963
rect 1250 1933 1269 1936
rect 1202 1896 1205 1916
rect 1198 1893 1205 1896
rect 1178 1873 1189 1876
rect 1154 1813 1165 1816
rect 1154 1733 1157 1746
rect 1170 1736 1173 1816
rect 1166 1733 1173 1736
rect 1146 1713 1153 1716
rect 1150 1586 1153 1713
rect 1166 1656 1169 1733
rect 1186 1726 1189 1873
rect 1198 1736 1201 1893
rect 1210 1813 1213 1923
rect 1198 1733 1205 1736
rect 1210 1733 1213 1796
rect 1178 1723 1189 1726
rect 1166 1653 1173 1656
rect 1162 1613 1165 1636
rect 1170 1616 1173 1653
rect 1178 1626 1181 1723
rect 1202 1716 1205 1733
rect 1202 1713 1209 1716
rect 1194 1633 1197 1706
rect 1206 1636 1209 1713
rect 1218 1696 1221 1916
rect 1230 1826 1233 1923
rect 1226 1823 1233 1826
rect 1226 1793 1229 1823
rect 1226 1713 1229 1736
rect 1234 1723 1237 1806
rect 1242 1803 1245 1876
rect 1250 1823 1253 1926
rect 1258 1803 1261 1906
rect 1266 1813 1269 1933
rect 1290 1903 1293 1926
rect 1298 1896 1301 2103
rect 1290 1893 1301 1896
rect 1274 1733 1277 1866
rect 1282 1793 1285 1816
rect 1282 1716 1285 1746
rect 1274 1713 1285 1716
rect 1218 1693 1229 1696
rect 1202 1633 1209 1636
rect 1178 1623 1197 1626
rect 1170 1613 1181 1616
rect 1162 1603 1173 1606
rect 1178 1586 1181 1613
rect 1150 1583 1157 1586
rect 1154 1506 1157 1583
rect 1146 1503 1157 1506
rect 1170 1583 1181 1586
rect 1146 1483 1149 1503
rect 1170 1436 1173 1583
rect 1186 1566 1189 1606
rect 1182 1563 1189 1566
rect 1182 1456 1185 1563
rect 1182 1453 1189 1456
rect 1170 1433 1181 1436
rect 1066 1123 1069 1146
rect 1082 1133 1085 1206
rect 1098 1203 1101 1296
rect 1110 1186 1113 1393
rect 1146 1356 1149 1426
rect 1154 1403 1165 1406
rect 1146 1353 1157 1356
rect 1106 1183 1113 1186
rect 1106 1166 1109 1183
rect 1098 1163 1109 1166
rect 1058 1103 1065 1106
rect 1062 1036 1065 1103
rect 1058 1033 1065 1036
rect 1034 933 1045 936
rect 1010 873 1021 876
rect 1018 756 1021 873
rect 994 513 1005 516
rect 1010 753 1021 756
rect 1010 513 1013 753
rect 1034 746 1037 933
rect 1050 906 1053 926
rect 1046 903 1053 906
rect 1046 836 1049 903
rect 1058 853 1061 1033
rect 1066 993 1069 1016
rect 1098 976 1101 1163
rect 1114 1096 1117 1156
rect 1110 1093 1117 1096
rect 1110 996 1113 1093
rect 1110 993 1117 996
rect 1098 973 1109 976
rect 1114 973 1117 993
rect 1046 833 1053 836
rect 1050 813 1053 833
rect 1058 813 1061 836
rect 1034 743 1045 746
rect 1018 696 1021 736
rect 1026 713 1029 726
rect 1018 693 1025 696
rect 1022 596 1025 693
rect 1018 593 1025 596
rect 1018 573 1021 593
rect 1034 533 1037 726
rect 1042 716 1045 743
rect 1050 736 1053 806
rect 1066 803 1069 906
rect 1074 883 1077 966
rect 1106 956 1109 973
rect 1106 953 1113 956
rect 1098 903 1101 926
rect 1110 876 1113 953
rect 1122 903 1125 1326
rect 1146 1323 1149 1346
rect 1154 1333 1157 1353
rect 1170 1253 1173 1416
rect 1178 1326 1181 1433
rect 1186 1353 1189 1453
rect 1194 1343 1197 1623
rect 1202 1406 1205 1633
rect 1210 1413 1213 1616
rect 1226 1566 1229 1693
rect 1274 1626 1277 1713
rect 1274 1623 1285 1626
rect 1282 1603 1285 1623
rect 1290 1586 1293 1893
rect 1306 1886 1309 1956
rect 1302 1883 1309 1886
rect 1302 1756 1305 1883
rect 1298 1753 1305 1756
rect 1298 1706 1301 1753
rect 1306 1723 1309 1736
rect 1298 1703 1305 1706
rect 1302 1636 1305 1703
rect 1298 1633 1305 1636
rect 1298 1596 1301 1633
rect 1306 1603 1309 1616
rect 1298 1593 1309 1596
rect 1218 1563 1229 1566
rect 1282 1583 1293 1586
rect 1202 1403 1213 1406
rect 1210 1383 1213 1403
rect 1218 1396 1221 1563
rect 1242 1533 1245 1546
rect 1226 1496 1229 1516
rect 1266 1513 1269 1526
rect 1226 1493 1237 1496
rect 1234 1436 1237 1493
rect 1282 1486 1285 1583
rect 1306 1503 1309 1593
rect 1226 1433 1237 1436
rect 1226 1403 1229 1433
rect 1258 1426 1261 1486
rect 1282 1483 1293 1486
rect 1258 1423 1269 1426
rect 1234 1413 1253 1416
rect 1218 1393 1229 1396
rect 1242 1393 1245 1406
rect 1178 1323 1189 1326
rect 1186 1266 1189 1323
rect 1202 1313 1205 1326
rect 1210 1316 1213 1336
rect 1226 1326 1229 1393
rect 1226 1323 1237 1326
rect 1210 1313 1217 1316
rect 1178 1263 1189 1266
rect 1178 1236 1181 1263
rect 1174 1233 1181 1236
rect 1214 1236 1217 1313
rect 1234 1266 1237 1323
rect 1226 1263 1237 1266
rect 1214 1233 1221 1236
rect 1138 1173 1141 1206
rect 1174 1166 1177 1233
rect 1186 1193 1189 1216
rect 1174 1163 1181 1166
rect 1130 1133 1133 1156
rect 1154 1133 1157 1146
rect 1178 1143 1181 1163
rect 1130 1123 1149 1126
rect 1138 1096 1141 1116
rect 1170 1103 1173 1136
rect 1178 1123 1181 1136
rect 1138 1093 1149 1096
rect 1146 1036 1149 1093
rect 1142 1033 1149 1036
rect 1130 973 1133 1006
rect 1142 886 1145 1033
rect 1154 1013 1173 1016
rect 1178 993 1181 1006
rect 1186 1003 1189 1126
rect 1138 883 1145 886
rect 1110 873 1117 876
rect 1074 813 1093 816
rect 1082 793 1085 806
rect 1098 786 1101 856
rect 1114 826 1117 873
rect 1106 823 1117 826
rect 1106 803 1109 823
rect 1090 783 1101 786
rect 1050 733 1061 736
rect 1042 713 1049 716
rect 1046 636 1049 713
rect 1042 633 1049 636
rect 978 503 989 506
rect 938 313 941 326
rect 962 323 965 426
rect 970 263 973 436
rect 986 413 989 503
rect 994 426 997 513
rect 1002 433 1005 506
rect 1042 493 1045 633
rect 1058 626 1061 733
rect 1058 623 1065 626
rect 1050 533 1053 616
rect 1062 506 1065 623
rect 1082 613 1085 736
rect 1090 733 1093 783
rect 1114 743 1133 746
rect 1098 733 1109 736
rect 1098 703 1101 726
rect 1058 503 1065 506
rect 1058 483 1061 503
rect 994 423 1005 426
rect 978 323 981 336
rect 986 333 989 346
rect 786 183 789 206
rect 802 133 805 146
rect 810 123 813 206
rect 818 133 821 156
rect 834 123 837 206
rect 962 173 965 206
rect 866 123 869 146
rect 914 133 917 166
rect 946 133 949 166
rect 994 153 997 206
rect 1002 163 1005 416
rect 1010 413 1013 446
rect 1010 393 1013 406
rect 1018 363 1021 416
rect 1026 323 1029 406
rect 1034 396 1037 416
rect 1050 396 1053 416
rect 1034 393 1053 396
rect 1034 343 1037 393
rect 1018 193 1021 216
rect 1042 213 1045 366
rect 994 123 997 136
rect 1026 133 1029 206
rect 1058 203 1061 216
rect 1042 123 1045 196
rect 1066 186 1069 436
rect 1074 306 1077 536
rect 1090 496 1093 546
rect 1098 523 1101 646
rect 1114 643 1117 743
rect 1122 723 1125 736
rect 1130 733 1133 743
rect 1138 726 1141 883
rect 1146 796 1149 816
rect 1154 803 1157 926
rect 1146 793 1157 796
rect 1154 733 1157 793
rect 1130 723 1141 726
rect 1130 683 1133 723
rect 1130 563 1133 676
rect 1146 633 1149 726
rect 1162 663 1165 986
rect 1194 963 1197 1126
rect 1202 1113 1205 1226
rect 1218 1213 1221 1233
rect 1226 1213 1229 1263
rect 1226 1126 1229 1146
rect 1210 1026 1213 1126
rect 1222 1123 1229 1126
rect 1222 1036 1225 1123
rect 1234 1113 1237 1126
rect 1222 1033 1229 1036
rect 1202 1023 1213 1026
rect 1202 983 1205 1023
rect 1122 533 1125 546
rect 1090 493 1101 496
rect 1098 436 1101 493
rect 1090 433 1101 436
rect 1090 413 1093 433
rect 1106 413 1117 416
rect 1082 323 1085 406
rect 1074 303 1081 306
rect 1078 186 1081 303
rect 1090 213 1093 336
rect 1098 313 1101 326
rect 1106 323 1109 413
rect 1114 193 1117 336
rect 1122 323 1125 526
rect 1146 523 1149 626
rect 1170 603 1173 946
rect 1186 913 1189 936
rect 1178 786 1181 906
rect 1210 896 1213 1016
rect 1206 893 1213 896
rect 1178 783 1185 786
rect 1182 656 1185 783
rect 1178 653 1185 656
rect 1178 566 1181 653
rect 1162 563 1181 566
rect 1162 486 1165 563
rect 1170 523 1173 546
rect 1154 483 1165 486
rect 1154 436 1157 483
rect 1178 466 1181 486
rect 1174 463 1181 466
rect 1154 433 1165 436
rect 1162 413 1165 433
rect 1174 376 1177 463
rect 1186 413 1189 636
rect 1194 626 1197 876
rect 1206 836 1209 893
rect 1202 833 1209 836
rect 1202 703 1205 833
rect 1210 713 1213 816
rect 1218 786 1221 1016
rect 1226 873 1229 1033
rect 1234 943 1237 1106
rect 1234 923 1237 936
rect 1218 783 1229 786
rect 1218 703 1221 726
rect 1194 623 1205 626
rect 1210 623 1213 696
rect 1194 413 1197 616
rect 1202 586 1205 623
rect 1218 613 1221 666
rect 1226 603 1229 783
rect 1234 673 1237 916
rect 1250 853 1253 1386
rect 1266 1356 1269 1423
rect 1258 1353 1269 1356
rect 1258 1296 1261 1353
rect 1266 1316 1269 1326
rect 1274 1323 1277 1336
rect 1290 1323 1293 1483
rect 1306 1333 1309 1416
rect 1266 1313 1277 1316
rect 1306 1313 1309 1326
rect 1258 1293 1265 1296
rect 1262 1226 1265 1293
rect 1258 1223 1265 1226
rect 1258 1093 1261 1223
rect 1274 1213 1277 1313
rect 1266 1193 1269 1206
rect 1282 1203 1285 1216
rect 1290 1213 1293 1246
rect 1266 1016 1269 1136
rect 1282 1123 1285 1156
rect 1290 1123 1293 1206
rect 1298 1203 1301 1236
rect 1290 1103 1293 1116
rect 1298 1113 1301 1126
rect 1306 1103 1309 1266
rect 1266 1013 1285 1016
rect 1258 933 1261 1006
rect 1266 916 1269 966
rect 1262 913 1269 916
rect 1262 836 1265 913
rect 1274 846 1277 1006
rect 1290 996 1293 1096
rect 1286 993 1293 996
rect 1286 936 1289 993
rect 1286 933 1293 936
rect 1290 916 1293 933
rect 1298 923 1301 1006
rect 1306 923 1309 996
rect 1314 976 1317 2203
rect 1322 1953 1325 2223
rect 1330 2213 1333 2226
rect 1346 2213 1349 2406
rect 1354 2393 1357 2433
rect 1362 2246 1365 2596
rect 1370 2413 1373 2426
rect 1378 2406 1381 2586
rect 1402 2546 1405 2653
rect 1466 2613 1469 2626
rect 1402 2543 1413 2546
rect 1394 2523 1405 2526
rect 1410 2516 1413 2543
rect 1402 2513 1413 2516
rect 1402 2496 1405 2513
rect 1418 2506 1421 2576
rect 1450 2543 1469 2546
rect 1394 2493 1405 2496
rect 1410 2503 1421 2506
rect 1394 2436 1397 2493
rect 1394 2433 1401 2436
rect 1370 2403 1381 2406
rect 1386 2403 1389 2416
rect 1370 2386 1373 2403
rect 1370 2383 1381 2386
rect 1358 2243 1365 2246
rect 1330 1973 1333 2126
rect 1338 2013 1341 2136
rect 1346 2133 1349 2176
rect 1358 2166 1361 2243
rect 1378 2236 1381 2383
rect 1398 2356 1401 2433
rect 1410 2376 1413 2503
rect 1418 2403 1421 2426
rect 1426 2413 1429 2526
rect 1450 2476 1453 2543
rect 1458 2526 1461 2536
rect 1466 2533 1469 2543
rect 1474 2526 1477 2616
rect 1482 2533 1485 2606
rect 1458 2523 1477 2526
rect 1482 2506 1485 2526
rect 1474 2503 1485 2506
rect 1450 2473 1461 2476
rect 1434 2413 1437 2436
rect 1426 2376 1429 2406
rect 1442 2403 1445 2416
rect 1410 2373 1429 2376
rect 1410 2356 1413 2373
rect 1398 2353 1405 2356
rect 1410 2353 1417 2356
rect 1394 2323 1397 2336
rect 1402 2306 1405 2353
rect 1370 2233 1381 2236
rect 1394 2303 1405 2306
rect 1394 2236 1397 2303
rect 1414 2296 1417 2353
rect 1426 2316 1429 2366
rect 1450 2333 1453 2416
rect 1458 2406 1461 2473
rect 1474 2436 1477 2503
rect 1474 2433 1485 2436
rect 1458 2403 1469 2406
rect 1426 2313 1437 2316
rect 1410 2293 1417 2296
rect 1394 2233 1401 2236
rect 1358 2163 1365 2166
rect 1362 2143 1365 2163
rect 1354 2133 1365 2136
rect 1354 2113 1357 2126
rect 1370 2036 1373 2233
rect 1378 2123 1381 2146
rect 1386 2113 1389 2216
rect 1398 2186 1401 2233
rect 1410 2193 1413 2293
rect 1434 2236 1437 2313
rect 1434 2233 1445 2236
rect 1426 2203 1429 2226
rect 1398 2183 1405 2186
rect 1362 2005 1365 2036
rect 1370 2033 1389 2036
rect 1378 1986 1381 2026
rect 1338 1933 1341 1956
rect 1354 1933 1357 1976
rect 1354 1913 1357 1926
rect 1322 1733 1325 1806
rect 1330 1803 1333 1826
rect 1354 1813 1357 1836
rect 1330 1666 1333 1766
rect 1346 1713 1349 1726
rect 1362 1723 1365 1986
rect 1370 1983 1381 1986
rect 1370 1686 1373 1983
rect 1386 1976 1389 2033
rect 1402 2023 1405 2183
rect 1434 2156 1437 2206
rect 1418 2153 1437 2156
rect 1418 2106 1421 2153
rect 1418 2103 1429 2106
rect 1426 2026 1429 2103
rect 1442 2033 1445 2233
rect 1458 2216 1461 2326
rect 1474 2323 1477 2416
rect 1458 2213 1477 2216
rect 1450 2166 1453 2206
rect 1466 2173 1469 2206
rect 1482 2186 1485 2433
rect 1490 2376 1493 2913
rect 1506 2886 1509 2906
rect 1502 2883 1509 2886
rect 1502 2766 1505 2883
rect 1502 2763 1509 2766
rect 1498 2533 1501 2746
rect 1506 2723 1509 2763
rect 1514 2756 1517 2986
rect 1522 2906 1525 3013
rect 1538 2996 1541 3016
rect 1534 2993 1541 2996
rect 1534 2926 1537 2993
rect 1546 2983 1549 3093
rect 1594 3046 1597 3173
rect 1602 3123 1605 3166
rect 1594 3043 1601 3046
rect 1554 2973 1557 3006
rect 1570 3005 1573 3016
rect 1598 2996 1601 3043
rect 1594 2993 1601 2996
rect 1534 2923 1541 2926
rect 1546 2923 1549 2936
rect 1554 2933 1557 2946
rect 1522 2903 1529 2906
rect 1526 2846 1529 2903
rect 1522 2843 1529 2846
rect 1522 2776 1525 2843
rect 1538 2783 1541 2923
rect 1554 2843 1557 2926
rect 1522 2773 1533 2776
rect 1562 2766 1565 2926
rect 1570 2813 1573 2936
rect 1578 2923 1581 2976
rect 1594 2943 1597 2993
rect 1610 2926 1613 3206
rect 1626 3143 1629 3206
rect 1642 3203 1645 3406
rect 1650 3403 1657 3406
rect 1654 3346 1657 3403
rect 1666 3393 1669 3406
rect 1654 3343 1661 3346
rect 1650 3303 1653 3326
rect 1626 3103 1629 3136
rect 1650 3076 1653 3286
rect 1658 3193 1661 3343
rect 1666 3216 1669 3386
rect 1674 3376 1677 3416
rect 1686 3406 1689 3513
rect 1686 3403 1693 3406
rect 1690 3383 1693 3403
rect 1674 3373 1685 3376
rect 1698 3373 1701 3606
rect 1706 3593 1709 3683
rect 1738 3616 1741 3636
rect 1730 3613 1741 3616
rect 1730 3556 1733 3613
rect 1730 3553 1741 3556
rect 1706 3383 1709 3406
rect 1674 3283 1677 3336
rect 1682 3323 1685 3373
rect 1690 3223 1693 3336
rect 1706 3333 1709 3346
rect 1714 3326 1717 3536
rect 1730 3413 1733 3526
rect 1698 3323 1717 3326
rect 1666 3213 1693 3216
rect 1682 3193 1685 3206
rect 1690 3143 1693 3213
rect 1674 3123 1677 3136
rect 1698 3133 1701 3206
rect 1706 3203 1709 3306
rect 1722 3233 1725 3406
rect 1642 3073 1653 3076
rect 1618 2983 1621 3016
rect 1642 2966 1645 3073
rect 1642 2963 1653 2966
rect 1618 2933 1621 2946
rect 1602 2923 1613 2926
rect 1602 2866 1605 2923
rect 1602 2863 1613 2866
rect 1578 2836 1581 2856
rect 1578 2833 1585 2836
rect 1554 2763 1565 2766
rect 1514 2753 1525 2756
rect 1498 2393 1501 2526
rect 1506 2523 1509 2716
rect 1522 2586 1525 2753
rect 1546 2603 1549 2616
rect 1514 2583 1525 2586
rect 1514 2503 1517 2583
rect 1490 2373 1497 2376
rect 1494 2276 1497 2373
rect 1514 2366 1517 2406
rect 1514 2363 1525 2366
rect 1522 2356 1525 2363
rect 1522 2353 1533 2356
rect 1522 2333 1525 2353
rect 1546 2296 1549 2526
rect 1554 2523 1557 2763
rect 1570 2646 1573 2806
rect 1582 2736 1585 2833
rect 1610 2803 1613 2863
rect 1626 2813 1629 2926
rect 1634 2923 1637 2936
rect 1642 2933 1645 2946
rect 1650 2906 1653 2963
rect 1642 2903 1653 2906
rect 1642 2806 1645 2903
rect 1642 2803 1653 2806
rect 1610 2756 1613 2796
rect 1578 2733 1585 2736
rect 1602 2753 1613 2756
rect 1578 2713 1581 2733
rect 1602 2706 1605 2753
rect 1602 2703 1613 2706
rect 1566 2643 1573 2646
rect 1566 2596 1569 2643
rect 1566 2593 1573 2596
rect 1570 2573 1573 2593
rect 1562 2506 1565 2536
rect 1578 2533 1581 2546
rect 1558 2503 1565 2506
rect 1558 2436 1561 2503
rect 1570 2456 1573 2526
rect 1586 2523 1589 2536
rect 1570 2453 1581 2456
rect 1558 2433 1565 2436
rect 1562 2413 1565 2433
rect 1578 2423 1581 2453
rect 1538 2293 1549 2296
rect 1494 2273 1501 2276
rect 1478 2183 1485 2186
rect 1450 2163 1469 2166
rect 1466 2123 1469 2163
rect 1478 2086 1481 2183
rect 1498 2176 1501 2273
rect 1538 2226 1541 2293
rect 1538 2223 1549 2226
rect 1490 2173 1501 2176
rect 1490 2093 1493 2173
rect 1522 2123 1525 2206
rect 1530 2143 1533 2206
rect 1478 2083 1485 2086
rect 1426 2023 1445 2026
rect 1378 1743 1381 1976
rect 1386 1973 1393 1976
rect 1390 1896 1393 1973
rect 1402 1916 1405 2006
rect 1426 1933 1429 2016
rect 1434 1923 1437 1996
rect 1442 1973 1445 2023
rect 1458 1956 1461 1976
rect 1458 1953 1465 1956
rect 1402 1913 1413 1916
rect 1390 1893 1397 1896
rect 1394 1826 1397 1893
rect 1386 1823 1397 1826
rect 1386 1763 1389 1823
rect 1410 1806 1413 1913
rect 1442 1846 1445 1936
rect 1450 1913 1453 1926
rect 1462 1906 1465 1953
rect 1394 1803 1413 1806
rect 1434 1843 1445 1846
rect 1458 1903 1465 1906
rect 1394 1733 1397 1803
rect 1434 1796 1437 1843
rect 1450 1796 1453 1826
rect 1458 1813 1461 1903
rect 1482 1873 1485 2083
rect 1506 1856 1509 2086
rect 1546 2073 1549 2223
rect 1562 2193 1565 2406
rect 1578 2356 1581 2396
rect 1574 2353 1581 2356
rect 1574 2266 1577 2353
rect 1594 2333 1597 2656
rect 1610 2636 1613 2703
rect 1634 2653 1637 2786
rect 1650 2743 1653 2803
rect 1610 2633 1617 2636
rect 1634 2633 1637 2646
rect 1602 2533 1605 2586
rect 1614 2566 1617 2633
rect 1626 2613 1629 2626
rect 1642 2616 1645 2676
rect 1638 2613 1645 2616
rect 1610 2563 1617 2566
rect 1610 2543 1613 2563
rect 1638 2546 1641 2613
rect 1638 2543 1645 2546
rect 1634 2506 1637 2526
rect 1626 2503 1637 2506
rect 1610 2413 1613 2426
rect 1626 2366 1629 2503
rect 1642 2373 1645 2543
rect 1650 2383 1653 2626
rect 1658 2366 1661 3086
rect 1666 3003 1669 3016
rect 1666 2906 1669 2996
rect 1674 2963 1677 3096
rect 1714 3093 1717 3206
rect 1682 2923 1685 3006
rect 1698 3005 1701 3016
rect 1722 2993 1725 3136
rect 1690 2933 1693 2986
rect 1730 2976 1733 3386
rect 1738 3106 1741 3553
rect 1746 3533 1749 3626
rect 1770 3596 1773 3693
rect 1786 3603 1789 3726
rect 1802 3723 1805 3936
rect 1810 3896 1813 4003
rect 1826 3953 1829 4006
rect 1818 3943 1837 3946
rect 1818 3933 1821 3943
rect 1818 3913 1821 3926
rect 1826 3923 1829 3936
rect 1834 3923 1837 3943
rect 1810 3893 1817 3896
rect 1814 3716 1817 3893
rect 1842 3766 1845 3926
rect 1850 3923 1853 3936
rect 1842 3763 1853 3766
rect 1826 3743 1845 3746
rect 1826 3733 1829 3743
rect 1810 3713 1817 3716
rect 1826 3713 1829 3726
rect 1834 3723 1837 3736
rect 1842 3723 1845 3743
rect 1850 3723 1853 3763
rect 1858 3736 1861 3936
rect 1874 3913 1877 4043
rect 1898 3936 1901 4136
rect 1906 4093 1909 4126
rect 1914 4076 1917 4153
rect 1922 4116 1925 4226
rect 1930 4213 1933 4246
rect 1938 4203 1941 4256
rect 1946 4196 1949 4216
rect 1954 4203 1957 4216
rect 1970 4213 1973 4526
rect 1978 4513 1981 4526
rect 1994 4523 1997 4583
rect 2010 4513 2013 4526
rect 1986 4363 1989 4406
rect 1986 4343 2005 4346
rect 1986 4333 1989 4343
rect 1994 4303 1997 4336
rect 2002 4323 2005 4343
rect 2010 4253 2013 4436
rect 2018 4413 2021 4616
rect 2026 4503 2029 4526
rect 2034 4513 2037 4536
rect 2058 4523 2061 4616
rect 2098 4573 2101 4606
rect 2138 4583 2141 4606
rect 2034 4413 2037 4496
rect 2066 4493 2069 4526
rect 2098 4516 2101 4536
rect 2106 4533 2109 4566
rect 2122 4543 2141 4546
rect 2094 4513 2101 4516
rect 2082 4413 2085 4506
rect 2094 4466 2097 4513
rect 2106 4476 2109 4526
rect 2122 4523 2125 4543
rect 2130 4523 2133 4536
rect 2138 4533 2141 4543
rect 2146 4513 2149 4526
rect 2162 4523 2165 4616
rect 2210 4546 2213 4566
rect 2202 4543 2213 4546
rect 2106 4473 2117 4476
rect 2094 4463 2101 4466
rect 2098 4413 2101 4463
rect 2090 4373 2093 4406
rect 2018 4233 2021 4326
rect 1962 4196 1965 4206
rect 1930 4133 1933 4186
rect 1922 4113 1929 4116
rect 1910 4073 1917 4076
rect 1910 3956 1913 4073
rect 1926 4066 1929 4113
rect 1938 4076 1941 4196
rect 1946 4193 1965 4196
rect 1994 4123 1997 4216
rect 2026 4213 2029 4326
rect 2042 4246 2045 4366
rect 2106 4353 2109 4406
rect 2114 4336 2117 4473
rect 2170 4446 2173 4526
rect 2202 4466 2205 4543
rect 2202 4463 2213 4466
rect 2170 4443 2181 4446
rect 2146 4366 2149 4406
rect 2178 4396 2181 4443
rect 2194 4413 2197 4426
rect 2170 4393 2181 4396
rect 2106 4333 2117 4336
rect 2138 4363 2149 4366
rect 2138 4333 2141 4363
rect 2154 4333 2157 4376
rect 2170 4336 2173 4393
rect 2162 4333 2173 4336
rect 2042 4243 2049 4246
rect 2010 4183 2013 4206
rect 2018 4133 2021 4176
rect 1938 4073 1949 4076
rect 1922 4063 1929 4066
rect 1910 3953 1917 3956
rect 1898 3933 1909 3936
rect 1874 3803 1877 3816
rect 1898 3813 1901 3926
rect 1858 3733 1869 3736
rect 1866 3716 1869 3733
rect 1858 3713 1869 3716
rect 1770 3593 1781 3596
rect 1746 3406 1749 3526
rect 1746 3403 1757 3406
rect 1746 3213 1749 3336
rect 1754 3313 1757 3403
rect 1762 3386 1765 3566
rect 1778 3526 1781 3593
rect 1774 3523 1781 3526
rect 1774 3456 1777 3523
rect 1774 3453 1781 3456
rect 1778 3433 1781 3453
rect 1778 3403 1781 3426
rect 1762 3383 1773 3386
rect 1770 3306 1773 3383
rect 1786 3333 1789 3516
rect 1794 3413 1797 3536
rect 1794 3316 1797 3406
rect 1802 3376 1805 3606
rect 1810 3393 1813 3713
rect 1858 3636 1861 3713
rect 1858 3633 1865 3636
rect 1818 3413 1821 3626
rect 1826 3613 1845 3616
rect 1842 3603 1845 3613
rect 1842 3583 1845 3596
rect 1802 3373 1813 3376
rect 1762 3303 1773 3306
rect 1786 3313 1797 3316
rect 1746 3123 1749 3146
rect 1754 3123 1757 3206
rect 1762 3166 1765 3303
rect 1786 3246 1789 3313
rect 1810 3306 1813 3373
rect 1826 3323 1829 3526
rect 1842 3386 1845 3436
rect 1850 3423 1853 3626
rect 1862 3556 1865 3633
rect 1874 3583 1877 3796
rect 1906 3793 1909 3933
rect 1882 3733 1885 3776
rect 1914 3773 1917 3953
rect 1898 3743 1917 3746
rect 1882 3713 1885 3726
rect 1890 3706 1893 3736
rect 1898 3723 1901 3743
rect 1906 3723 1909 3736
rect 1914 3733 1917 3743
rect 1922 3723 1925 4063
rect 1946 4026 1949 4073
rect 1938 4023 1949 4026
rect 1938 4003 1941 4023
rect 1938 3943 1957 3946
rect 1930 3923 1933 3936
rect 1938 3933 1941 3943
rect 1946 3876 1949 3936
rect 1954 3923 1957 3943
rect 1962 3923 1965 3946
rect 1994 3923 1997 4046
rect 1946 3873 1957 3876
rect 1954 3763 1957 3873
rect 1962 3736 1965 3796
rect 1978 3793 1981 3816
rect 2002 3813 2005 3926
rect 2018 3826 2021 4126
rect 2034 4123 2037 4236
rect 2046 4196 2049 4243
rect 2058 4203 2061 4326
rect 2106 4286 2109 4333
rect 2098 4283 2109 4286
rect 2042 4193 2049 4196
rect 2066 4196 2069 4216
rect 2074 4203 2077 4256
rect 2082 4213 2085 4226
rect 2082 4196 2085 4206
rect 2066 4193 2085 4196
rect 2042 4173 2045 4193
rect 2082 4156 2085 4176
rect 2058 4113 2061 4156
rect 2082 4153 2089 4156
rect 2086 4096 2089 4153
rect 2082 4093 2089 4096
rect 2082 4076 2085 4093
rect 2074 4073 2085 4076
rect 2074 3966 2077 4073
rect 2098 4056 2101 4283
rect 2114 4213 2117 4326
rect 2162 4213 2165 4333
rect 2170 4223 2173 4326
rect 2178 4233 2181 4336
rect 2186 4253 2189 4326
rect 2202 4313 2205 4326
rect 2146 4133 2149 4206
rect 2170 4143 2173 4206
rect 2178 4203 2181 4216
rect 2194 4213 2197 4246
rect 2202 4213 2205 4226
rect 2210 4193 2213 4463
rect 2218 4333 2221 4616
rect 2230 4576 2233 4623
rect 2250 4613 2253 4626
rect 2226 4573 2233 4576
rect 2242 4576 2245 4606
rect 2242 4573 2253 4576
rect 2226 4433 2229 4573
rect 2234 4523 2237 4556
rect 2226 4203 2229 4416
rect 2234 4413 2237 4426
rect 2242 4396 2245 4546
rect 2250 4523 2253 4573
rect 2258 4543 2261 4616
rect 2290 4613 2293 4626
rect 2306 4596 2309 4643
rect 2386 4613 2389 4626
rect 2394 4613 2405 4616
rect 2426 4613 2429 4626
rect 2306 4593 2317 4596
rect 2274 4533 2277 4566
rect 2238 4393 2245 4396
rect 2238 4316 2241 4393
rect 2250 4323 2253 4406
rect 2238 4313 2245 4316
rect 2242 4266 2245 4313
rect 2258 4276 2261 4436
rect 2266 4323 2269 4526
rect 2282 4383 2285 4406
rect 2274 4333 2277 4356
rect 2282 4306 2285 4326
rect 2282 4303 2289 4306
rect 2258 4273 2277 4276
rect 2242 4263 2269 4266
rect 2090 4053 2101 4056
rect 2090 4006 2093 4053
rect 2106 4013 2109 4126
rect 2146 4036 2149 4126
rect 2154 4123 2157 4136
rect 2130 4033 2149 4036
rect 2090 4003 2101 4006
rect 2074 3963 2085 3966
rect 2034 3943 2053 3946
rect 2026 3923 2029 3936
rect 2034 3913 2037 3943
rect 2042 3923 2045 3936
rect 2050 3933 2053 3943
rect 2074 3933 2077 3946
rect 2058 3923 2069 3926
rect 2082 3916 2085 3963
rect 2098 3923 2101 4003
rect 2106 3923 2109 3936
rect 2058 3896 2061 3916
rect 2050 3893 2061 3896
rect 2074 3913 2085 3916
rect 2050 3836 2053 3893
rect 2074 3866 2077 3913
rect 2130 3876 2133 4033
rect 2154 4006 2157 4026
rect 2146 4003 2157 4006
rect 2146 3926 2149 4003
rect 2162 3933 2165 4016
rect 2170 3996 2173 4136
rect 2194 4123 2197 4136
rect 2194 3996 2197 4006
rect 2202 4003 2205 4106
rect 2210 3996 2213 4016
rect 2234 4013 2237 4246
rect 2242 4163 2245 4216
rect 2250 4156 2253 4206
rect 2242 4153 2253 4156
rect 2170 3993 2177 3996
rect 2194 3993 2213 3996
rect 2174 3926 2177 3993
rect 2146 3923 2157 3926
rect 2130 3873 2149 3876
rect 2066 3863 2077 3866
rect 2050 3833 2061 3836
rect 2018 3823 2025 3826
rect 1954 3733 1965 3736
rect 1890 3703 1901 3706
rect 1898 3636 1901 3703
rect 1954 3666 1957 3733
rect 1954 3663 1965 3666
rect 1890 3633 1901 3636
rect 1882 3613 1885 3626
rect 1890 3613 1893 3633
rect 1962 3613 1965 3663
rect 1970 3613 1973 3726
rect 1994 3633 1997 3736
rect 2010 3726 2013 3816
rect 2022 3766 2025 3823
rect 2058 3773 2061 3833
rect 2018 3763 2025 3766
rect 2018 3743 2021 3763
rect 2010 3723 2021 3726
rect 2018 3626 2021 3723
rect 2050 3696 2053 3716
rect 2042 3693 2053 3696
rect 2042 3646 2045 3693
rect 2042 3643 2053 3646
rect 2010 3623 2021 3626
rect 1994 3603 1997 3616
rect 1858 3553 1865 3556
rect 1858 3533 1861 3553
rect 1858 3393 1861 3416
rect 1842 3383 1861 3386
rect 1842 3306 1845 3336
rect 1802 3303 1813 3306
rect 1834 3303 1845 3306
rect 1786 3243 1797 3246
rect 1778 3213 1781 3226
rect 1762 3163 1773 3166
rect 1770 3116 1773 3163
rect 1786 3126 1789 3216
rect 1794 3183 1797 3243
rect 1794 3133 1797 3166
rect 1802 3133 1805 3303
rect 1834 3246 1837 3303
rect 1834 3243 1845 3246
rect 1826 3203 1829 3216
rect 1786 3123 1797 3126
rect 1762 3113 1773 3116
rect 1738 3103 1745 3106
rect 1742 3036 1745 3103
rect 1762 3056 1765 3113
rect 1762 3053 1769 3056
rect 1706 2973 1733 2976
rect 1738 3033 1745 3036
rect 1666 2903 1677 2906
rect 1674 2786 1677 2903
rect 1698 2836 1701 2926
rect 1690 2833 1701 2836
rect 1706 2833 1709 2973
rect 1714 2863 1717 2966
rect 1722 2926 1725 2946
rect 1722 2923 1729 2926
rect 1726 2846 1729 2923
rect 1722 2843 1729 2846
rect 1690 2813 1693 2833
rect 1698 2823 1701 2833
rect 1706 2813 1717 2816
rect 1670 2783 1677 2786
rect 1670 2706 1673 2783
rect 1698 2766 1701 2806
rect 1722 2793 1725 2843
rect 1730 2813 1733 2826
rect 1738 2776 1741 3033
rect 1746 2933 1749 3016
rect 1766 2956 1769 3053
rect 1766 2953 1773 2956
rect 1762 2933 1765 2946
rect 1770 2936 1773 2953
rect 1778 2943 1781 3016
rect 1794 2993 1797 3123
rect 1802 3093 1805 3126
rect 1810 3066 1813 3136
rect 1826 3133 1829 3196
rect 1818 3103 1821 3126
rect 1842 3103 1845 3243
rect 1850 3213 1853 3336
rect 1858 3196 1861 3383
rect 1854 3193 1861 3196
rect 1854 3096 1857 3193
rect 1866 3106 1869 3456
rect 1874 3323 1877 3536
rect 1930 3533 1933 3596
rect 2010 3593 2013 3623
rect 2018 3563 2021 3606
rect 2042 3593 2045 3626
rect 1898 3513 1901 3526
rect 1906 3513 1909 3526
rect 1946 3486 1949 3536
rect 2018 3533 2021 3556
rect 2050 3553 2053 3643
rect 1970 3513 1973 3526
rect 1978 3513 1981 3526
rect 1946 3483 1957 3486
rect 1914 3413 1917 3426
rect 1954 3413 1957 3483
rect 2026 3433 2029 3536
rect 2050 3513 2053 3526
rect 2058 3513 2061 3526
rect 2002 3413 2021 3416
rect 1938 3346 1941 3406
rect 1954 3393 1957 3406
rect 1922 3343 1941 3346
rect 1882 3306 1885 3326
rect 1882 3303 1893 3306
rect 1890 3236 1893 3303
rect 1922 3266 1925 3343
rect 2002 3336 2005 3406
rect 2018 3346 2021 3406
rect 2026 3403 2029 3426
rect 2042 3406 2045 3446
rect 2034 3403 2045 3406
rect 2050 3396 2053 3436
rect 2034 3393 2053 3396
rect 2018 3343 2025 3346
rect 1922 3263 1933 3266
rect 1886 3233 1893 3236
rect 1886 3156 1889 3233
rect 1882 3153 1889 3156
rect 1874 3133 1877 3146
rect 1882 3123 1885 3153
rect 1898 3136 1901 3216
rect 1930 3193 1933 3263
rect 1890 3133 1901 3136
rect 1906 3153 1925 3156
rect 1906 3133 1909 3153
rect 1914 3133 1917 3146
rect 1866 3103 1877 3106
rect 1854 3093 1861 3096
rect 1810 3063 1821 3066
rect 1818 3013 1821 3063
rect 1858 3056 1861 3093
rect 1858 3053 1865 3056
rect 1862 2966 1865 3053
rect 1858 2963 1865 2966
rect 1770 2933 1781 2936
rect 1842 2933 1845 2946
rect 1858 2943 1861 2963
rect 1874 2946 1877 3103
rect 1898 3013 1901 3106
rect 1906 3093 1909 3126
rect 1922 3083 1925 3153
rect 1946 3123 1949 3326
rect 1962 3243 1965 3336
rect 1978 3256 1981 3336
rect 2002 3333 2013 3336
rect 1986 3313 1989 3326
rect 2002 3313 2005 3326
rect 2010 3296 2013 3333
rect 2002 3293 2013 3296
rect 1978 3253 1989 3256
rect 1986 3213 1989 3253
rect 1962 3193 1965 3206
rect 2002 3166 2005 3293
rect 2022 3276 2025 3343
rect 2018 3273 2025 3276
rect 2018 3253 2021 3273
rect 2002 3163 2013 3166
rect 1970 3116 1973 3136
rect 1962 3113 1973 3116
rect 1962 3036 1965 3113
rect 1962 3033 1973 3036
rect 1970 3013 1973 3033
rect 1930 2993 1933 3006
rect 1870 2943 1877 2946
rect 1746 2923 1773 2926
rect 1778 2916 1781 2933
rect 1762 2913 1781 2916
rect 1682 2763 1701 2766
rect 1730 2773 1741 2776
rect 1682 2723 1685 2763
rect 1666 2703 1673 2706
rect 1666 2496 1669 2703
rect 1730 2696 1733 2773
rect 1730 2693 1741 2696
rect 1674 2666 1677 2686
rect 1738 2673 1741 2693
rect 1674 2663 1685 2666
rect 1682 2586 1685 2663
rect 1714 2613 1717 2626
rect 1674 2583 1685 2586
rect 1674 2523 1677 2583
rect 1682 2513 1685 2536
rect 1690 2523 1693 2566
rect 1698 2533 1701 2556
rect 1666 2493 1677 2496
rect 1722 2493 1725 2626
rect 1746 2603 1749 2806
rect 1754 2793 1757 2806
rect 1762 2776 1765 2913
rect 1870 2896 1873 2943
rect 1978 2936 1981 3136
rect 1986 3133 1997 3136
rect 2010 3133 2013 3163
rect 2002 3103 2005 3126
rect 2018 3086 2021 3166
rect 2010 3083 2021 3086
rect 2010 2976 2013 3083
rect 2026 3066 2029 3216
rect 2034 3196 2037 3393
rect 2042 3213 2045 3336
rect 2050 3323 2053 3376
rect 2058 3323 2061 3406
rect 2050 3213 2053 3226
rect 2058 3196 2061 3256
rect 2034 3193 2045 3196
rect 2042 3126 2045 3193
rect 2022 3063 2029 3066
rect 2034 3123 2045 3126
rect 2054 3193 2061 3196
rect 2022 3006 2025 3063
rect 2034 3013 2037 3123
rect 2054 3106 2057 3193
rect 2050 3103 2057 3106
rect 2050 3006 2053 3103
rect 2022 3003 2029 3006
rect 2050 3003 2061 3006
rect 2010 2973 2021 2976
rect 1866 2893 1873 2896
rect 1758 2773 1765 2776
rect 1758 2726 1761 2773
rect 1770 2733 1773 2816
rect 1758 2723 1765 2726
rect 1762 2633 1765 2723
rect 1802 2716 1805 2736
rect 1794 2713 1805 2716
rect 1810 2716 1813 2766
rect 1826 2733 1829 2816
rect 1866 2813 1869 2893
rect 1874 2813 1877 2826
rect 1850 2753 1853 2806
rect 1866 2746 1869 2806
rect 1882 2803 1885 2926
rect 1890 2776 1893 2816
rect 1850 2743 1869 2746
rect 1874 2773 1893 2776
rect 1850 2733 1853 2743
rect 1858 2733 1869 2736
rect 1842 2723 1861 2726
rect 1810 2713 1821 2716
rect 1858 2713 1861 2723
rect 1794 2646 1797 2713
rect 1794 2643 1805 2646
rect 1770 2613 1773 2636
rect 1786 2613 1789 2626
rect 1794 2563 1797 2606
rect 1802 2536 1805 2643
rect 1738 2523 1741 2534
rect 1802 2533 1809 2536
rect 1762 2513 1765 2526
rect 1674 2406 1677 2493
rect 1738 2426 1741 2486
rect 1738 2423 1745 2426
rect 1666 2403 1677 2406
rect 1666 2383 1669 2403
rect 1626 2363 1637 2366
rect 1658 2363 1665 2366
rect 1574 2263 1581 2266
rect 1570 2213 1573 2246
rect 1578 2213 1581 2263
rect 1586 2203 1589 2306
rect 1618 2303 1621 2326
rect 1594 2213 1597 2226
rect 1610 2213 1613 2226
rect 1618 2193 1621 2206
rect 1594 2123 1597 2136
rect 1562 2033 1565 2096
rect 1626 2076 1629 2126
rect 1634 2113 1637 2363
rect 1662 2286 1665 2363
rect 1658 2283 1665 2286
rect 1658 2216 1661 2283
rect 1658 2213 1665 2216
rect 1642 2096 1645 2146
rect 1618 2073 1629 2076
rect 1638 2093 1645 2096
rect 1522 1993 1525 2016
rect 1530 1973 1533 2026
rect 1570 2013 1573 2046
rect 1514 1906 1517 1926
rect 1514 1903 1525 1906
rect 1498 1853 1509 1856
rect 1466 1833 1477 1836
rect 1474 1803 1477 1826
rect 1434 1793 1445 1796
rect 1450 1793 1461 1796
rect 1394 1696 1397 1726
rect 1394 1693 1405 1696
rect 1370 1683 1389 1686
rect 1322 1663 1333 1666
rect 1322 1603 1325 1663
rect 1330 1623 1357 1626
rect 1322 1403 1325 1526
rect 1330 1513 1333 1623
rect 1354 1616 1357 1623
rect 1338 1566 1341 1606
rect 1346 1603 1349 1616
rect 1354 1613 1365 1616
rect 1370 1613 1381 1616
rect 1354 1593 1357 1606
rect 1370 1583 1373 1606
rect 1338 1563 1357 1566
rect 1322 1206 1325 1396
rect 1330 1223 1333 1506
rect 1354 1456 1357 1563
rect 1378 1516 1381 1536
rect 1342 1453 1357 1456
rect 1370 1513 1381 1516
rect 1370 1456 1373 1513
rect 1370 1453 1381 1456
rect 1342 1336 1345 1453
rect 1362 1413 1365 1436
rect 1338 1333 1345 1336
rect 1338 1233 1341 1333
rect 1322 1203 1329 1206
rect 1326 1136 1329 1203
rect 1338 1183 1341 1216
rect 1346 1203 1349 1316
rect 1354 1306 1357 1406
rect 1370 1333 1373 1416
rect 1378 1396 1381 1453
rect 1386 1413 1389 1683
rect 1402 1556 1405 1693
rect 1426 1686 1429 1776
rect 1442 1753 1445 1793
rect 1458 1696 1461 1793
rect 1498 1786 1501 1853
rect 1522 1846 1525 1903
rect 1538 1866 1541 1936
rect 1546 1873 1549 1926
rect 1554 1923 1557 1936
rect 1562 1913 1565 1966
rect 1538 1863 1557 1866
rect 1514 1843 1525 1846
rect 1498 1783 1509 1786
rect 1506 1763 1509 1783
rect 1474 1723 1477 1736
rect 1514 1723 1517 1843
rect 1554 1813 1557 1863
rect 1594 1856 1597 2026
rect 1618 2003 1621 2073
rect 1638 2006 1641 2093
rect 1634 2003 1641 2006
rect 1594 1853 1605 1856
rect 1530 1793 1533 1806
rect 1602 1776 1605 1853
rect 1594 1773 1605 1776
rect 1522 1706 1525 1766
rect 1394 1553 1405 1556
rect 1418 1683 1429 1686
rect 1450 1693 1461 1696
rect 1514 1703 1525 1706
rect 1394 1533 1397 1553
rect 1418 1526 1421 1683
rect 1450 1616 1453 1693
rect 1514 1636 1517 1703
rect 1514 1633 1525 1636
rect 1434 1593 1437 1616
rect 1450 1613 1457 1616
rect 1394 1403 1397 1516
rect 1410 1433 1413 1526
rect 1418 1523 1429 1526
rect 1442 1523 1445 1606
rect 1454 1556 1457 1613
rect 1450 1553 1457 1556
rect 1426 1466 1429 1523
rect 1418 1463 1429 1466
rect 1378 1393 1385 1396
rect 1382 1326 1385 1393
rect 1378 1323 1385 1326
rect 1354 1303 1365 1306
rect 1362 1236 1365 1303
rect 1378 1236 1381 1323
rect 1354 1233 1365 1236
rect 1374 1233 1381 1236
rect 1354 1213 1357 1233
rect 1362 1203 1365 1216
rect 1374 1186 1377 1233
rect 1374 1183 1381 1186
rect 1378 1146 1381 1183
rect 1394 1173 1397 1326
rect 1402 1303 1405 1416
rect 1418 1403 1421 1463
rect 1450 1393 1453 1553
rect 1482 1543 1485 1606
rect 1498 1603 1501 1616
rect 1458 1503 1461 1536
rect 1474 1456 1477 1536
rect 1506 1533 1509 1606
rect 1522 1586 1525 1633
rect 1530 1603 1533 1756
rect 1594 1746 1597 1773
rect 1594 1743 1605 1746
rect 1554 1733 1565 1736
rect 1546 1713 1549 1726
rect 1554 1596 1557 1726
rect 1562 1613 1565 1726
rect 1570 1703 1573 1726
rect 1578 1706 1581 1736
rect 1586 1713 1589 1736
rect 1578 1703 1589 1706
rect 1554 1593 1565 1596
rect 1578 1593 1581 1606
rect 1522 1583 1533 1586
rect 1466 1453 1477 1456
rect 1466 1413 1469 1453
rect 1418 1313 1421 1326
rect 1466 1323 1469 1356
rect 1482 1323 1485 1526
rect 1490 1296 1493 1506
rect 1506 1426 1509 1526
rect 1530 1446 1533 1583
rect 1554 1533 1557 1546
rect 1562 1523 1565 1593
rect 1522 1443 1533 1446
rect 1506 1423 1513 1426
rect 1498 1333 1501 1416
rect 1510 1326 1513 1423
rect 1482 1293 1493 1296
rect 1506 1323 1513 1326
rect 1442 1193 1445 1216
rect 1378 1143 1389 1146
rect 1322 1133 1329 1136
rect 1322 1113 1325 1133
rect 1322 993 1325 1006
rect 1314 973 1321 976
rect 1318 916 1321 973
rect 1290 913 1301 916
rect 1298 856 1301 913
rect 1314 913 1321 916
rect 1298 853 1305 856
rect 1274 843 1281 846
rect 1262 833 1269 836
rect 1234 613 1237 626
rect 1202 583 1213 586
rect 1210 526 1213 583
rect 1242 553 1245 776
rect 1258 733 1261 816
rect 1266 773 1269 833
rect 1278 756 1281 843
rect 1302 776 1305 853
rect 1274 753 1281 756
rect 1298 773 1305 776
rect 1274 733 1277 753
rect 1266 723 1285 726
rect 1290 723 1293 736
rect 1298 726 1301 773
rect 1306 733 1309 746
rect 1298 723 1309 726
rect 1250 613 1253 686
rect 1258 613 1261 626
rect 1266 603 1269 723
rect 1298 633 1301 646
rect 1290 613 1293 626
rect 1306 623 1309 723
rect 1314 693 1317 913
rect 1322 743 1325 816
rect 1330 776 1333 1106
rect 1354 966 1357 1136
rect 1386 1096 1389 1143
rect 1402 1113 1405 1126
rect 1346 963 1357 966
rect 1378 1093 1389 1096
rect 1346 946 1349 963
rect 1378 953 1381 1093
rect 1434 1056 1437 1126
rect 1442 1123 1445 1186
rect 1482 1156 1485 1293
rect 1506 1196 1509 1323
rect 1522 1206 1525 1443
rect 1546 1403 1549 1416
rect 1570 1413 1573 1536
rect 1586 1533 1589 1703
rect 1602 1626 1605 1743
rect 1594 1623 1605 1626
rect 1578 1513 1581 1526
rect 1594 1506 1597 1623
rect 1602 1543 1605 1606
rect 1586 1503 1597 1506
rect 1586 1446 1589 1503
rect 1610 1456 1613 1526
rect 1618 1503 1621 1976
rect 1626 1703 1629 1726
rect 1634 1686 1637 2003
rect 1642 1903 1645 1926
rect 1650 1886 1653 2206
rect 1662 2106 1665 2213
rect 1674 2143 1677 2386
rect 1706 2363 1709 2406
rect 1698 2336 1701 2356
rect 1694 2333 1701 2336
rect 1682 2213 1685 2326
rect 1694 2256 1697 2333
rect 1694 2253 1701 2256
rect 1690 2213 1693 2236
rect 1698 2203 1701 2253
rect 1706 2223 1709 2356
rect 1730 2353 1733 2416
rect 1742 2346 1745 2423
rect 1738 2343 1745 2346
rect 1714 2303 1717 2316
rect 1706 2213 1725 2216
rect 1714 2193 1717 2206
rect 1722 2196 1725 2213
rect 1722 2193 1729 2196
rect 1682 2133 1693 2136
rect 1714 2133 1717 2176
rect 1658 2103 1665 2106
rect 1658 2083 1661 2103
rect 1658 1996 1661 2056
rect 1666 2013 1669 2036
rect 1698 2033 1701 2126
rect 1714 2113 1717 2126
rect 1726 2106 1729 2193
rect 1722 2103 1729 2106
rect 1722 2086 1725 2103
rect 1714 2083 1725 2086
rect 1682 2023 1701 2026
rect 1658 1993 1669 1996
rect 1682 1993 1685 2023
rect 1698 2016 1701 2023
rect 1666 1926 1669 1993
rect 1690 1926 1693 2016
rect 1698 2013 1709 2016
rect 1714 2003 1717 2083
rect 1738 2066 1741 2343
rect 1754 2236 1757 2496
rect 1806 2486 1809 2533
rect 1802 2483 1809 2486
rect 1770 2413 1789 2416
rect 1770 2366 1773 2413
rect 1766 2363 1773 2366
rect 1766 2256 1769 2363
rect 1766 2253 1773 2256
rect 1754 2233 1761 2236
rect 1730 2063 1741 2066
rect 1658 1923 1669 1926
rect 1682 1923 1693 1926
rect 1714 1923 1717 1996
rect 1730 1936 1733 2063
rect 1738 2013 1741 2026
rect 1746 2023 1749 2226
rect 1758 2166 1761 2233
rect 1770 2203 1773 2253
rect 1754 2163 1761 2166
rect 1746 1996 1749 2016
rect 1722 1933 1733 1936
rect 1742 1993 1749 1996
rect 1658 1903 1661 1923
rect 1682 1906 1685 1923
rect 1678 1903 1685 1906
rect 1630 1683 1637 1686
rect 1646 1883 1653 1886
rect 1610 1453 1621 1456
rect 1578 1443 1589 1446
rect 1530 1316 1533 1336
rect 1530 1313 1541 1316
rect 1538 1236 1541 1313
rect 1502 1193 1509 1196
rect 1514 1203 1525 1206
rect 1530 1233 1541 1236
rect 1482 1153 1493 1156
rect 1426 1053 1437 1056
rect 1418 1003 1421 1016
rect 1426 1003 1429 1053
rect 1442 1046 1445 1096
rect 1450 1083 1453 1136
rect 1490 1133 1493 1153
rect 1502 1126 1505 1193
rect 1498 1123 1505 1126
rect 1482 1096 1485 1116
rect 1474 1093 1485 1096
rect 1434 1043 1445 1046
rect 1346 943 1357 946
rect 1354 886 1357 943
rect 1370 923 1373 946
rect 1394 913 1397 936
rect 1410 923 1413 936
rect 1346 883 1357 886
rect 1346 803 1349 883
rect 1394 793 1397 816
rect 1330 773 1341 776
rect 1322 613 1325 716
rect 1338 616 1341 773
rect 1362 733 1365 756
rect 1410 713 1413 726
rect 1330 613 1341 616
rect 1386 613 1389 706
rect 1234 533 1245 536
rect 1258 533 1261 546
rect 1202 523 1213 526
rect 1234 523 1261 526
rect 1202 503 1205 523
rect 1274 443 1277 526
rect 1130 313 1133 336
rect 1138 333 1141 376
rect 1174 373 1181 376
rect 1138 303 1141 326
rect 1154 313 1157 326
rect 1162 266 1165 336
rect 1170 323 1173 356
rect 1154 263 1165 266
rect 1154 213 1157 263
rect 1178 213 1181 373
rect 1186 316 1189 406
rect 1194 333 1197 376
rect 1186 313 1197 316
rect 1178 193 1181 206
rect 1058 183 1069 186
rect 1074 183 1081 186
rect 1058 106 1061 183
rect 1074 153 1077 183
rect 1082 133 1085 166
rect 1130 123 1133 146
rect 1194 126 1197 313
rect 1210 303 1213 426
rect 1282 423 1285 526
rect 1226 323 1229 406
rect 1226 216 1229 236
rect 1218 213 1229 216
rect 1202 133 1205 186
rect 1218 166 1221 213
rect 1218 163 1229 166
rect 1218 133 1221 146
rect 1194 123 1213 126
rect 1226 123 1229 163
rect 1234 133 1237 216
rect 1242 213 1245 336
rect 1258 193 1261 406
rect 1282 366 1285 416
rect 1274 363 1285 366
rect 1274 316 1277 363
rect 1290 333 1293 376
rect 1298 333 1301 606
rect 1314 456 1317 556
rect 1322 513 1325 536
rect 1330 523 1333 613
rect 1338 523 1341 536
rect 1346 523 1349 596
rect 1370 593 1373 606
rect 1314 453 1333 456
rect 1306 393 1309 416
rect 1290 323 1309 326
rect 1274 313 1285 316
rect 1282 256 1285 313
rect 1314 266 1317 336
rect 1322 323 1325 356
rect 1306 263 1317 266
rect 1282 253 1293 256
rect 1290 176 1293 253
rect 1306 213 1309 263
rect 1330 213 1333 453
rect 1346 376 1349 506
rect 1354 413 1357 536
rect 1362 456 1365 526
rect 1370 503 1373 536
rect 1386 533 1389 546
rect 1378 513 1381 526
rect 1362 453 1373 456
rect 1370 413 1373 453
rect 1394 416 1397 526
rect 1410 493 1413 626
rect 1386 413 1397 416
rect 1402 413 1405 436
rect 1378 393 1381 406
rect 1338 373 1349 376
rect 1346 343 1349 373
rect 1330 193 1333 206
rect 1346 183 1349 206
rect 1282 173 1293 176
rect 1258 133 1261 166
rect 1282 146 1285 173
rect 1282 143 1293 146
rect 1058 103 1069 106
rect 1066 33 1069 103
rect 1290 96 1293 143
rect 1306 123 1309 136
rect 1354 126 1357 376
rect 1370 296 1373 366
rect 1386 353 1389 413
rect 1378 303 1381 326
rect 1386 306 1389 336
rect 1394 333 1397 406
rect 1402 333 1405 386
rect 1410 326 1413 406
rect 1418 363 1421 656
rect 1434 533 1437 1043
rect 1474 1036 1477 1093
rect 1474 1033 1485 1036
rect 1458 1013 1477 1016
rect 1442 973 1445 1006
rect 1450 923 1453 1006
rect 1482 1003 1485 1033
rect 1458 933 1461 946
rect 1466 886 1469 926
rect 1458 883 1469 886
rect 1458 826 1461 883
rect 1458 823 1469 826
rect 1458 786 1461 806
rect 1450 783 1461 786
rect 1450 736 1453 783
rect 1450 733 1461 736
rect 1450 696 1453 716
rect 1446 693 1453 696
rect 1446 626 1449 693
rect 1458 653 1461 733
rect 1466 703 1469 823
rect 1446 623 1453 626
rect 1474 623 1477 936
rect 1482 916 1485 996
rect 1490 936 1493 1026
rect 1498 943 1501 1123
rect 1506 1003 1509 1016
rect 1514 993 1517 1203
rect 1522 1133 1525 1196
rect 1530 1123 1533 1233
rect 1538 1133 1541 1216
rect 1554 1186 1557 1326
rect 1578 1323 1581 1443
rect 1586 1333 1589 1346
rect 1554 1183 1565 1186
rect 1546 1126 1549 1176
rect 1538 1123 1549 1126
rect 1538 1056 1541 1123
rect 1562 1116 1565 1183
rect 1530 1053 1541 1056
rect 1554 1113 1565 1116
rect 1530 1006 1533 1053
rect 1546 1013 1549 1046
rect 1530 1003 1541 1006
rect 1490 933 1501 936
rect 1482 913 1489 916
rect 1486 846 1489 913
rect 1482 843 1489 846
rect 1482 803 1485 843
rect 1490 813 1493 826
rect 1498 813 1501 933
rect 1514 913 1517 936
rect 1538 876 1541 1003
rect 1530 873 1541 876
rect 1530 826 1533 873
rect 1506 793 1509 806
rect 1514 733 1517 826
rect 1530 823 1541 826
rect 1538 783 1541 823
rect 1546 766 1549 956
rect 1554 906 1557 1113
rect 1562 1013 1565 1026
rect 1578 1013 1581 1316
rect 1594 1303 1597 1426
rect 1618 1376 1621 1453
rect 1610 1373 1621 1376
rect 1610 1286 1613 1373
rect 1630 1336 1633 1683
rect 1646 1676 1649 1883
rect 1658 1813 1661 1876
rect 1666 1813 1669 1896
rect 1678 1836 1681 1903
rect 1678 1833 1685 1836
rect 1642 1673 1649 1676
rect 1642 1603 1645 1673
rect 1650 1613 1653 1646
rect 1658 1603 1661 1716
rect 1626 1333 1633 1336
rect 1626 1316 1629 1333
rect 1602 1283 1613 1286
rect 1622 1313 1629 1316
rect 1602 1156 1605 1283
rect 1622 1236 1625 1313
rect 1622 1233 1629 1236
rect 1602 1153 1613 1156
rect 1594 1116 1597 1136
rect 1590 1113 1597 1116
rect 1590 1036 1593 1113
rect 1590 1033 1597 1036
rect 1602 1033 1605 1126
rect 1594 1013 1597 1033
rect 1562 1003 1573 1006
rect 1562 923 1565 946
rect 1594 916 1597 936
rect 1586 913 1597 916
rect 1554 903 1561 906
rect 1558 846 1561 903
rect 1538 763 1549 766
rect 1554 843 1561 846
rect 1450 603 1453 623
rect 1458 613 1477 616
rect 1482 573 1485 726
rect 1490 603 1493 726
rect 1498 673 1501 726
rect 1538 636 1541 763
rect 1538 633 1549 636
rect 1514 613 1517 626
rect 1434 413 1437 526
rect 1458 523 1461 546
rect 1498 536 1501 556
rect 1498 533 1505 536
rect 1502 486 1505 533
rect 1514 523 1517 606
rect 1522 513 1525 616
rect 1530 593 1533 616
rect 1498 483 1505 486
rect 1442 373 1445 406
rect 1498 366 1501 483
rect 1546 453 1549 633
rect 1554 613 1557 843
rect 1570 803 1573 886
rect 1586 866 1589 913
rect 1602 896 1605 1026
rect 1610 933 1613 1153
rect 1618 1133 1621 1216
rect 1626 1116 1629 1233
rect 1634 1203 1637 1326
rect 1622 1113 1629 1116
rect 1622 1036 1625 1113
rect 1634 1043 1637 1166
rect 1642 1093 1645 1566
rect 1650 1486 1653 1556
rect 1666 1533 1669 1616
rect 1674 1613 1677 1816
rect 1682 1783 1685 1833
rect 1690 1766 1693 1916
rect 1698 1896 1701 1916
rect 1722 1903 1725 1933
rect 1730 1903 1733 1916
rect 1698 1893 1709 1896
rect 1706 1826 1709 1893
rect 1686 1763 1693 1766
rect 1698 1823 1709 1826
rect 1686 1636 1689 1763
rect 1698 1646 1701 1823
rect 1730 1813 1733 1896
rect 1742 1876 1745 1993
rect 1754 1893 1757 2163
rect 1770 2153 1773 2196
rect 1778 2146 1781 2406
rect 1786 2203 1789 2396
rect 1794 2253 1797 2426
rect 1802 2336 1805 2483
rect 1818 2436 1821 2713
rect 1842 2613 1845 2626
rect 1850 2603 1853 2636
rect 1858 2603 1861 2706
rect 1874 2683 1877 2773
rect 1882 2733 1885 2766
rect 1898 2756 1901 2806
rect 1906 2796 1909 2826
rect 1922 2803 1925 2926
rect 1954 2923 1957 2934
rect 1978 2933 1989 2936
rect 1978 2866 1981 2926
rect 1986 2876 1989 2933
rect 2018 2876 2021 2973
rect 1986 2873 1997 2876
rect 1962 2863 1981 2866
rect 1906 2793 1913 2796
rect 1930 2793 1933 2806
rect 1954 2796 1957 2826
rect 1962 2803 1965 2863
rect 1946 2793 1957 2796
rect 1894 2753 1901 2756
rect 1866 2613 1877 2616
rect 1882 2613 1885 2726
rect 1894 2686 1897 2753
rect 1910 2746 1913 2793
rect 1906 2743 1913 2746
rect 1946 2746 1949 2793
rect 1946 2743 1957 2746
rect 1906 2696 1909 2743
rect 1922 2713 1925 2736
rect 1906 2693 1913 2696
rect 1894 2683 1901 2686
rect 1898 2646 1901 2683
rect 1894 2643 1901 2646
rect 1874 2596 1877 2613
rect 1870 2593 1877 2596
rect 1842 2503 1845 2576
rect 1850 2573 1861 2576
rect 1810 2433 1821 2436
rect 1810 2353 1813 2433
rect 1802 2333 1813 2336
rect 1810 2246 1813 2333
rect 1802 2243 1813 2246
rect 1794 2213 1797 2236
rect 1802 2196 1805 2243
rect 1810 2203 1813 2226
rect 1802 2193 1813 2196
rect 1766 2143 1781 2146
rect 1766 2046 1769 2143
rect 1762 2043 1769 2046
rect 1742 1873 1749 1876
rect 1746 1853 1749 1873
rect 1754 1836 1757 1876
rect 1750 1833 1757 1836
rect 1706 1706 1709 1786
rect 1714 1723 1717 1806
rect 1738 1803 1741 1826
rect 1750 1776 1753 1833
rect 1750 1773 1757 1776
rect 1754 1733 1757 1773
rect 1722 1723 1741 1726
rect 1706 1703 1717 1706
rect 1698 1643 1705 1646
rect 1686 1633 1693 1636
rect 1674 1573 1677 1606
rect 1682 1603 1685 1616
rect 1690 1553 1693 1633
rect 1702 1566 1705 1643
rect 1698 1563 1705 1566
rect 1666 1523 1677 1526
rect 1666 1503 1669 1523
rect 1682 1486 1685 1536
rect 1650 1483 1661 1486
rect 1658 1376 1661 1483
rect 1674 1483 1685 1486
rect 1674 1436 1677 1483
rect 1674 1433 1685 1436
rect 1682 1413 1685 1433
rect 1690 1423 1693 1526
rect 1698 1503 1701 1563
rect 1714 1546 1717 1703
rect 1738 1603 1741 1723
rect 1754 1713 1757 1726
rect 1746 1613 1749 1636
rect 1754 1606 1757 1706
rect 1746 1603 1757 1606
rect 1706 1543 1717 1546
rect 1706 1506 1709 1543
rect 1730 1523 1741 1526
rect 1706 1503 1717 1506
rect 1714 1436 1717 1503
rect 1706 1433 1717 1436
rect 1650 1373 1661 1376
rect 1650 1276 1653 1373
rect 1650 1273 1661 1276
rect 1658 1196 1661 1273
rect 1650 1193 1661 1196
rect 1618 1033 1625 1036
rect 1642 1033 1645 1066
rect 1618 993 1621 1033
rect 1610 913 1613 926
rect 1618 923 1621 936
rect 1626 923 1629 1016
rect 1634 1013 1637 1026
rect 1650 1023 1653 1193
rect 1658 1126 1661 1136
rect 1666 1133 1669 1176
rect 1682 1133 1685 1326
rect 1690 1313 1693 1406
rect 1706 1403 1709 1433
rect 1730 1393 1733 1416
rect 1738 1413 1741 1523
rect 1746 1506 1749 1603
rect 1754 1523 1757 1596
rect 1762 1553 1765 2043
rect 1770 1983 1773 2026
rect 1778 1973 1781 2136
rect 1786 2123 1789 2156
rect 1794 2133 1805 2136
rect 1810 2133 1813 2193
rect 1802 2003 1805 2126
rect 1810 2013 1813 2046
rect 1818 2003 1821 2216
rect 1826 2186 1829 2416
rect 1842 2413 1845 2446
rect 1850 2433 1853 2573
rect 1858 2523 1861 2566
rect 1870 2456 1873 2593
rect 1870 2453 1877 2456
rect 1874 2433 1877 2453
rect 1850 2413 1853 2426
rect 1858 2403 1861 2426
rect 1850 2383 1861 2386
rect 1850 2326 1853 2383
rect 1882 2356 1885 2606
rect 1894 2596 1897 2643
rect 1910 2626 1913 2693
rect 1906 2623 1913 2626
rect 1906 2603 1909 2623
rect 1894 2593 1901 2596
rect 1914 2593 1917 2606
rect 1898 2383 1901 2593
rect 1922 2433 1925 2676
rect 1930 2423 1933 2446
rect 1938 2413 1941 2616
rect 1946 2606 1949 2726
rect 1954 2703 1957 2743
rect 1962 2713 1965 2776
rect 1970 2766 1973 2836
rect 1994 2826 1997 2873
rect 1978 2813 1981 2826
rect 1986 2823 1997 2826
rect 2010 2873 2021 2876
rect 1986 2806 1989 2823
rect 1978 2803 1989 2806
rect 1978 2783 1981 2803
rect 2010 2766 2013 2873
rect 1970 2763 1981 2766
rect 2010 2763 2021 2766
rect 1978 2716 1981 2763
rect 1970 2713 1981 2716
rect 1970 2693 1973 2713
rect 2002 2676 2005 2716
rect 1986 2673 2005 2676
rect 1962 2616 1965 2656
rect 1962 2613 1973 2616
rect 1946 2603 1957 2606
rect 1954 2523 1957 2603
rect 1970 2536 1973 2613
rect 1986 2546 1989 2673
rect 2010 2656 2013 2746
rect 2002 2653 2013 2656
rect 2002 2566 2005 2653
rect 2002 2563 2013 2566
rect 1986 2543 2005 2546
rect 1962 2533 1973 2536
rect 1954 2496 1957 2516
rect 1962 2503 1965 2533
rect 1950 2493 1957 2496
rect 1882 2353 1893 2356
rect 1842 2323 1853 2326
rect 1842 2236 1845 2323
rect 1866 2316 1869 2336
rect 1858 2246 1861 2316
rect 1866 2313 1877 2316
rect 1858 2243 1865 2246
rect 1842 2233 1853 2236
rect 1834 2203 1837 2216
rect 1842 2193 1845 2206
rect 1826 2183 1833 2186
rect 1830 2036 1833 2183
rect 1850 2136 1853 2233
rect 1862 2196 1865 2243
rect 1842 2133 1853 2136
rect 1858 2193 1865 2196
rect 1842 2043 1845 2133
rect 1850 2083 1853 2126
rect 1858 2076 1861 2193
rect 1874 2176 1877 2313
rect 1850 2073 1861 2076
rect 1866 2173 1877 2176
rect 1830 2033 1845 2036
rect 1834 2013 1837 2026
rect 1842 2006 1845 2033
rect 1826 2003 1845 2006
rect 1778 1866 1781 1956
rect 1802 1946 1805 1996
rect 1802 1943 1809 1946
rect 1806 1896 1809 1943
rect 1818 1913 1821 1926
rect 1802 1893 1809 1896
rect 1778 1863 1789 1866
rect 1746 1503 1753 1506
rect 1750 1426 1753 1503
rect 1746 1423 1753 1426
rect 1746 1376 1749 1423
rect 1730 1373 1749 1376
rect 1730 1356 1733 1373
rect 1754 1356 1757 1406
rect 1730 1353 1741 1356
rect 1714 1276 1717 1336
rect 1710 1273 1717 1276
rect 1658 1123 1677 1126
rect 1666 1056 1669 1116
rect 1690 1106 1693 1126
rect 1682 1103 1693 1106
rect 1666 1053 1673 1056
rect 1658 1016 1661 1046
rect 1650 1013 1661 1016
rect 1634 933 1637 946
rect 1650 933 1653 1013
rect 1670 1006 1673 1053
rect 1682 1046 1685 1103
rect 1682 1043 1693 1046
rect 1698 1043 1701 1236
rect 1710 1186 1713 1273
rect 1706 1183 1713 1186
rect 1706 1126 1709 1183
rect 1706 1123 1713 1126
rect 1710 1066 1713 1123
rect 1722 1113 1725 1306
rect 1738 1246 1741 1353
rect 1730 1243 1741 1246
rect 1750 1353 1757 1356
rect 1750 1246 1753 1353
rect 1762 1303 1765 1536
rect 1770 1403 1773 1856
rect 1786 1776 1789 1863
rect 1778 1773 1789 1776
rect 1778 1743 1781 1773
rect 1778 1696 1781 1736
rect 1802 1733 1805 1893
rect 1810 1803 1813 1816
rect 1778 1693 1789 1696
rect 1778 1323 1781 1646
rect 1786 1533 1789 1693
rect 1794 1613 1797 1686
rect 1802 1603 1805 1716
rect 1818 1683 1821 1816
rect 1810 1576 1813 1616
rect 1818 1583 1821 1606
rect 1794 1573 1813 1576
rect 1794 1533 1797 1573
rect 1786 1506 1789 1526
rect 1802 1523 1805 1556
rect 1810 1506 1813 1536
rect 1786 1503 1797 1506
rect 1794 1426 1797 1503
rect 1790 1423 1797 1426
rect 1806 1503 1813 1506
rect 1806 1426 1809 1503
rect 1806 1423 1813 1426
rect 1790 1316 1793 1423
rect 1802 1333 1805 1406
rect 1786 1313 1793 1316
rect 1810 1313 1813 1423
rect 1750 1243 1757 1246
rect 1730 1213 1733 1243
rect 1746 1213 1749 1226
rect 1706 1063 1713 1066
rect 1690 1016 1693 1043
rect 1666 1003 1673 1006
rect 1682 1013 1693 1016
rect 1642 903 1645 926
rect 1658 913 1661 936
rect 1666 906 1669 1003
rect 1650 903 1669 906
rect 1602 893 1609 896
rect 1586 863 1597 866
rect 1562 723 1565 746
rect 1570 626 1573 796
rect 1594 793 1597 863
rect 1606 786 1609 893
rect 1618 803 1621 816
rect 1650 806 1653 903
rect 1658 813 1661 826
rect 1666 813 1669 856
rect 1682 853 1685 1013
rect 1706 1003 1709 1063
rect 1730 1026 1733 1206
rect 1738 1113 1741 1206
rect 1746 1053 1749 1186
rect 1754 1153 1757 1243
rect 1762 1163 1765 1256
rect 1762 1056 1765 1136
rect 1770 1126 1773 1206
rect 1778 1133 1781 1176
rect 1786 1136 1789 1313
rect 1810 1233 1813 1276
rect 1794 1146 1797 1226
rect 1802 1213 1805 1226
rect 1818 1213 1821 1576
rect 1826 1196 1829 2003
rect 1842 1886 1845 1986
rect 1850 1923 1853 2073
rect 1834 1883 1845 1886
rect 1834 1753 1837 1883
rect 1842 1813 1845 1866
rect 1850 1803 1853 1916
rect 1858 1873 1861 2046
rect 1866 1993 1869 2173
rect 1882 2123 1885 2136
rect 1874 2013 1877 2086
rect 1890 2083 1893 2353
rect 1906 2323 1909 2356
rect 1950 2346 1953 2493
rect 1950 2343 1957 2346
rect 1906 2146 1909 2316
rect 1938 2213 1941 2226
rect 1902 2143 1909 2146
rect 1930 2156 1933 2166
rect 1946 2156 1949 2326
rect 1954 2286 1957 2343
rect 1962 2303 1965 2466
rect 1970 2353 1973 2516
rect 1978 2403 1981 2416
rect 1986 2403 1989 2526
rect 2002 2516 2005 2543
rect 2010 2523 2013 2563
rect 2002 2513 2013 2516
rect 1994 2413 2005 2416
rect 1978 2323 1981 2386
rect 1954 2283 1961 2286
rect 1958 2166 1961 2283
rect 2002 2236 2005 2406
rect 2010 2313 2013 2513
rect 2018 2483 2021 2763
rect 2026 2673 2029 3003
rect 2058 2983 2061 3003
rect 2034 2906 2037 2926
rect 2034 2903 2045 2906
rect 2042 2826 2045 2903
rect 2034 2823 2045 2826
rect 2034 2803 2037 2823
rect 2058 2813 2061 2926
rect 2066 2923 2069 3863
rect 2082 3793 2085 3806
rect 2090 3733 2093 3776
rect 2122 3746 2125 3856
rect 2130 3813 2133 3826
rect 2122 3743 2129 3746
rect 2082 3713 2101 3716
rect 2082 3533 2085 3713
rect 2090 3516 2093 3536
rect 2082 3513 2093 3516
rect 2082 3446 2085 3513
rect 2082 3443 2093 3446
rect 2074 3123 2077 3416
rect 2082 3276 2085 3426
rect 2090 3373 2093 3443
rect 2098 3383 2101 3656
rect 2106 3613 2109 3726
rect 2114 3613 2117 3736
rect 2126 3646 2129 3743
rect 2146 3733 2149 3873
rect 2138 3673 2141 3726
rect 2154 3716 2157 3923
rect 2170 3923 2177 3926
rect 2170 3853 2173 3923
rect 2162 3796 2165 3836
rect 2170 3813 2173 3826
rect 2162 3793 2169 3796
rect 2150 3713 2157 3716
rect 2122 3643 2129 3646
rect 2082 3273 2093 3276
rect 2082 3203 2085 3266
rect 2090 3163 2093 3273
rect 2098 3203 2101 3326
rect 2106 3213 2109 3476
rect 2114 3213 2117 3536
rect 2122 3496 2125 3643
rect 2150 3626 2153 3713
rect 2166 3706 2169 3793
rect 2162 3703 2169 3706
rect 2130 3603 2133 3626
rect 2150 3623 2157 3626
rect 2162 3623 2165 3703
rect 2178 3646 2181 3736
rect 2186 3706 2189 3966
rect 2218 3943 2221 4006
rect 2242 3996 2245 4153
rect 2250 4123 2253 4146
rect 2258 4133 2261 4256
rect 2266 4203 2269 4263
rect 2234 3993 2245 3996
rect 2202 3813 2205 3936
rect 2210 3743 2213 3896
rect 2234 3856 2237 3993
rect 2250 3953 2253 4086
rect 2266 4003 2269 4116
rect 2274 4063 2277 4273
rect 2286 4246 2289 4303
rect 2282 4243 2289 4246
rect 2282 4083 2285 4243
rect 2298 4176 2301 4386
rect 2306 4323 2309 4416
rect 2314 4366 2317 4593
rect 2338 4583 2341 4606
rect 2378 4603 2397 4606
rect 2370 4403 2373 4526
rect 2394 4523 2397 4603
rect 2402 4466 2405 4613
rect 2410 4533 2413 4556
rect 2402 4463 2413 4466
rect 2386 4413 2389 4426
rect 2402 4413 2405 4436
rect 2314 4363 2321 4366
rect 2318 4316 2321 4363
rect 2314 4313 2321 4316
rect 2314 4246 2317 4313
rect 2330 4256 2333 4366
rect 2370 4326 2373 4336
rect 2378 4333 2381 4406
rect 2394 4363 2397 4406
rect 2402 4366 2405 4406
rect 2410 4403 2413 4463
rect 2426 4383 2429 4596
rect 2474 4593 2477 4606
rect 2490 4576 2493 4646
rect 2506 4593 2509 4606
rect 2490 4573 2501 4576
rect 2498 4546 2501 4573
rect 2490 4543 2501 4546
rect 2442 4513 2445 4526
rect 2450 4423 2453 4526
rect 2490 4466 2493 4543
rect 2490 4463 2497 4466
rect 2474 4413 2477 4426
rect 2494 4376 2497 4463
rect 2494 4373 2501 4376
rect 2402 4363 2413 4366
rect 2362 4316 2365 4326
rect 2370 4323 2389 4326
rect 2354 4313 2365 4316
rect 2330 4253 2337 4256
rect 2314 4243 2325 4246
rect 2290 4173 2301 4176
rect 2290 4023 2293 4173
rect 2298 4123 2301 4156
rect 2250 3916 2253 3946
rect 2250 3913 2261 3916
rect 2234 3853 2245 3856
rect 2218 3796 2221 3806
rect 2226 3803 2229 3836
rect 2234 3796 2237 3816
rect 2242 3813 2245 3853
rect 2218 3793 2237 3796
rect 2210 3726 2213 3736
rect 2194 3723 2213 3726
rect 2226 3706 2229 3786
rect 2186 3703 2197 3706
rect 2174 3643 2181 3646
rect 2138 3533 2141 3606
rect 2130 3513 2133 3526
rect 2138 3513 2141 3526
rect 2122 3493 2129 3496
rect 2126 3356 2129 3493
rect 2146 3423 2149 3606
rect 2154 3466 2157 3623
rect 2162 3533 2165 3616
rect 2174 3586 2177 3643
rect 2194 3636 2197 3703
rect 2218 3703 2229 3706
rect 2218 3646 2221 3703
rect 2218 3643 2229 3646
rect 2186 3633 2197 3636
rect 2186 3593 2189 3633
rect 2194 3613 2213 3616
rect 2218 3613 2221 3626
rect 2210 3603 2213 3613
rect 2226 3593 2229 3643
rect 2174 3583 2181 3586
rect 2170 3473 2173 3536
rect 2154 3463 2173 3466
rect 2122 3353 2129 3356
rect 2122 3276 2125 3353
rect 2146 3323 2149 3406
rect 2162 3313 2165 3326
rect 2170 3296 2173 3463
rect 2162 3293 2173 3296
rect 2122 3273 2133 3276
rect 2082 3123 2085 3136
rect 2098 3066 2101 3136
rect 2114 3133 2117 3206
rect 2130 3146 2133 3273
rect 2162 3226 2165 3293
rect 2162 3223 2173 3226
rect 2122 3143 2133 3146
rect 2106 3103 2109 3126
rect 2098 3063 2109 3066
rect 2106 3013 2109 3063
rect 2082 2993 2085 3006
rect 2074 2933 2077 2946
rect 2090 2933 2093 2956
rect 2098 2853 2101 2986
rect 2098 2813 2101 2826
rect 2042 2743 2045 2806
rect 2034 2703 2037 2726
rect 2042 2713 2045 2736
rect 2050 2733 2053 2796
rect 2082 2746 2085 2806
rect 2106 2796 2109 2946
rect 2102 2793 2109 2796
rect 2090 2753 2093 2766
rect 2082 2743 2093 2746
rect 2066 2733 2077 2736
rect 2058 2703 2061 2726
rect 2074 2693 2077 2726
rect 2082 2713 2085 2726
rect 2090 2706 2093 2743
rect 2082 2703 2093 2706
rect 2102 2706 2105 2793
rect 2114 2763 2117 3126
rect 2122 3013 2125 3143
rect 2130 3103 2133 3126
rect 2146 3056 2149 3216
rect 2170 3193 2173 3223
rect 2170 3116 2173 3136
rect 2162 3113 2173 3116
rect 2146 3053 2153 3056
rect 2150 2996 2153 3053
rect 2162 3036 2165 3113
rect 2162 3033 2173 3036
rect 2146 2993 2153 2996
rect 2146 2976 2149 2993
rect 2138 2973 2149 2976
rect 2122 2906 2125 2936
rect 2138 2906 2141 2973
rect 2162 2933 2165 3016
rect 2170 3013 2173 3033
rect 2178 2916 2181 3583
rect 2234 3533 2237 3716
rect 2186 3523 2197 3526
rect 2186 3506 2189 3523
rect 2202 3513 2205 3526
rect 2186 3503 2193 3506
rect 2190 3436 2193 3503
rect 2242 3476 2245 3796
rect 2250 3573 2253 3906
rect 2258 3803 2261 3913
rect 2266 3906 2269 3946
rect 2274 3933 2277 3976
rect 2290 3923 2293 4016
rect 2266 3903 2277 3906
rect 2274 3846 2277 3903
rect 2298 3853 2301 4066
rect 2306 3963 2309 4136
rect 2314 4123 2317 4166
rect 2322 4056 2325 4243
rect 2334 4206 2337 4253
rect 2346 4213 2349 4226
rect 2330 4203 2337 4206
rect 2330 4146 2333 4203
rect 2338 4166 2341 4186
rect 2338 4163 2349 4166
rect 2330 4143 2337 4146
rect 2334 4066 2337 4143
rect 2314 4053 2325 4056
rect 2330 4063 2337 4066
rect 2314 4043 2317 4053
rect 2330 3946 2333 4063
rect 2346 4046 2349 4163
rect 2362 4123 2365 4313
rect 2394 4256 2397 4356
rect 2402 4333 2405 4363
rect 2418 4296 2421 4326
rect 2418 4293 2425 4296
rect 2386 4253 2397 4256
rect 2378 4196 2381 4216
rect 2370 4193 2381 4196
rect 2370 4133 2373 4193
rect 2386 4133 2389 4253
rect 2394 4133 2397 4246
rect 2402 4213 2405 4226
rect 2402 4126 2405 4206
rect 2378 4123 2405 4126
rect 2410 4106 2413 4286
rect 2422 4166 2425 4293
rect 2434 4183 2437 4346
rect 2458 4213 2461 4326
rect 2338 4043 2349 4046
rect 2402 4103 2413 4106
rect 2418 4163 2425 4166
rect 2338 4013 2341 4043
rect 2402 4036 2405 4103
rect 2402 4033 2413 4036
rect 2326 3943 2333 3946
rect 2346 3943 2349 4016
rect 2306 3923 2309 3936
rect 2270 3843 2277 3846
rect 2270 3796 2273 3843
rect 2314 3813 2317 3926
rect 2326 3806 2329 3943
rect 2354 3936 2357 4026
rect 2394 3973 2397 4016
rect 2410 4013 2413 4033
rect 2338 3873 2341 3936
rect 2346 3933 2357 3936
rect 2346 3913 2349 3933
rect 2354 3923 2365 3926
rect 2266 3793 2273 3796
rect 2290 3793 2293 3806
rect 2326 3803 2333 3806
rect 2266 3733 2269 3793
rect 2330 3783 2333 3803
rect 2338 3743 2341 3866
rect 2258 3706 2261 3726
rect 2274 3716 2277 3736
rect 2274 3713 2285 3716
rect 2314 3713 2317 3726
rect 2258 3703 2265 3706
rect 2262 3636 2265 3703
rect 2282 3636 2285 3713
rect 2258 3633 2265 3636
rect 2274 3633 2285 3636
rect 2258 3583 2261 3633
rect 2274 3536 2277 3633
rect 2322 3616 2325 3736
rect 2330 3713 2333 3736
rect 2258 3533 2277 3536
rect 2250 3513 2253 3526
rect 2242 3473 2249 3476
rect 2186 3433 2193 3436
rect 2186 3123 2189 3433
rect 2194 3393 2197 3416
rect 2194 3316 2197 3386
rect 2202 3333 2205 3346
rect 2194 3313 2201 3316
rect 2198 3246 2201 3313
rect 2194 3243 2201 3246
rect 2194 3193 2197 3243
rect 2194 3123 2197 3136
rect 2202 3116 2205 3186
rect 2194 3113 2205 3116
rect 2210 3116 2213 3406
rect 2234 3383 2237 3466
rect 2246 3406 2249 3473
rect 2242 3403 2249 3406
rect 2242 3353 2245 3403
rect 2218 3266 2221 3336
rect 2226 3323 2245 3326
rect 2250 3306 2253 3386
rect 2246 3303 2253 3306
rect 2218 3263 2237 3266
rect 2234 3213 2237 3263
rect 2218 3133 2221 3146
rect 2210 3113 2217 3116
rect 2194 3096 2197 3113
rect 2190 3093 2197 3096
rect 2190 2946 2193 3093
rect 2190 2943 2197 2946
rect 2170 2913 2181 2916
rect 2122 2903 2129 2906
rect 2138 2903 2149 2906
rect 2126 2846 2129 2903
rect 2146 2846 2149 2903
rect 2122 2843 2129 2846
rect 2138 2843 2149 2846
rect 2122 2793 2125 2843
rect 2138 2826 2141 2843
rect 2170 2836 2173 2913
rect 2170 2833 2181 2836
rect 2130 2823 2141 2826
rect 2130 2806 2133 2823
rect 2138 2813 2165 2816
rect 2130 2803 2149 2806
rect 2102 2703 2109 2706
rect 2026 2533 2029 2616
rect 2042 2613 2045 2686
rect 2058 2616 2061 2686
rect 2054 2613 2061 2616
rect 2034 2603 2045 2606
rect 2054 2556 2057 2613
rect 2066 2563 2069 2606
rect 2054 2553 2061 2556
rect 2002 2233 2009 2236
rect 1986 2203 1989 2226
rect 2006 2186 2009 2233
rect 2002 2183 2009 2186
rect 1958 2163 1973 2166
rect 1930 2153 1957 2156
rect 1902 2096 1905 2143
rect 1930 2096 1933 2153
rect 1954 2133 1957 2153
rect 1970 2143 1973 2163
rect 2002 2146 2005 2183
rect 1986 2143 2005 2146
rect 1902 2093 1909 2096
rect 1930 2093 1937 2096
rect 1906 2046 1909 2093
rect 1906 2043 1917 2046
rect 1866 1966 1869 1986
rect 1866 1963 1873 1966
rect 1870 1876 1873 1963
rect 1866 1873 1873 1876
rect 1858 1813 1861 1826
rect 1842 1733 1845 1766
rect 1834 1613 1837 1646
rect 1842 1603 1845 1726
rect 1822 1193 1829 1196
rect 1794 1143 1813 1146
rect 1786 1133 1797 1136
rect 1770 1123 1789 1126
rect 1794 1116 1797 1133
rect 1754 1053 1765 1056
rect 1730 1023 1741 1026
rect 1690 923 1693 936
rect 1706 906 1709 996
rect 1698 903 1709 906
rect 1698 836 1701 903
rect 1698 833 1709 836
rect 1682 813 1701 816
rect 1650 803 1661 806
rect 1666 803 1677 806
rect 1602 783 1609 786
rect 1658 786 1661 803
rect 1658 783 1669 786
rect 1690 783 1693 806
rect 1578 713 1581 726
rect 1570 623 1581 626
rect 1586 623 1589 736
rect 1602 716 1605 783
rect 1598 713 1605 716
rect 1598 656 1601 713
rect 1594 653 1601 656
rect 1578 603 1581 623
rect 1594 616 1597 653
rect 1586 613 1597 616
rect 1602 613 1605 636
rect 1570 513 1573 526
rect 1562 416 1565 446
rect 1530 413 1565 416
rect 1394 323 1413 326
rect 1386 303 1397 306
rect 1370 293 1381 296
rect 1362 133 1365 206
rect 1370 203 1373 236
rect 1378 203 1381 293
rect 1394 256 1397 303
rect 1386 253 1397 256
rect 1386 233 1389 253
rect 1418 213 1421 336
rect 1434 333 1437 366
rect 1498 363 1505 366
rect 1482 323 1485 356
rect 1502 286 1505 363
rect 1498 283 1505 286
rect 1450 213 1453 236
rect 1498 173 1501 283
rect 1514 193 1517 346
rect 1522 323 1525 406
rect 1570 403 1573 426
rect 1578 413 1581 596
rect 1586 523 1589 613
rect 1594 576 1597 606
rect 1594 573 1605 576
rect 1586 406 1589 456
rect 1594 413 1597 566
rect 1602 523 1605 573
rect 1610 523 1613 716
rect 1626 696 1629 756
rect 1634 723 1637 736
rect 1650 713 1653 726
rect 1658 703 1661 776
rect 1666 706 1669 783
rect 1674 723 1677 736
rect 1706 713 1709 833
rect 1714 733 1717 976
rect 1722 743 1725 966
rect 1730 883 1733 1016
rect 1738 973 1741 1023
rect 1746 1006 1749 1046
rect 1754 1013 1757 1053
rect 1746 1003 1757 1006
rect 1738 903 1741 926
rect 1730 803 1733 826
rect 1666 703 1677 706
rect 1626 693 1637 696
rect 1634 626 1637 693
rect 1658 646 1661 696
rect 1626 623 1637 626
rect 1650 643 1661 646
rect 1618 443 1621 606
rect 1626 516 1629 623
rect 1650 596 1653 643
rect 1674 636 1677 703
rect 1666 633 1677 636
rect 1666 603 1669 633
rect 1650 593 1661 596
rect 1642 533 1645 546
rect 1626 513 1637 516
rect 1634 446 1637 513
rect 1626 443 1637 446
rect 1578 403 1589 406
rect 1538 333 1541 346
rect 1522 183 1525 206
rect 1418 133 1421 166
rect 1354 123 1373 126
rect 1466 123 1469 166
rect 1538 123 1541 326
rect 1562 296 1565 336
rect 1554 293 1565 296
rect 1546 163 1549 206
rect 1554 203 1557 293
rect 1554 133 1557 196
rect 1570 183 1573 396
rect 1578 316 1581 403
rect 1586 323 1589 346
rect 1578 313 1589 316
rect 1586 183 1589 313
rect 1602 213 1605 406
rect 1610 323 1613 436
rect 1626 416 1629 443
rect 1650 433 1653 536
rect 1658 523 1661 593
rect 1690 553 1693 616
rect 1698 613 1701 706
rect 1698 586 1701 606
rect 1714 603 1717 716
rect 1722 706 1725 736
rect 1730 723 1733 796
rect 1738 733 1741 816
rect 1746 803 1749 986
rect 1746 733 1749 746
rect 1754 716 1757 1003
rect 1762 823 1765 936
rect 1770 926 1773 1116
rect 1786 1113 1797 1116
rect 1778 983 1781 1056
rect 1786 933 1789 1113
rect 1770 923 1789 926
rect 1746 713 1757 716
rect 1722 703 1733 706
rect 1730 636 1733 703
rect 1722 633 1733 636
rect 1722 616 1725 633
rect 1722 613 1741 616
rect 1698 583 1709 586
rect 1666 496 1669 536
rect 1674 513 1677 526
rect 1682 523 1685 546
rect 1706 516 1709 583
rect 1730 573 1733 606
rect 1746 533 1749 713
rect 1762 673 1765 806
rect 1754 603 1757 656
rect 1762 533 1765 616
rect 1770 593 1773 826
rect 1778 683 1781 846
rect 1778 586 1781 676
rect 1770 583 1781 586
rect 1770 516 1773 583
rect 1786 563 1789 916
rect 1794 906 1797 1026
rect 1802 1013 1805 1136
rect 1802 923 1805 996
rect 1794 903 1801 906
rect 1798 836 1801 903
rect 1810 843 1813 1143
rect 1822 1126 1825 1193
rect 1822 1123 1829 1126
rect 1818 963 1821 1106
rect 1826 1006 1829 1123
rect 1834 1043 1837 1596
rect 1842 1333 1845 1526
rect 1842 1313 1845 1326
rect 1842 1103 1845 1306
rect 1850 1096 1853 1686
rect 1858 1183 1861 1696
rect 1866 1506 1869 1873
rect 1874 1733 1877 1856
rect 1874 1713 1877 1726
rect 1882 1683 1885 1976
rect 1890 1953 1893 2006
rect 1914 1983 1917 2043
rect 1922 1976 1925 2086
rect 1934 2036 1937 2093
rect 1954 2056 1957 2126
rect 1954 2053 1961 2056
rect 1930 2033 1937 2036
rect 1930 2013 1933 2033
rect 1938 2003 1941 2016
rect 1958 1996 1961 2053
rect 1986 2046 1989 2143
rect 2002 2123 2005 2136
rect 2018 2126 2021 2426
rect 2042 2366 2045 2406
rect 2050 2383 2053 2446
rect 2058 2433 2061 2553
rect 2082 2443 2085 2703
rect 2106 2683 2109 2703
rect 2106 2603 2109 2616
rect 2114 2566 2117 2756
rect 2130 2723 2133 2736
rect 2122 2666 2125 2686
rect 2154 2683 2157 2806
rect 2178 2803 2181 2833
rect 2186 2803 2189 2926
rect 2122 2663 2129 2666
rect 2106 2563 2117 2566
rect 2106 2446 2109 2563
rect 2126 2556 2129 2663
rect 2146 2613 2165 2616
rect 2146 2576 2149 2613
rect 2122 2553 2129 2556
rect 2138 2573 2149 2576
rect 2122 2506 2125 2553
rect 2138 2533 2141 2573
rect 2146 2523 2149 2536
rect 2162 2533 2165 2606
rect 2178 2603 2181 2796
rect 2194 2756 2197 2943
rect 2202 2916 2205 3106
rect 2214 3046 2217 3113
rect 2210 3043 2217 3046
rect 2210 2933 2213 3043
rect 2226 3013 2229 3196
rect 2246 3186 2249 3303
rect 2246 3183 2253 3186
rect 2258 3183 2261 3533
rect 2266 3496 2269 3516
rect 2274 3513 2277 3526
rect 2266 3493 2273 3496
rect 2270 3426 2273 3493
rect 2266 3423 2273 3426
rect 2266 3253 2269 3423
rect 2234 3076 2237 3136
rect 2242 3123 2245 3136
rect 2250 3133 2253 3183
rect 2234 3073 2253 3076
rect 2258 3073 2261 3126
rect 2274 3103 2277 3406
rect 2282 3323 2285 3526
rect 2290 3513 2293 3616
rect 2306 3603 2309 3616
rect 2322 3613 2329 3616
rect 2306 3533 2309 3566
rect 2290 3413 2293 3426
rect 2306 3416 2309 3436
rect 2298 3413 2309 3416
rect 2314 3413 2317 3606
rect 2326 3546 2329 3613
rect 2338 3556 2341 3626
rect 2346 3563 2349 3716
rect 2354 3623 2357 3846
rect 2354 3603 2357 3616
rect 2338 3553 2349 3556
rect 2322 3543 2329 3546
rect 2306 3393 2309 3406
rect 2282 3096 2285 3236
rect 2290 3213 2293 3336
rect 2298 3296 2301 3356
rect 2306 3313 2309 3326
rect 2298 3293 2305 3296
rect 2302 3226 2305 3293
rect 2298 3223 2305 3226
rect 2274 3093 2285 3096
rect 2250 3013 2253 3073
rect 2266 3036 2269 3056
rect 2262 3033 2269 3036
rect 2226 2993 2229 3006
rect 2202 2913 2209 2916
rect 2206 2836 2209 2913
rect 2202 2833 2209 2836
rect 2202 2796 2205 2833
rect 2210 2803 2213 2816
rect 2218 2813 2221 2936
rect 2250 2903 2253 3006
rect 2262 2956 2265 3033
rect 2262 2953 2269 2956
rect 2258 2876 2261 2936
rect 2242 2873 2261 2876
rect 2242 2813 2245 2873
rect 2266 2823 2269 2953
rect 2274 2916 2277 3093
rect 2290 2983 2293 3186
rect 2298 2976 2301 3223
rect 2306 3026 2309 3206
rect 2314 3033 2317 3366
rect 2322 3176 2325 3543
rect 2330 3513 2333 3526
rect 2346 3496 2349 3553
rect 2342 3493 2349 3496
rect 2330 3323 2333 3436
rect 2342 3426 2345 3493
rect 2342 3423 2349 3426
rect 2338 3383 2341 3406
rect 2346 3366 2349 3423
rect 2342 3363 2349 3366
rect 2342 3316 2345 3363
rect 2354 3353 2357 3526
rect 2362 3516 2365 3856
rect 2370 3613 2373 3876
rect 2378 3796 2381 3956
rect 2394 3923 2397 3936
rect 2402 3923 2405 4006
rect 2418 3933 2421 4163
rect 2434 4036 2437 4136
rect 2430 4033 2437 4036
rect 2430 3986 2433 4033
rect 2442 4003 2445 4026
rect 2458 4013 2461 4126
rect 2466 4063 2469 4216
rect 2474 4046 2477 4166
rect 2470 4043 2477 4046
rect 2430 3983 2437 3986
rect 2434 3963 2437 3983
rect 2434 3943 2453 3946
rect 2410 3913 2413 3926
rect 2426 3906 2429 3936
rect 2434 3923 2437 3943
rect 2442 3923 2445 3936
rect 2450 3933 2453 3943
rect 2418 3903 2429 3906
rect 2386 3813 2405 3816
rect 2402 3806 2405 3813
rect 2378 3793 2385 3796
rect 2382 3716 2385 3793
rect 2394 3733 2397 3806
rect 2402 3803 2413 3806
rect 2402 3733 2405 3786
rect 2410 3733 2413 3803
rect 2418 3783 2421 3903
rect 2426 3876 2429 3896
rect 2458 3876 2461 4006
rect 2470 3976 2473 4043
rect 2470 3973 2477 3976
rect 2466 3923 2469 3956
rect 2426 3873 2437 3876
rect 2434 3816 2437 3873
rect 2450 3873 2461 3876
rect 2450 3856 2453 3873
rect 2474 3863 2477 3973
rect 2482 3903 2485 4336
rect 2498 4213 2501 4373
rect 2506 4336 2509 4536
rect 2522 4493 2525 4526
rect 2530 4476 2533 4536
rect 2526 4473 2533 4476
rect 2526 4426 2529 4473
rect 2538 4433 2541 4526
rect 2546 4523 2549 4606
rect 2554 4523 2557 4616
rect 2586 4603 2589 4616
rect 2658 4613 2661 4626
rect 2610 4593 2613 4606
rect 2578 4543 2597 4546
rect 2578 4533 2581 4543
rect 2578 4513 2581 4526
rect 2586 4523 2589 4536
rect 2594 4523 2597 4543
rect 2514 4413 2517 4426
rect 2526 4423 2533 4426
rect 2506 4333 2525 4336
rect 2530 4333 2533 4423
rect 2522 4303 2525 4326
rect 2530 4293 2533 4326
rect 2546 4323 2549 4406
rect 2554 4333 2557 4356
rect 2562 4283 2565 4446
rect 2610 4443 2613 4566
rect 2618 4523 2621 4536
rect 2634 4533 2637 4546
rect 2658 4536 2661 4596
rect 2690 4576 2693 4616
rect 2698 4613 2701 4626
rect 2682 4573 2693 4576
rect 2626 4463 2629 4526
rect 2650 4456 2653 4536
rect 2658 4533 2669 4536
rect 2682 4533 2685 4573
rect 2698 4556 2701 4606
rect 2690 4553 2701 4556
rect 2658 4473 2661 4526
rect 2630 4453 2653 4456
rect 2594 4343 2597 4406
rect 2602 4333 2613 4336
rect 2618 4323 2621 4416
rect 2630 4316 2633 4453
rect 2666 4426 2669 4533
rect 2674 4513 2677 4526
rect 2690 4523 2693 4553
rect 2714 4543 2717 4616
rect 2802 4613 2805 4626
rect 2842 4613 2845 4626
rect 2698 4523 2701 4536
rect 2706 4516 2709 4536
rect 2698 4513 2709 4516
rect 2662 4423 2669 4426
rect 2626 4313 2633 4316
rect 2522 4203 2525 4226
rect 2514 4056 2517 4126
rect 2522 4123 2525 4136
rect 2538 4113 2541 4206
rect 2546 4083 2549 4126
rect 2554 4066 2557 4146
rect 2562 4106 2565 4276
rect 2570 4123 2573 4216
rect 2602 4166 2605 4286
rect 2594 4163 2605 4166
rect 2562 4103 2569 4106
rect 2506 4053 2517 4056
rect 2550 4063 2557 4066
rect 2498 3936 2501 4016
rect 2506 4003 2509 4053
rect 2514 4013 2517 4026
rect 2530 4013 2533 4026
rect 2522 3993 2525 4006
rect 2538 4003 2541 4016
rect 2550 3996 2553 4063
rect 2566 4056 2569 4103
rect 2562 4053 2569 4056
rect 2550 3993 2557 3996
rect 2498 3933 2505 3936
rect 2426 3813 2437 3816
rect 2446 3853 2453 3856
rect 2426 3793 2429 3813
rect 2446 3776 2449 3853
rect 2490 3813 2493 3926
rect 2502 3876 2505 3933
rect 2498 3873 2505 3876
rect 2498 3853 2501 3873
rect 2446 3773 2453 3776
rect 2382 3713 2389 3716
rect 2378 3603 2381 3646
rect 2378 3533 2381 3556
rect 2362 3513 2373 3516
rect 2370 3446 2373 3513
rect 2386 3473 2389 3713
rect 2394 3523 2397 3606
rect 2362 3443 2373 3446
rect 2362 3376 2365 3443
rect 2402 3426 2405 3626
rect 2410 3553 2413 3716
rect 2418 3713 2421 3726
rect 2426 3646 2429 3746
rect 2450 3733 2453 3773
rect 2498 3746 2501 3796
rect 2474 3733 2477 3746
rect 2498 3743 2505 3746
rect 2514 3743 2517 3966
rect 2522 3913 2525 3976
rect 2554 3973 2557 3993
rect 2530 3793 2533 3946
rect 2562 3943 2565 4053
rect 2570 4003 2573 4016
rect 2578 4013 2581 4136
rect 2594 4056 2597 4163
rect 2610 4146 2613 4256
rect 2606 4143 2613 4146
rect 2606 4076 2609 4143
rect 2606 4073 2613 4076
rect 2594 4053 2605 4056
rect 2586 3976 2589 4006
rect 2582 3973 2589 3976
rect 2546 3923 2549 3936
rect 2538 3803 2541 3826
rect 2434 3663 2437 3726
rect 2502 3696 2505 3743
rect 2498 3693 2505 3696
rect 2426 3643 2437 3646
rect 2418 3593 2421 3626
rect 2434 3566 2437 3643
rect 2458 3603 2461 3616
rect 2466 3613 2485 3616
rect 2490 3613 2493 3626
rect 2426 3563 2437 3566
rect 2402 3423 2413 3426
rect 2378 3393 2381 3406
rect 2362 3373 2369 3376
rect 2354 3323 2357 3336
rect 2366 3316 2369 3373
rect 2378 3333 2381 3376
rect 2386 3323 2389 3356
rect 2394 3333 2397 3386
rect 2402 3373 2405 3416
rect 2342 3313 2349 3316
rect 2330 3196 2333 3286
rect 2338 3216 2341 3256
rect 2346 3226 2349 3313
rect 2362 3313 2369 3316
rect 2346 3223 2357 3226
rect 2338 3213 2357 3216
rect 2330 3193 2341 3196
rect 2322 3173 2329 3176
rect 2326 3106 2329 3173
rect 2322 3103 2329 3106
rect 2306 3023 2317 3026
rect 2282 2973 2301 2976
rect 2282 2923 2285 2973
rect 2290 2933 2301 2936
rect 2306 2933 2309 3016
rect 2274 2913 2293 2916
rect 2250 2813 2261 2816
rect 2266 2813 2277 2816
rect 2202 2793 2213 2796
rect 2194 2753 2201 2756
rect 2198 2706 2201 2753
rect 2194 2703 2201 2706
rect 2194 2653 2197 2703
rect 2202 2603 2205 2616
rect 2122 2503 2133 2506
rect 2106 2443 2117 2446
rect 2058 2403 2061 2426
rect 2066 2413 2077 2416
rect 2098 2403 2101 2426
rect 2042 2363 2049 2366
rect 2026 2293 2029 2326
rect 2046 2296 2049 2363
rect 2074 2356 2077 2376
rect 2070 2353 2077 2356
rect 2042 2293 2049 2296
rect 2042 2276 2045 2293
rect 2034 2273 2045 2276
rect 2034 2136 2037 2273
rect 2058 2266 2061 2326
rect 2070 2306 2073 2353
rect 2070 2303 2077 2306
rect 2050 2263 2061 2266
rect 2050 2213 2053 2263
rect 2074 2186 2077 2303
rect 2090 2223 2093 2356
rect 2114 2333 2117 2443
rect 2130 2376 2133 2503
rect 2154 2423 2157 2526
rect 2170 2413 2173 2526
rect 2178 2496 2181 2596
rect 2186 2533 2189 2566
rect 2186 2513 2189 2526
rect 2178 2493 2189 2496
rect 2126 2373 2133 2376
rect 2126 2326 2129 2373
rect 2122 2323 2129 2326
rect 2138 2323 2141 2336
rect 2082 2213 2101 2216
rect 2058 2183 2077 2186
rect 2034 2133 2045 2136
rect 2018 2123 2029 2126
rect 2002 2056 2005 2076
rect 2026 2056 2029 2123
rect 2002 2053 2013 2056
rect 1986 2043 1997 2046
rect 1954 1993 1961 1996
rect 1954 1976 1957 1993
rect 1914 1973 1925 1976
rect 1946 1973 1957 1976
rect 1914 1946 1917 1973
rect 1914 1943 1925 1946
rect 1890 1803 1893 1926
rect 1906 1856 1909 1936
rect 1902 1853 1909 1856
rect 1902 1776 1905 1853
rect 1922 1846 1925 1943
rect 1938 1933 1941 1956
rect 1914 1843 1925 1846
rect 1902 1773 1909 1776
rect 1890 1693 1893 1756
rect 1906 1703 1909 1773
rect 1874 1656 1877 1676
rect 1914 1673 1917 1843
rect 1930 1813 1933 1826
rect 1938 1806 1941 1926
rect 1946 1813 1949 1973
rect 1970 1953 1973 2016
rect 1978 1943 1981 2026
rect 1954 1853 1957 1936
rect 1986 1933 1989 2006
rect 1994 1933 1997 2043
rect 2010 1956 2013 2053
rect 2022 2053 2029 2056
rect 2022 2006 2025 2053
rect 2042 2046 2045 2133
rect 2058 2056 2061 2183
rect 2090 2133 2093 2206
rect 2098 2203 2101 2213
rect 2106 2203 2109 2296
rect 2122 2243 2125 2323
rect 2130 2236 2133 2256
rect 2122 2233 2133 2236
rect 2098 2133 2109 2136
rect 2082 2123 2101 2126
rect 2114 2123 2117 2216
rect 2058 2053 2077 2056
rect 2034 2043 2045 2046
rect 2034 2013 2037 2043
rect 2022 2003 2029 2006
rect 2002 1953 2013 1956
rect 1962 1923 1981 1926
rect 1978 1873 1981 1923
rect 1994 1863 1997 1926
rect 2002 1856 2005 1953
rect 2010 1906 2013 1936
rect 2010 1903 2017 1906
rect 1986 1853 2005 1856
rect 1874 1653 1881 1656
rect 1878 1556 1881 1653
rect 1898 1613 1901 1636
rect 1874 1553 1881 1556
rect 1890 1553 1893 1606
rect 1906 1573 1909 1606
rect 1914 1603 1917 1616
rect 1922 1593 1925 1806
rect 1934 1803 1941 1806
rect 1934 1746 1937 1803
rect 1930 1743 1937 1746
rect 1930 1586 1933 1743
rect 1938 1603 1941 1726
rect 1954 1666 1957 1806
rect 1962 1803 1965 1816
rect 1986 1766 1989 1853
rect 2014 1846 2017 1903
rect 2010 1843 2017 1846
rect 2010 1786 2013 1843
rect 2026 1813 2029 2003
rect 2050 1996 2053 2026
rect 2042 1993 2053 1996
rect 2042 1896 2045 1993
rect 2058 1973 2061 2026
rect 2066 2023 2069 2036
rect 2074 2016 2077 2053
rect 2066 2013 2077 2016
rect 2082 2013 2085 2116
rect 2042 1893 2053 1896
rect 2018 1793 2021 1806
rect 2034 1803 2037 1876
rect 2042 1803 2045 1826
rect 2010 1783 2021 1786
rect 1986 1763 1997 1766
rect 1994 1733 1997 1763
rect 2018 1696 2021 1783
rect 2010 1693 2021 1696
rect 1946 1663 1957 1666
rect 1946 1613 1949 1663
rect 1970 1613 1973 1646
rect 1930 1583 1941 1586
rect 1874 1523 1877 1553
rect 1882 1513 1885 1536
rect 1866 1503 1873 1506
rect 1870 1436 1873 1503
rect 1898 1466 1901 1536
rect 1922 1523 1925 1556
rect 1938 1516 1941 1583
rect 1978 1523 1981 1606
rect 1890 1463 1901 1466
rect 1930 1513 1941 1516
rect 1890 1446 1893 1463
rect 1930 1446 1933 1513
rect 1866 1433 1873 1436
rect 1886 1443 1893 1446
rect 1922 1443 1933 1446
rect 1866 1223 1869 1433
rect 1874 1333 1877 1416
rect 1886 1376 1889 1443
rect 1906 1403 1909 1416
rect 1922 1396 1925 1443
rect 1922 1393 1933 1396
rect 1886 1373 1893 1376
rect 1890 1353 1893 1373
rect 1874 1213 1877 1326
rect 1930 1253 1933 1393
rect 1954 1353 1957 1406
rect 1978 1336 1981 1426
rect 1986 1376 1989 1416
rect 1994 1413 1997 1436
rect 2002 1423 2005 1686
rect 2010 1586 2013 1693
rect 2026 1603 2029 1726
rect 2034 1613 2037 1796
rect 2050 1766 2053 1893
rect 2042 1763 2053 1766
rect 2042 1683 2045 1763
rect 2050 1613 2053 1646
rect 2010 1583 2021 1586
rect 2018 1456 2021 1583
rect 2042 1573 2045 1606
rect 2050 1556 2053 1606
rect 2042 1553 2053 1556
rect 2042 1506 2045 1553
rect 2058 1543 2061 1896
rect 2066 1773 2069 2013
rect 2090 2003 2093 2036
rect 2098 2023 2101 2066
rect 2122 2036 2125 2233
rect 2130 2206 2133 2226
rect 2130 2203 2141 2206
rect 2138 2136 2141 2203
rect 2130 2133 2141 2136
rect 2130 2113 2133 2133
rect 2114 2033 2125 2036
rect 2114 2006 2117 2033
rect 2106 2003 2117 2006
rect 2130 2005 2133 2016
rect 2106 1956 2109 2003
rect 2154 1966 2157 2246
rect 2162 2116 2165 2406
rect 2186 2256 2189 2493
rect 2210 2403 2213 2793
rect 2218 2716 2221 2806
rect 2226 2733 2229 2746
rect 2266 2726 2269 2813
rect 2290 2753 2293 2913
rect 2298 2813 2301 2826
rect 2282 2733 2293 2736
rect 2218 2713 2225 2716
rect 2222 2636 2225 2713
rect 2250 2683 2253 2726
rect 2266 2723 2293 2726
rect 2274 2666 2277 2716
rect 2218 2633 2225 2636
rect 2270 2663 2277 2666
rect 2218 2593 2221 2633
rect 2226 2566 2229 2616
rect 2226 2563 2237 2566
rect 2234 2496 2237 2563
rect 2258 2533 2261 2616
rect 2226 2493 2237 2496
rect 2226 2473 2229 2493
rect 2218 2316 2221 2406
rect 2234 2363 2237 2416
rect 2242 2403 2245 2416
rect 2250 2413 2253 2446
rect 2258 2406 2261 2526
rect 2270 2416 2273 2663
rect 2282 2423 2285 2656
rect 2306 2653 2309 2926
rect 2314 2923 2317 3023
rect 2322 2943 2325 3103
rect 2330 2936 2333 3076
rect 2322 2933 2333 2936
rect 2338 2933 2341 3193
rect 2362 3053 2365 3313
rect 2378 3246 2381 3266
rect 2374 3243 2381 3246
rect 2374 3196 2377 3243
rect 2386 3233 2405 3236
rect 2386 3223 2389 3233
rect 2386 3203 2389 3216
rect 2374 3193 2381 3196
rect 2378 3146 2381 3193
rect 2374 3143 2381 3146
rect 2322 2816 2325 2926
rect 2338 2906 2341 2926
rect 2334 2903 2341 2906
rect 2334 2826 2337 2903
rect 2334 2823 2341 2826
rect 2346 2823 2349 3036
rect 2374 3026 2377 3143
rect 2386 3073 2389 3136
rect 2354 3013 2357 3026
rect 2374 3023 2381 3026
rect 2362 3003 2365 3016
rect 2354 2916 2357 2936
rect 2370 2933 2373 3006
rect 2354 2913 2365 2916
rect 2318 2813 2325 2816
rect 2318 2756 2321 2813
rect 2318 2753 2325 2756
rect 2298 2566 2301 2646
rect 2314 2643 2317 2736
rect 2322 2733 2325 2753
rect 2330 2713 2333 2806
rect 2338 2803 2341 2823
rect 2362 2816 2365 2913
rect 2378 2833 2381 3023
rect 2354 2813 2365 2816
rect 2378 2813 2381 2826
rect 2354 2723 2357 2813
rect 2378 2716 2381 2736
rect 2370 2713 2381 2716
rect 2370 2636 2373 2713
rect 2370 2633 2381 2636
rect 2346 2613 2349 2626
rect 2378 2613 2381 2633
rect 2386 2596 2389 3056
rect 2394 2923 2397 3226
rect 2402 3213 2405 3233
rect 2410 3223 2413 3423
rect 2402 3013 2405 3166
rect 2410 3096 2413 3206
rect 2418 3183 2421 3476
rect 2426 3233 2429 3563
rect 2434 3483 2437 3536
rect 2450 3496 2453 3536
rect 2446 3493 2453 3496
rect 2446 3406 2449 3493
rect 2474 3486 2477 3606
rect 2482 3603 2485 3613
rect 2458 3413 2461 3486
rect 2470 3483 2477 3486
rect 2446 3403 2453 3406
rect 2426 3133 2429 3226
rect 2450 3223 2453 3403
rect 2470 3356 2473 3483
rect 2482 3383 2485 3576
rect 2490 3496 2493 3606
rect 2498 3593 2501 3693
rect 2514 3566 2517 3686
rect 2522 3676 2525 3726
rect 2522 3673 2541 3676
rect 2530 3613 2533 3666
rect 2538 3613 2541 3673
rect 2538 3593 2541 3606
rect 2514 3563 2525 3566
rect 2498 3513 2501 3526
rect 2490 3493 2497 3496
rect 2494 3366 2497 3493
rect 2522 3486 2525 3563
rect 2546 3536 2549 3916
rect 2570 3866 2573 3926
rect 2554 3863 2573 3866
rect 2554 3813 2557 3863
rect 2562 3786 2565 3856
rect 2582 3846 2585 3973
rect 2582 3843 2589 3846
rect 2570 3796 2573 3836
rect 2578 3813 2581 3826
rect 2586 3803 2589 3843
rect 2594 3813 2597 4036
rect 2602 4013 2605 4053
rect 2610 3903 2613 4073
rect 2618 4013 2621 4216
rect 2626 4126 2629 4313
rect 2642 4296 2645 4406
rect 2662 4356 2665 4423
rect 2638 4293 2645 4296
rect 2638 4226 2641 4293
rect 2650 4233 2653 4356
rect 2662 4353 2669 4356
rect 2658 4323 2661 4336
rect 2666 4306 2669 4353
rect 2674 4333 2677 4416
rect 2682 4413 2685 4446
rect 2698 4413 2701 4513
rect 2714 4436 2717 4526
rect 2706 4433 2717 4436
rect 2706 4406 2709 4433
rect 2730 4426 2733 4556
rect 2762 4533 2765 4546
rect 2826 4533 2829 4606
rect 2730 4423 2741 4426
rect 2682 4333 2685 4406
rect 2690 4403 2709 4406
rect 2662 4303 2669 4306
rect 2662 4236 2665 4303
rect 2674 4263 2677 4326
rect 2682 4266 2685 4326
rect 2682 4263 2693 4266
rect 2662 4233 2669 4236
rect 2638 4223 2645 4226
rect 2634 4143 2637 4206
rect 2626 4123 2633 4126
rect 2630 4036 2633 4123
rect 2626 4033 2633 4036
rect 2626 3986 2629 4033
rect 2642 4023 2645 4223
rect 2650 4213 2661 4216
rect 2650 4203 2653 4213
rect 2666 4206 2669 4233
rect 2658 4203 2669 4206
rect 2658 4133 2661 4203
rect 2674 4193 2677 4236
rect 2634 3993 2637 4016
rect 2642 3996 2645 4016
rect 2642 3993 2649 3996
rect 2626 3983 2637 3986
rect 2626 3833 2629 3926
rect 2570 3793 2581 3796
rect 2562 3783 2573 3786
rect 2554 3593 2557 3726
rect 2570 3723 2573 3783
rect 2578 3706 2581 3793
rect 2574 3703 2581 3706
rect 2574 3646 2577 3703
rect 2562 3623 2565 3646
rect 2570 3643 2577 3646
rect 2546 3533 2557 3536
rect 2514 3483 2525 3486
rect 2506 3373 2509 3406
rect 2490 3363 2497 3366
rect 2470 3353 2477 3356
rect 2474 3286 2477 3353
rect 2470 3283 2477 3286
rect 2450 3173 2453 3206
rect 2458 3193 2461 3226
rect 2470 3206 2473 3283
rect 2466 3203 2473 3206
rect 2482 3203 2485 3346
rect 2458 3143 2461 3186
rect 2410 3093 2417 3096
rect 2414 3006 2417 3093
rect 2410 3003 2417 3006
rect 2410 2966 2413 3003
rect 2406 2963 2413 2966
rect 2426 2966 2429 3106
rect 2466 3103 2469 3203
rect 2490 3196 2493 3363
rect 2498 3323 2501 3346
rect 2514 3283 2517 3483
rect 2498 3213 2501 3226
rect 2474 3193 2493 3196
rect 2498 3186 2501 3206
rect 2498 3183 2509 3186
rect 2490 3156 2493 3176
rect 2490 3153 2497 3156
rect 2474 3123 2477 3146
rect 2494 3096 2497 3153
rect 2490 3093 2497 3096
rect 2490 3076 2493 3093
rect 2482 3073 2493 3076
rect 2466 3013 2469 3036
rect 2482 3026 2485 3073
rect 2506 3046 2509 3183
rect 2522 3053 2525 3436
rect 2530 3403 2533 3416
rect 2538 3403 2541 3526
rect 2554 3436 2557 3533
rect 2546 3433 2557 3436
rect 2530 3323 2533 3376
rect 2538 3263 2541 3336
rect 2546 3246 2549 3433
rect 2570 3416 2573 3643
rect 2586 3636 2589 3726
rect 2594 3696 2597 3806
rect 2626 3753 2629 3816
rect 2634 3743 2637 3983
rect 2646 3866 2649 3993
rect 2642 3863 2649 3866
rect 2602 3713 2605 3726
rect 2594 3693 2601 3696
rect 2578 3633 2589 3636
rect 2578 3603 2581 3633
rect 2586 3603 2589 3626
rect 2598 3596 2601 3693
rect 2610 3623 2613 3726
rect 2618 3716 2621 3736
rect 2618 3713 2629 3716
rect 2626 3626 2629 3713
rect 2622 3623 2629 3626
rect 2554 3413 2573 3416
rect 2594 3593 2601 3596
rect 2594 3416 2597 3593
rect 2610 3583 2613 3616
rect 2622 3576 2625 3623
rect 2642 3613 2645 3863
rect 2658 3856 2661 3936
rect 2666 3873 2669 4016
rect 2682 3953 2685 4263
rect 2698 4223 2701 4326
rect 2706 4303 2709 4336
rect 2714 4333 2717 4346
rect 2722 4326 2725 4416
rect 2738 4356 2741 4423
rect 2794 4413 2797 4526
rect 2826 4513 2829 4526
rect 2842 4523 2845 4606
rect 2850 4523 2853 4536
rect 2858 4533 2861 4556
rect 2866 4516 2869 4536
rect 2890 4533 2893 4616
rect 2946 4553 2949 4616
rect 2970 4593 2973 4606
rect 2946 4543 2965 4546
rect 2858 4513 2869 4516
rect 2858 4496 2861 4513
rect 2850 4493 2861 4496
rect 2850 4436 2853 4493
rect 2874 4446 2877 4526
rect 2874 4443 2885 4446
rect 2850 4433 2861 4436
rect 2754 4373 2757 4406
rect 2770 4383 2773 4406
rect 2786 4363 2789 4386
rect 2714 4323 2725 4326
rect 2730 4353 2741 4356
rect 2690 4123 2693 4216
rect 2714 4213 2717 4323
rect 2730 4283 2733 4353
rect 2738 4313 2741 4326
rect 2746 4253 2749 4336
rect 2754 4323 2757 4336
rect 2762 4333 2765 4356
rect 2770 4323 2773 4336
rect 2778 4313 2781 4326
rect 2786 4296 2789 4336
rect 2794 4323 2797 4336
rect 2778 4293 2789 4296
rect 2730 4213 2749 4216
rect 2730 4203 2733 4213
rect 2738 4123 2741 4206
rect 2754 4203 2757 4236
rect 2778 4226 2781 4293
rect 2802 4246 2805 4366
rect 2818 4333 2821 4346
rect 2826 4333 2829 4376
rect 2850 4373 2853 4416
rect 2834 4313 2837 4326
rect 2842 4273 2845 4336
rect 2850 4323 2853 4336
rect 2858 4333 2861 4433
rect 2866 4403 2869 4416
rect 2882 4366 2885 4443
rect 2874 4363 2885 4366
rect 2866 4333 2869 4346
rect 2874 4326 2877 4363
rect 2866 4323 2877 4326
rect 2882 4343 2901 4346
rect 2882 4323 2885 4343
rect 2798 4243 2805 4246
rect 2778 4223 2789 4226
rect 2762 4106 2765 4206
rect 2786 4163 2789 4223
rect 2798 4176 2801 4243
rect 2810 4213 2813 4226
rect 2826 4213 2829 4236
rect 2834 4193 2837 4206
rect 2794 4173 2801 4176
rect 2754 4103 2765 4106
rect 2754 4056 2757 4103
rect 2794 4096 2797 4173
rect 2842 4133 2845 4256
rect 2850 4213 2853 4226
rect 2866 4213 2869 4323
rect 2890 4316 2893 4336
rect 2898 4333 2901 4343
rect 2906 4316 2909 4526
rect 2914 4396 2917 4416
rect 2922 4403 2925 4436
rect 2930 4413 2933 4526
rect 2946 4523 2949 4543
rect 2954 4523 2957 4536
rect 2962 4533 2965 4543
rect 2962 4443 2965 4526
rect 2970 4523 2973 4556
rect 3002 4503 3005 4526
rect 2954 4413 2957 4426
rect 2930 4396 2933 4406
rect 2914 4393 2933 4396
rect 2962 4353 2965 4436
rect 2994 4413 2997 4426
rect 3042 4356 3045 4596
rect 3098 4573 3101 4616
rect 3114 4543 3133 4546
rect 3058 4513 3061 4526
rect 3082 4483 3085 4536
rect 3114 4533 3117 4543
rect 3098 4513 3101 4526
rect 3106 4493 3109 4526
rect 3026 4353 3045 4356
rect 2890 4313 2909 4316
rect 2890 4253 2893 4313
rect 2914 4263 2917 4326
rect 2938 4313 2941 4326
rect 2946 4323 2949 4346
rect 2978 4313 2981 4326
rect 2874 4206 2877 4216
rect 2906 4213 2909 4236
rect 2866 4203 2877 4206
rect 2954 4203 2957 4226
rect 2866 4163 2869 4203
rect 2882 4133 2885 4146
rect 2770 4093 2797 4096
rect 2754 4053 2765 4056
rect 2762 4033 2765 4053
rect 2682 3933 2685 3946
rect 2714 3866 2717 4006
rect 2730 3993 2733 4006
rect 2746 3926 2749 4016
rect 2770 3973 2773 4093
rect 2818 4003 2821 4016
rect 2730 3913 2733 3926
rect 2746 3923 2757 3926
rect 2706 3863 2717 3866
rect 2658 3853 2665 3856
rect 2662 3776 2665 3853
rect 2658 3773 2665 3776
rect 2618 3573 2625 3576
rect 2618 3526 2621 3573
rect 2610 3523 2621 3526
rect 2634 3526 2637 3606
rect 2634 3523 2641 3526
rect 2610 3456 2613 3523
rect 2610 3453 2621 3456
rect 2618 3433 2621 3453
rect 2594 3413 2605 3416
rect 2610 3413 2613 3426
rect 2554 3316 2557 3413
rect 2562 3333 2565 3406
rect 2554 3313 2565 3316
rect 2562 3246 2565 3313
rect 2538 3243 2549 3246
rect 2554 3243 2565 3246
rect 2538 3196 2541 3243
rect 2554 3203 2557 3243
rect 2538 3193 2549 3196
rect 2546 3173 2549 3193
rect 2498 3043 2509 3046
rect 2554 3043 2557 3136
rect 2562 3103 2565 3126
rect 2570 3056 2573 3226
rect 2578 3123 2581 3356
rect 2586 3333 2589 3346
rect 2594 3323 2597 3406
rect 2602 3306 2605 3413
rect 2598 3303 2605 3306
rect 2586 3213 2589 3256
rect 2598 3236 2601 3303
rect 2598 3233 2605 3236
rect 2594 3196 2597 3216
rect 2590 3193 2597 3196
rect 2590 3106 2593 3193
rect 2602 3116 2605 3233
rect 2610 3173 2613 3386
rect 2618 3353 2621 3416
rect 2626 3403 2629 3516
rect 2638 3466 2641 3523
rect 2634 3463 2641 3466
rect 2634 3443 2637 3463
rect 2634 3413 2637 3426
rect 2626 3213 2629 3336
rect 2642 3333 2645 3406
rect 2650 3393 2653 3616
rect 2658 3603 2661 3773
rect 2674 3613 2677 3826
rect 2682 3736 2685 3816
rect 2706 3803 2709 3863
rect 2730 3813 2733 3826
rect 2706 3766 2709 3796
rect 2722 3786 2725 3806
rect 2738 3803 2741 3876
rect 2754 3846 2757 3923
rect 2778 3896 2781 3916
rect 2746 3843 2757 3846
rect 2770 3893 2781 3896
rect 2770 3846 2773 3893
rect 2770 3843 2781 3846
rect 2746 3813 2749 3843
rect 2762 3813 2765 3826
rect 2754 3793 2757 3806
rect 2722 3783 2733 3786
rect 2702 3763 2709 3766
rect 2682 3733 2693 3736
rect 2690 3603 2693 3733
rect 2702 3646 2705 3763
rect 2702 3643 2709 3646
rect 2698 3613 2701 3626
rect 2674 3466 2677 3536
rect 2706 3516 2709 3643
rect 2714 3603 2717 3756
rect 2730 3706 2733 3783
rect 2762 3756 2765 3806
rect 2778 3803 2781 3843
rect 2786 3813 2789 3926
rect 2802 3813 2805 3926
rect 2794 3793 2797 3806
rect 2722 3703 2733 3706
rect 2746 3753 2765 3756
rect 2722 3683 2725 3703
rect 2722 3613 2725 3626
rect 2746 3576 2749 3753
rect 2746 3573 2757 3576
rect 2706 3513 2717 3516
rect 2714 3486 2717 3513
rect 2706 3483 2717 3486
rect 2674 3463 2685 3466
rect 2658 3246 2661 3406
rect 2658 3243 2669 3246
rect 2642 3203 2645 3226
rect 2618 3133 2621 3146
rect 2602 3113 2613 3116
rect 2590 3103 2597 3106
rect 2566 3053 2573 3056
rect 2482 3023 2493 3026
rect 2442 3003 2453 3006
rect 2426 2963 2433 2966
rect 2406 2906 2409 2963
rect 2406 2903 2413 2906
rect 2410 2883 2413 2903
rect 2430 2886 2433 2963
rect 2426 2883 2433 2886
rect 2394 2813 2397 2866
rect 2394 2783 2397 2806
rect 2402 2616 2405 2836
rect 2410 2803 2413 2856
rect 2410 2713 2413 2726
rect 2418 2663 2421 2816
rect 2426 2646 2429 2883
rect 2434 2776 2437 2826
rect 2442 2803 2445 2926
rect 2450 2813 2453 3003
rect 2474 2933 2477 2946
rect 2490 2933 2493 3023
rect 2466 2813 2469 2886
rect 2490 2823 2493 2926
rect 2498 2916 2501 3043
rect 2506 2933 2509 3006
rect 2498 2913 2505 2916
rect 2502 2816 2505 2913
rect 2498 2813 2505 2816
rect 2434 2773 2445 2776
rect 2434 2716 2437 2766
rect 2442 2723 2445 2773
rect 2434 2713 2445 2716
rect 2422 2643 2429 2646
rect 2402 2613 2413 2616
rect 2378 2593 2389 2596
rect 2298 2563 2309 2566
rect 2306 2496 2309 2563
rect 2354 2523 2357 2546
rect 2378 2516 2381 2593
rect 2394 2523 2397 2606
rect 2410 2516 2413 2613
rect 2378 2513 2389 2516
rect 2298 2493 2309 2496
rect 2298 2436 2301 2493
rect 2290 2433 2301 2436
rect 2270 2413 2277 2416
rect 2250 2403 2261 2406
rect 2242 2333 2253 2336
rect 2226 2323 2245 2326
rect 2258 2323 2261 2366
rect 2178 2253 2189 2256
rect 2210 2313 2221 2316
rect 2178 2233 2181 2253
rect 2186 2213 2189 2226
rect 2210 2216 2213 2313
rect 2210 2213 2221 2216
rect 2218 2193 2221 2213
rect 2162 2113 2169 2116
rect 2166 1996 2169 2113
rect 2194 2066 2197 2136
rect 2210 2133 2213 2146
rect 2202 2113 2205 2126
rect 2218 2123 2221 2136
rect 2226 2126 2229 2226
rect 2234 2203 2237 2323
rect 2242 2133 2245 2316
rect 2266 2253 2269 2386
rect 2258 2213 2261 2226
rect 2258 2203 2269 2206
rect 2226 2123 2237 2126
rect 2226 2096 2229 2116
rect 2178 2063 2197 2066
rect 2218 2093 2229 2096
rect 2178 2013 2181 2063
rect 2194 2026 2197 2046
rect 2218 2036 2221 2093
rect 2234 2043 2237 2123
rect 2218 2033 2229 2036
rect 2194 2023 2205 2026
rect 2166 1993 2173 1996
rect 2146 1963 2157 1966
rect 2106 1953 2117 1956
rect 2074 1756 2077 1806
rect 2066 1753 2077 1756
rect 2066 1603 2069 1753
rect 2074 1676 2077 1746
rect 2082 1696 2085 1806
rect 2090 1803 2093 1936
rect 2114 1933 2117 1953
rect 2098 1813 2101 1866
rect 2106 1796 2109 1856
rect 2114 1803 2117 1926
rect 2146 1916 2149 1963
rect 2146 1913 2157 1916
rect 2154 1893 2157 1913
rect 2170 1896 2173 1993
rect 2202 1976 2205 2023
rect 2226 2013 2229 2033
rect 2234 1996 2237 2026
rect 2194 1973 2205 1976
rect 2226 1993 2237 1996
rect 2162 1893 2173 1896
rect 2162 1873 2165 1893
rect 2186 1876 2189 1926
rect 2178 1873 2189 1876
rect 2178 1826 2181 1873
rect 2122 1813 2141 1816
rect 2130 1796 2133 1806
rect 2138 1803 2141 1813
rect 2090 1723 2093 1796
rect 2106 1793 2133 1796
rect 2146 1776 2149 1826
rect 2178 1823 2189 1826
rect 2138 1773 2149 1776
rect 2106 1733 2109 1746
rect 2138 1706 2141 1773
rect 2154 1753 2157 1816
rect 2186 1803 2189 1823
rect 2194 1813 2197 1973
rect 2226 1916 2229 1993
rect 2202 1896 2205 1916
rect 2226 1913 2237 1916
rect 2202 1893 2213 1896
rect 2210 1846 2213 1893
rect 2202 1843 2213 1846
rect 2202 1813 2205 1843
rect 2154 1713 2157 1726
rect 2138 1703 2149 1706
rect 2082 1693 2093 1696
rect 2074 1673 2081 1676
rect 2078 1616 2081 1673
rect 2074 1613 2081 1616
rect 2042 1503 2053 1506
rect 2010 1453 2021 1456
rect 1986 1373 1997 1376
rect 1978 1333 1989 1336
rect 1970 1223 1973 1326
rect 1978 1253 1981 1326
rect 1986 1246 1989 1333
rect 1994 1323 1997 1373
rect 2010 1356 2013 1453
rect 2050 1436 2053 1503
rect 2026 1433 2053 1436
rect 2026 1376 2029 1433
rect 2050 1393 2053 1406
rect 2074 1393 2077 1613
rect 2090 1596 2093 1693
rect 2090 1593 2101 1596
rect 2098 1546 2101 1593
rect 2098 1543 2105 1546
rect 2102 1496 2105 1543
rect 2114 1523 2117 1606
rect 2122 1603 2125 1616
rect 2138 1613 2141 1646
rect 2130 1573 2133 1606
rect 2146 1573 2149 1703
rect 2154 1556 2157 1606
rect 2162 1576 2165 1616
rect 2170 1593 2173 1736
rect 2218 1733 2221 1816
rect 2226 1813 2229 1826
rect 2178 1603 2181 1636
rect 2162 1573 2169 1576
rect 2098 1493 2105 1496
rect 2098 1423 2101 1493
rect 2138 1486 2141 1556
rect 2150 1553 2157 1556
rect 2150 1506 2153 1553
rect 2166 1516 2169 1573
rect 2166 1513 2173 1516
rect 2150 1503 2157 1506
rect 2122 1483 2141 1486
rect 2098 1393 2101 1416
rect 2026 1373 2037 1376
rect 2010 1353 2029 1356
rect 2002 1306 2005 1336
rect 1978 1243 1989 1246
rect 1998 1303 2005 1306
rect 1930 1193 1933 1216
rect 1866 1133 1869 1146
rect 1954 1143 1957 1206
rect 1970 1173 1973 1206
rect 1978 1126 1981 1243
rect 1998 1236 2001 1303
rect 1834 1013 1837 1036
rect 1842 1033 1845 1096
rect 1850 1093 1861 1096
rect 1858 1046 1861 1093
rect 1850 1043 1861 1046
rect 1850 1023 1853 1043
rect 1826 1003 1845 1006
rect 1818 876 1821 936
rect 1826 883 1829 936
rect 1842 886 1845 1003
rect 1866 903 1869 1016
rect 1890 943 1893 1126
rect 1914 1113 1917 1126
rect 1970 1123 1981 1126
rect 1986 1233 2001 1236
rect 1970 1026 1973 1123
rect 1986 1106 1989 1233
rect 1982 1103 1989 1106
rect 1982 1046 1985 1103
rect 1982 1043 1989 1046
rect 1970 1023 1981 1026
rect 1914 1013 1933 1016
rect 1978 1006 1981 1023
rect 1986 1013 1989 1043
rect 1906 946 1909 1006
rect 1922 993 1925 1006
rect 1906 943 1917 946
rect 1874 913 1877 926
rect 1834 883 1845 886
rect 1818 873 1829 876
rect 1794 833 1801 836
rect 1794 756 1797 833
rect 1802 793 1805 816
rect 1810 783 1813 836
rect 1818 823 1821 866
rect 1826 813 1829 873
rect 1834 863 1837 883
rect 1890 876 1893 936
rect 1914 923 1917 943
rect 1938 906 1941 946
rect 1970 923 1973 1006
rect 1978 1003 1985 1006
rect 1930 903 1941 906
rect 1890 873 1909 876
rect 1858 813 1861 826
rect 1906 786 1909 873
rect 1930 846 1933 903
rect 1930 843 1941 846
rect 1922 786 1925 806
rect 1906 783 1925 786
rect 1794 753 1805 756
rect 1794 733 1797 746
rect 1794 653 1797 726
rect 1802 693 1805 753
rect 1882 733 1885 756
rect 1906 753 1909 783
rect 1938 736 1941 843
rect 1938 733 1945 736
rect 1954 733 1957 916
rect 1982 906 1985 1003
rect 1994 916 1997 1216
rect 2002 1213 2005 1226
rect 2010 1213 2013 1336
rect 2010 1193 2013 1206
rect 2002 1156 2005 1176
rect 2018 1173 2021 1346
rect 2002 1153 2009 1156
rect 2006 1026 2009 1153
rect 2026 1123 2029 1353
rect 2034 1233 2037 1373
rect 2002 1023 2009 1026
rect 2002 1003 2005 1023
rect 2018 1013 2021 1116
rect 2026 1003 2029 1116
rect 2034 1013 2037 1206
rect 2042 1116 2045 1386
rect 2050 1323 2053 1336
rect 2058 1333 2061 1356
rect 2058 1306 2061 1326
rect 2050 1123 2053 1306
rect 2058 1303 2065 1306
rect 2062 1246 2065 1303
rect 2058 1243 2065 1246
rect 2058 1213 2061 1243
rect 2074 1223 2077 1336
rect 2090 1333 2093 1346
rect 2098 1326 2101 1336
rect 2082 1323 2101 1326
rect 2098 1313 2101 1323
rect 2098 1213 2101 1226
rect 2074 1143 2077 1206
rect 2042 1113 2053 1116
rect 2026 933 2029 946
rect 1994 913 2001 916
rect 1982 903 1989 906
rect 1978 803 1981 886
rect 1978 746 1981 766
rect 1970 743 1981 746
rect 1834 713 1837 726
rect 1802 666 1805 686
rect 1802 663 1813 666
rect 1810 576 1813 663
rect 1802 573 1813 576
rect 1698 513 1709 516
rect 1762 513 1773 516
rect 1778 513 1781 526
rect 1786 523 1789 536
rect 1666 493 1677 496
rect 1674 426 1677 493
rect 1618 413 1629 416
rect 1634 413 1637 426
rect 1618 363 1621 413
rect 1626 393 1629 406
rect 1618 306 1621 326
rect 1614 303 1621 306
rect 1614 236 1617 303
rect 1614 233 1621 236
rect 1626 233 1629 386
rect 1642 353 1645 406
rect 1650 333 1653 426
rect 1666 423 1677 426
rect 1658 353 1661 416
rect 1658 333 1661 346
rect 1666 333 1669 423
rect 1674 333 1677 406
rect 1698 403 1701 513
rect 1762 426 1765 513
rect 1794 506 1797 536
rect 1802 523 1805 573
rect 1826 536 1829 616
rect 1786 503 1797 506
rect 1706 383 1709 406
rect 1722 393 1725 416
rect 1738 413 1741 426
rect 1762 423 1773 426
rect 1690 333 1693 366
rect 1650 313 1653 326
rect 1610 166 1613 216
rect 1618 203 1621 233
rect 1634 213 1637 306
rect 1658 226 1661 326
rect 1666 303 1669 326
rect 1730 323 1733 406
rect 1746 366 1749 406
rect 1770 403 1773 423
rect 1778 383 1781 406
rect 1738 363 1749 366
rect 1642 223 1669 226
rect 1642 213 1645 223
rect 1650 213 1661 216
rect 1666 213 1669 223
rect 1674 213 1685 216
rect 1610 163 1621 166
rect 1618 153 1621 163
rect 1626 146 1629 206
rect 1642 203 1653 206
rect 1642 183 1645 203
rect 1626 143 1637 146
rect 1602 123 1605 136
rect 1634 123 1637 143
rect 1658 133 1661 206
rect 1682 133 1685 196
rect 1690 183 1693 236
rect 1738 203 1741 363
rect 1786 323 1789 503
rect 1794 266 1797 346
rect 1786 263 1797 266
rect 1778 216 1781 256
rect 1762 213 1781 216
rect 1730 123 1733 136
rect 1754 133 1757 206
rect 1770 183 1773 206
rect 1778 123 1781 206
rect 1786 183 1789 263
rect 1810 253 1813 536
rect 1826 533 1837 536
rect 1818 503 1821 526
rect 1834 516 1837 533
rect 1826 413 1829 516
rect 1834 513 1841 516
rect 1850 513 1853 606
rect 1838 446 1841 513
rect 1834 443 1841 446
rect 1834 403 1837 443
rect 1842 413 1845 426
rect 1850 403 1853 496
rect 1866 366 1869 576
rect 1882 436 1885 556
rect 1898 526 1901 646
rect 1894 523 1901 526
rect 1930 523 1933 726
rect 1942 636 1945 733
rect 1970 676 1973 743
rect 1986 696 1989 903
rect 1998 816 2001 913
rect 1994 813 2001 816
rect 2010 813 2013 926
rect 2034 923 2037 1006
rect 2042 933 2045 1086
rect 2050 906 2053 1113
rect 2058 1106 2061 1126
rect 2058 1103 2069 1106
rect 2066 1046 2069 1103
rect 2090 1066 2093 1126
rect 2098 1123 2101 1136
rect 2106 1123 2109 1366
rect 2122 1346 2125 1483
rect 2138 1353 2141 1446
rect 2154 1383 2157 1503
rect 2162 1396 2165 1416
rect 2170 1413 2173 1513
rect 2178 1506 2181 1586
rect 2186 1523 2189 1606
rect 2194 1603 2197 1716
rect 2218 1696 2221 1726
rect 2210 1693 2221 1696
rect 2210 1636 2213 1693
rect 2210 1633 2221 1636
rect 2218 1616 2221 1633
rect 2202 1613 2221 1616
rect 2210 1583 2213 1606
rect 2226 1603 2229 1806
rect 2234 1596 2237 1913
rect 2250 1886 2253 2126
rect 2274 2093 2277 2413
rect 2290 2373 2293 2433
rect 2282 2213 2285 2326
rect 2298 2296 2301 2426
rect 2314 2356 2317 2476
rect 2362 2426 2365 2446
rect 2338 2413 2341 2426
rect 2354 2423 2365 2426
rect 2354 2376 2357 2423
rect 2354 2373 2365 2376
rect 2314 2353 2325 2356
rect 2322 2333 2325 2353
rect 2298 2293 2309 2296
rect 2306 2226 2309 2293
rect 2346 2266 2349 2326
rect 2298 2223 2309 2226
rect 2330 2263 2349 2266
rect 2298 2153 2301 2223
rect 2282 2056 2285 2126
rect 2298 2123 2301 2136
rect 2306 2123 2309 2206
rect 2314 2173 2317 2206
rect 2330 2203 2333 2263
rect 2338 2213 2357 2216
rect 2282 2053 2293 2056
rect 2274 1923 2277 2016
rect 2290 2013 2293 2053
rect 2298 2033 2301 2066
rect 2306 2013 2309 2026
rect 2250 1883 2257 1886
rect 2242 1633 2245 1876
rect 2254 1786 2257 1883
rect 2250 1783 2257 1786
rect 2250 1723 2253 1783
rect 2258 1716 2261 1766
rect 2254 1713 2261 1716
rect 2254 1666 2257 1713
rect 2250 1663 2257 1666
rect 2250 1603 2253 1663
rect 2266 1643 2269 1856
rect 2274 1793 2277 1806
rect 2274 1723 2277 1756
rect 2282 1733 2285 1826
rect 2290 1803 2293 1816
rect 2194 1523 2197 1576
rect 2218 1566 2221 1596
rect 2214 1563 2221 1566
rect 2226 1593 2237 1596
rect 2178 1503 2189 1506
rect 2186 1436 2189 1503
rect 2202 1443 2205 1546
rect 2214 1496 2217 1563
rect 2226 1503 2229 1593
rect 2250 1533 2253 1596
rect 2274 1593 2277 1616
rect 2258 1523 2277 1526
rect 2214 1493 2221 1496
rect 2178 1433 2189 1436
rect 2178 1403 2181 1433
rect 2194 1413 2213 1416
rect 2162 1393 2181 1396
rect 2186 1393 2189 1406
rect 2194 1403 2205 1406
rect 2210 1403 2213 1413
rect 2122 1343 2133 1346
rect 2114 1303 2117 1326
rect 2130 1316 2133 1343
rect 2122 1313 2133 1316
rect 2122 1256 2125 1313
rect 2138 1303 2141 1326
rect 2118 1253 2125 1256
rect 2118 1166 2121 1253
rect 2118 1163 2125 1166
rect 2122 1146 2125 1163
rect 2122 1143 2133 1146
rect 2090 1063 2101 1066
rect 2114 1063 2117 1136
rect 2042 903 2053 906
rect 2058 1043 2069 1046
rect 1994 793 1997 813
rect 2018 763 2021 826
rect 2002 733 2005 756
rect 1986 693 1997 696
rect 1970 673 1981 676
rect 1938 633 1945 636
rect 1894 436 1897 523
rect 1938 516 1941 633
rect 1946 576 1949 616
rect 1946 573 1965 576
rect 1946 523 1949 536
rect 1954 523 1957 566
rect 1962 533 1965 573
rect 1978 533 1981 673
rect 1994 636 1997 693
rect 1990 633 1997 636
rect 1990 546 1993 633
rect 2002 563 2005 616
rect 1986 543 1993 546
rect 1938 513 1965 516
rect 1874 433 1885 436
rect 1890 433 1897 436
rect 1874 413 1877 433
rect 1890 416 1893 433
rect 1886 413 1893 416
rect 1862 363 1869 366
rect 1826 313 1829 326
rect 1834 213 1837 336
rect 1842 303 1845 326
rect 1850 313 1853 326
rect 1862 316 1865 363
rect 1886 356 1889 413
rect 1886 353 1893 356
rect 1874 323 1877 336
rect 1862 313 1869 316
rect 1866 256 1869 313
rect 1866 253 1873 256
rect 1870 206 1873 253
rect 1882 213 1885 336
rect 1890 306 1893 353
rect 1898 316 1901 416
rect 1906 323 1909 506
rect 1922 403 1925 416
rect 1922 323 1925 396
rect 1946 386 1949 506
rect 1962 466 1965 513
rect 1942 383 1949 386
rect 1954 463 1965 466
rect 1898 313 1909 316
rect 1890 303 1901 306
rect 1802 193 1805 206
rect 1866 203 1873 206
rect 1866 183 1869 203
rect 1794 133 1797 146
rect 1842 123 1845 136
rect 1890 123 1893 206
rect 1898 193 1901 303
rect 1906 296 1909 313
rect 1906 293 1917 296
rect 1914 236 1917 293
rect 1906 233 1917 236
rect 1906 133 1909 233
rect 1930 216 1933 336
rect 1942 236 1945 383
rect 1942 233 1949 236
rect 1914 213 1933 216
rect 1914 163 1917 206
rect 1938 133 1941 206
rect 1946 173 1949 233
rect 1954 203 1957 463
rect 1962 323 1965 436
rect 1970 413 1973 426
rect 1986 393 1989 543
rect 1994 486 1997 526
rect 2002 503 2005 526
rect 1994 483 2001 486
rect 1998 416 2001 483
rect 1994 413 2001 416
rect 1994 386 1997 413
rect 1986 383 1997 386
rect 1970 313 1973 336
rect 1986 326 1989 383
rect 1978 323 1989 326
rect 1978 303 1981 323
rect 1994 213 1997 336
rect 2002 323 2005 396
rect 2010 333 2013 526
rect 2018 413 2021 546
rect 2026 443 2029 866
rect 2042 846 2045 903
rect 2042 843 2053 846
rect 2050 823 2053 843
rect 2058 816 2061 1043
rect 2042 813 2061 816
rect 2034 723 2037 806
rect 2026 413 2029 436
rect 2026 356 2029 406
rect 2018 353 2029 356
rect 2002 296 2005 316
rect 2002 293 2009 296
rect 2006 226 2009 293
rect 2002 223 2009 226
rect 2002 206 2005 223
rect 1970 193 1973 206
rect 1994 203 2005 206
rect 1946 113 1949 126
rect 1986 123 1989 146
rect 1282 93 1293 96
rect 1282 53 1285 93
rect 1994 83 1997 203
rect 2002 123 2005 176
rect 2010 113 2013 136
rect 2018 126 2021 353
rect 2034 313 2037 716
rect 2042 613 2045 806
rect 2058 796 2061 806
rect 2066 803 2069 1026
rect 2098 1013 2101 1063
rect 2130 1056 2133 1143
rect 2122 1053 2133 1056
rect 2106 1033 2109 1046
rect 2122 1023 2125 1053
rect 2122 1003 2125 1016
rect 2146 1013 2149 1336
rect 2154 1323 2157 1336
rect 2162 1313 2165 1326
rect 2170 1316 2173 1336
rect 2178 1333 2181 1393
rect 2218 1376 2221 1493
rect 2202 1373 2221 1376
rect 2170 1313 2181 1316
rect 2162 1266 2165 1286
rect 2158 1263 2165 1266
rect 2158 1206 2161 1263
rect 2178 1246 2181 1313
rect 2202 1266 2205 1373
rect 2226 1323 2229 1406
rect 2234 1396 2237 1416
rect 2234 1393 2241 1396
rect 2238 1316 2241 1393
rect 2250 1336 2253 1426
rect 2258 1413 2261 1506
rect 2266 1403 2269 1523
rect 2274 1413 2277 1426
rect 2250 1333 2269 1336
rect 2282 1333 2285 1726
rect 2290 1723 2293 1756
rect 2298 1746 2301 1916
rect 2314 1763 2317 2156
rect 2338 2133 2341 2213
rect 2346 2193 2349 2206
rect 2330 1986 2333 2126
rect 2346 2113 2349 2136
rect 2362 2133 2365 2373
rect 2386 2366 2389 2513
rect 2402 2513 2413 2516
rect 2402 2456 2405 2513
rect 2398 2453 2405 2456
rect 2398 2406 2401 2453
rect 2410 2413 2413 2446
rect 2422 2436 2425 2643
rect 2434 2526 2437 2706
rect 2442 2533 2445 2713
rect 2450 2623 2453 2736
rect 2466 2733 2469 2806
rect 2482 2746 2485 2806
rect 2478 2743 2485 2746
rect 2498 2746 2501 2813
rect 2498 2743 2505 2746
rect 2458 2713 2461 2726
rect 2458 2576 2461 2616
rect 2466 2583 2469 2686
rect 2458 2573 2469 2576
rect 2458 2533 2461 2546
rect 2434 2523 2445 2526
rect 2422 2433 2429 2436
rect 2398 2403 2405 2406
rect 2402 2383 2405 2403
rect 2418 2383 2421 2416
rect 2426 2386 2429 2433
rect 2434 2403 2437 2486
rect 2426 2383 2433 2386
rect 2386 2363 2393 2366
rect 2390 2286 2393 2363
rect 2386 2283 2393 2286
rect 2386 2216 2389 2283
rect 2378 2213 2389 2216
rect 2346 2076 2349 2096
rect 2342 2073 2349 2076
rect 2342 1996 2345 2073
rect 2354 2033 2357 2126
rect 2370 2123 2373 2136
rect 2378 2033 2381 2213
rect 2402 2203 2405 2326
rect 2410 2323 2413 2336
rect 2418 2306 2421 2356
rect 2414 2303 2421 2306
rect 2414 2236 2417 2303
rect 2430 2296 2433 2383
rect 2426 2293 2433 2296
rect 2414 2233 2421 2236
rect 2410 2193 2413 2216
rect 2402 2096 2405 2146
rect 2418 2123 2421 2233
rect 2394 2093 2405 2096
rect 2394 2046 2397 2093
rect 2394 2043 2405 2046
rect 2354 2006 2357 2026
rect 2394 2006 2397 2026
rect 2402 2013 2405 2043
rect 2354 2003 2365 2006
rect 2342 1993 2349 1996
rect 2326 1983 2333 1986
rect 2326 1896 2329 1983
rect 2338 1903 2341 1976
rect 2326 1893 2333 1896
rect 2330 1873 2333 1893
rect 2338 1793 2341 1816
rect 2338 1756 2341 1776
rect 2334 1753 2341 1756
rect 2298 1743 2317 1746
rect 2298 1713 2301 1736
rect 2306 1723 2309 1736
rect 2314 1706 2317 1743
rect 2298 1703 2317 1706
rect 2290 1533 2293 1646
rect 2298 1516 2301 1703
rect 2322 1626 2325 1716
rect 2334 1706 2337 1753
rect 2346 1713 2349 1993
rect 2362 1946 2365 2003
rect 2354 1943 2365 1946
rect 2386 2003 2397 2006
rect 2386 1946 2389 2003
rect 2386 1943 2397 1946
rect 2354 1753 2357 1943
rect 2362 1773 2365 1876
rect 2370 1853 2373 1926
rect 2394 1886 2397 1943
rect 2402 1933 2405 1946
rect 2386 1883 2397 1886
rect 2386 1723 2389 1883
rect 2410 1843 2413 2086
rect 2426 2063 2429 2293
rect 2434 2106 2437 2216
rect 2442 2146 2445 2523
rect 2450 2506 2453 2526
rect 2466 2523 2469 2573
rect 2478 2506 2481 2743
rect 2450 2503 2461 2506
rect 2458 2436 2461 2503
rect 2450 2433 2461 2436
rect 2474 2503 2481 2506
rect 2450 2413 2453 2433
rect 2474 2396 2477 2503
rect 2490 2443 2493 2736
rect 2502 2626 2505 2743
rect 2514 2703 2517 2936
rect 2522 2906 2525 3026
rect 2554 2956 2557 3016
rect 2538 2953 2557 2956
rect 2538 2933 2541 2953
rect 2566 2946 2569 3053
rect 2566 2943 2573 2946
rect 2546 2923 2549 2936
rect 2522 2903 2533 2906
rect 2562 2903 2565 2926
rect 2570 2916 2573 2943
rect 2578 2933 2581 2946
rect 2594 2933 2597 3103
rect 2610 2956 2613 3113
rect 2626 3103 2629 3166
rect 2634 3133 2637 3146
rect 2642 3123 2645 3136
rect 2650 3123 2653 3136
rect 2602 2953 2613 2956
rect 2570 2913 2581 2916
rect 2530 2836 2533 2903
rect 2578 2856 2581 2913
rect 2522 2833 2533 2836
rect 2562 2853 2581 2856
rect 2522 2776 2525 2833
rect 2522 2773 2529 2776
rect 2526 2696 2529 2773
rect 2538 2733 2541 2816
rect 2554 2723 2557 2816
rect 2562 2766 2565 2853
rect 2594 2813 2597 2856
rect 2562 2763 2569 2766
rect 2566 2716 2569 2763
rect 2578 2723 2581 2736
rect 2498 2623 2505 2626
rect 2522 2693 2529 2696
rect 2562 2713 2569 2716
rect 2498 2563 2501 2623
rect 2506 2593 2509 2606
rect 2522 2566 2525 2693
rect 2562 2566 2565 2713
rect 2594 2693 2597 2736
rect 2602 2676 2605 2953
rect 2618 2853 2621 2936
rect 2626 2933 2629 3016
rect 2626 2906 2629 2926
rect 2634 2923 2637 2946
rect 2626 2903 2633 2906
rect 2630 2846 2633 2903
rect 2626 2843 2633 2846
rect 2626 2813 2629 2843
rect 2626 2793 2629 2806
rect 2642 2786 2645 2926
rect 2626 2783 2645 2786
rect 2610 2733 2613 2756
rect 2594 2673 2605 2676
rect 2570 2593 2573 2616
rect 2594 2576 2597 2673
rect 2610 2613 2613 2726
rect 2618 2716 2621 2726
rect 2626 2723 2629 2783
rect 2618 2713 2629 2716
rect 2610 2583 2613 2606
rect 2594 2573 2601 2576
rect 2514 2563 2525 2566
rect 2514 2523 2517 2563
rect 2466 2393 2477 2396
rect 2466 2306 2469 2393
rect 2490 2313 2493 2416
rect 2498 2403 2501 2516
rect 2538 2513 2541 2526
rect 2506 2413 2509 2426
rect 2466 2303 2485 2306
rect 2482 2246 2485 2303
rect 2458 2203 2461 2246
rect 2482 2243 2489 2246
rect 2486 2196 2489 2243
rect 2498 2213 2501 2336
rect 2514 2333 2517 2446
rect 2506 2303 2509 2326
rect 2522 2256 2525 2336
rect 2546 2333 2549 2566
rect 2558 2563 2565 2566
rect 2558 2506 2561 2563
rect 2558 2503 2565 2506
rect 2562 2486 2565 2503
rect 2562 2483 2573 2486
rect 2570 2336 2573 2483
rect 2586 2426 2589 2526
rect 2598 2436 2601 2573
rect 2618 2556 2621 2696
rect 2626 2616 2629 2713
rect 2634 2623 2637 2736
rect 2642 2713 2645 2726
rect 2650 2696 2653 2926
rect 2658 2803 2661 2836
rect 2666 2786 2669 3243
rect 2682 3223 2685 3463
rect 2706 3406 2709 3483
rect 2706 3403 2717 3406
rect 2722 3403 2725 3526
rect 2730 3413 2733 3486
rect 2754 3476 2757 3573
rect 2770 3556 2773 3746
rect 2802 3733 2805 3806
rect 2818 3743 2821 3936
rect 2834 3826 2837 4126
rect 2842 3933 2845 4006
rect 2866 3926 2869 4016
rect 2874 4003 2877 4126
rect 2914 4103 2917 4126
rect 2922 4026 2925 4136
rect 2938 4133 2941 4166
rect 2962 4116 2965 4176
rect 2954 4113 2965 4116
rect 2954 4036 2957 4113
rect 2954 4033 2961 4036
rect 2914 4023 2925 4026
rect 2874 3933 2877 3946
rect 2850 3923 2869 3926
rect 2834 3823 2845 3826
rect 2826 3686 2829 3806
rect 2842 3803 2845 3823
rect 2850 3813 2853 3916
rect 2858 3913 2869 3916
rect 2882 3913 2885 4016
rect 2890 3993 2893 4006
rect 2914 3956 2917 4023
rect 2914 3953 2925 3956
rect 2922 3933 2925 3953
rect 2938 3926 2941 4016
rect 2946 3933 2949 3996
rect 2958 3956 2961 4033
rect 2958 3953 2965 3956
rect 2922 3923 2941 3926
rect 2858 3793 2861 3913
rect 2938 3906 2941 3923
rect 2954 3916 2957 3936
rect 2930 3903 2941 3906
rect 2950 3913 2957 3916
rect 2930 3836 2933 3903
rect 2950 3836 2953 3913
rect 2930 3833 2941 3836
rect 2950 3833 2957 3836
rect 2866 3813 2869 3826
rect 2914 3813 2933 3816
rect 2874 3736 2877 3806
rect 2906 3766 2909 3806
rect 2922 3793 2925 3806
rect 2906 3763 2925 3766
rect 2870 3733 2877 3736
rect 2818 3683 2829 3686
rect 2818 3653 2821 3683
rect 2834 3636 2837 3726
rect 2870 3646 2873 3733
rect 2870 3643 2877 3646
rect 2826 3633 2837 3636
rect 2766 3553 2773 3556
rect 2766 3496 2769 3553
rect 2766 3493 2773 3496
rect 2754 3473 2765 3476
rect 2762 3456 2765 3473
rect 2770 3463 2773 3493
rect 2778 3483 2781 3576
rect 2826 3556 2829 3633
rect 2842 3596 2845 3626
rect 2866 3613 2869 3626
rect 2842 3593 2853 3596
rect 2826 3553 2837 3556
rect 2786 3533 2789 3546
rect 2834 3533 2837 3553
rect 2850 3546 2853 3593
rect 2842 3543 2853 3546
rect 2874 3546 2877 3643
rect 2882 3603 2885 3726
rect 2898 3696 2901 3756
rect 2922 3723 2925 3763
rect 2894 3693 2901 3696
rect 2894 3626 2897 3693
rect 2906 3636 2909 3656
rect 2906 3633 2917 3636
rect 2894 3623 2901 3626
rect 2874 3543 2885 3546
rect 2818 3503 2821 3526
rect 2842 3523 2845 3543
rect 2874 3516 2877 3536
rect 2754 3453 2765 3456
rect 2714 3383 2717 3403
rect 2738 3383 2741 3406
rect 2730 3323 2733 3346
rect 2770 3313 2773 3336
rect 2778 3323 2781 3406
rect 2690 3203 2693 3216
rect 2738 3206 2741 3286
rect 2722 3133 2725 3206
rect 2730 3203 2741 3206
rect 2730 3123 2733 3203
rect 2738 3133 2741 3146
rect 2746 3123 2749 3136
rect 2754 3133 2757 3186
rect 2786 3146 2789 3356
rect 2794 3323 2797 3416
rect 2818 3413 2821 3426
rect 2810 3333 2813 3406
rect 2834 3396 2837 3506
rect 2842 3496 2845 3516
rect 2866 3513 2877 3516
rect 2842 3493 2853 3496
rect 2850 3436 2853 3493
rect 2842 3433 2853 3436
rect 2866 3436 2869 3513
rect 2866 3433 2877 3436
rect 2842 3403 2845 3433
rect 2850 3413 2869 3416
rect 2834 3393 2845 3396
rect 2818 3333 2821 3346
rect 2778 3143 2789 3146
rect 2778 3076 2781 3143
rect 2802 3116 2805 3136
rect 2810 3123 2813 3326
rect 2818 3323 2829 3326
rect 2834 3256 2837 3386
rect 2842 3313 2845 3393
rect 2858 3383 2861 3406
rect 2874 3403 2877 3433
rect 2882 3363 2885 3543
rect 2898 3536 2901 3623
rect 2914 3576 2917 3633
rect 2938 3613 2941 3833
rect 2954 3813 2957 3833
rect 2946 3606 2949 3736
rect 2962 3703 2965 3953
rect 2970 3653 2973 4186
rect 2986 4133 2989 4276
rect 3026 4223 3029 4353
rect 3058 4346 3061 4416
rect 3074 4376 3077 4446
rect 3122 4443 3125 4536
rect 3130 4523 3133 4543
rect 3138 4503 3141 4536
rect 3074 4373 3085 4376
rect 3054 4343 3061 4346
rect 3042 4193 3045 4326
rect 3054 4296 3057 4343
rect 3054 4293 3061 4296
rect 3058 4273 3061 4293
rect 3050 4203 3053 4226
rect 3066 4213 3069 4336
rect 2978 4113 2981 4126
rect 2994 4103 2997 4126
rect 2978 4023 2989 4026
rect 2978 3913 2981 4023
rect 2994 3913 2997 4016
rect 2890 3533 2901 3536
rect 2906 3573 2917 3576
rect 2938 3603 2949 3606
rect 2890 3353 2893 3533
rect 2898 3403 2901 3526
rect 2906 3396 2909 3573
rect 2930 3513 2933 3526
rect 2914 3413 2917 3506
rect 2938 3496 2941 3603
rect 2954 3556 2957 3646
rect 2962 3613 2965 3626
rect 2970 3613 2973 3636
rect 2934 3493 2941 3496
rect 2946 3553 2957 3556
rect 2830 3253 2837 3256
rect 2818 3133 2821 3216
rect 2830 3166 2833 3253
rect 2850 3166 2853 3336
rect 2890 3333 2893 3346
rect 2898 3323 2901 3396
rect 2906 3393 2917 3396
rect 2922 3393 2925 3416
rect 2906 3333 2909 3386
rect 2914 3376 2917 3393
rect 2914 3373 2925 3376
rect 2922 3326 2925 3373
rect 2914 3323 2925 3326
rect 2874 3206 2877 3256
rect 2914 3226 2917 3323
rect 2934 3276 2937 3493
rect 2946 3286 2949 3553
rect 2962 3546 2965 3606
rect 2978 3556 2981 3816
rect 2986 3623 2989 3736
rect 2994 3723 2997 3806
rect 3002 3736 3005 4136
rect 3042 4133 3045 4146
rect 3010 4096 3013 4126
rect 3050 4123 3053 4136
rect 3010 4093 3021 4096
rect 3018 4036 3021 4093
rect 3010 4033 3021 4036
rect 3010 3936 3013 4033
rect 3018 4003 3021 4016
rect 3034 4006 3037 4106
rect 3042 4023 3053 4026
rect 3026 3973 3029 4006
rect 3034 4003 3041 4006
rect 3010 3933 3021 3936
rect 3010 3893 3013 3926
rect 3018 3813 3021 3933
rect 3026 3913 3029 3926
rect 3038 3916 3041 4003
rect 3058 3953 3061 4206
rect 3066 4106 3069 4156
rect 3074 4143 3077 4236
rect 3082 4123 3085 4373
rect 3090 4333 3093 4416
rect 3090 4223 3093 4326
rect 3098 4273 3101 4336
rect 3114 4323 3117 4436
rect 3138 4403 3141 4486
rect 3146 4433 3149 4526
rect 3154 4523 3157 4616
rect 3178 4566 3181 4606
rect 3174 4563 3181 4566
rect 3162 4523 3165 4546
rect 3154 4333 3157 4506
rect 3174 4476 3177 4563
rect 3186 4486 3189 4576
rect 3194 4543 3213 4546
rect 3194 4533 3197 4543
rect 3202 4503 3205 4536
rect 3210 4523 3213 4543
rect 3218 4533 3221 4576
rect 3186 4483 3197 4486
rect 3174 4473 3181 4476
rect 3162 4413 3165 4466
rect 3178 4396 3181 4473
rect 3194 4426 3197 4483
rect 3186 4423 3197 4426
rect 3186 4403 3189 4423
rect 3218 4413 3221 4476
rect 3178 4393 3189 4396
rect 3154 4323 3165 4326
rect 3130 4236 3133 4256
rect 3170 4253 3173 4336
rect 3178 4323 3181 4346
rect 3186 4316 3189 4393
rect 3210 4346 3213 4406
rect 3234 4403 3237 4426
rect 3242 4416 3245 4526
rect 3250 4483 3253 4606
rect 3266 4513 3269 4536
rect 3274 4523 3277 4616
rect 3282 4523 3285 4536
rect 3290 4523 3293 4546
rect 3314 4506 3317 4536
rect 3322 4513 3325 4526
rect 3242 4413 3253 4416
rect 3210 4343 3221 4346
rect 3210 4323 3213 4336
rect 3178 4313 3189 4316
rect 3130 4233 3141 4236
rect 3138 4176 3141 4233
rect 3154 4213 3157 4226
rect 3178 4203 3181 4313
rect 3218 4226 3221 4343
rect 3242 4333 3245 4406
rect 3250 4306 3253 4413
rect 3258 4396 3261 4416
rect 3266 4403 3269 4506
rect 3306 4503 3317 4506
rect 3274 4413 3277 4496
rect 3306 4436 3309 4503
rect 3306 4433 3317 4436
rect 3274 4396 3277 4406
rect 3258 4393 3277 4396
rect 3258 4333 3261 4386
rect 3282 4376 3285 4416
rect 3298 4403 3301 4416
rect 3266 4373 3285 4376
rect 3266 4323 3269 4373
rect 3242 4303 3253 4306
rect 3194 4213 3197 4226
rect 3218 4223 3229 4226
rect 3130 4173 3141 4176
rect 3066 4103 3077 4106
rect 3074 3936 3077 4103
rect 3050 3923 3053 3936
rect 3034 3913 3041 3916
rect 3010 3803 3021 3806
rect 3002 3733 3021 3736
rect 3002 3626 3005 3716
rect 3010 3643 3013 3726
rect 3018 3706 3021 3733
rect 3026 3713 3029 3806
rect 3034 3733 3037 3913
rect 3058 3903 3061 3936
rect 3066 3933 3077 3936
rect 3042 3876 3045 3896
rect 3042 3873 3053 3876
rect 3050 3756 3053 3873
rect 3066 3816 3069 3933
rect 3082 3893 3085 3916
rect 3062 3813 3069 3816
rect 3062 3766 3065 3813
rect 3074 3773 3077 3806
rect 3082 3786 3085 3816
rect 3090 3796 3093 4136
rect 3106 4083 3109 4126
rect 3098 4003 3101 4026
rect 3114 4013 3117 4076
rect 3130 4036 3133 4173
rect 3138 4123 3141 4136
rect 3122 4033 3133 4036
rect 3106 3933 3109 3976
rect 3114 3903 3117 3926
rect 3122 3886 3125 4033
rect 3130 4013 3133 4026
rect 3138 4003 3141 4016
rect 3146 4003 3149 4126
rect 3154 3956 3157 4006
rect 3170 4003 3173 4046
rect 3178 4043 3205 4046
rect 3178 4033 3181 4043
rect 3186 4003 3189 4016
rect 3150 3953 3157 3956
rect 3118 3883 3125 3886
rect 3118 3816 3121 3883
rect 3118 3813 3125 3816
rect 3090 3793 3101 3796
rect 3122 3793 3125 3813
rect 3130 3796 3133 3936
rect 3150 3896 3153 3953
rect 3150 3893 3157 3896
rect 3154 3873 3157 3893
rect 3138 3813 3141 3836
rect 3162 3803 3165 3946
rect 3194 3933 3197 4036
rect 3202 4023 3205 4043
rect 3202 4003 3205 4016
rect 3210 3933 3213 4216
rect 3226 4156 3229 4223
rect 3242 4213 3245 4303
rect 3290 4263 3293 4336
rect 3242 4196 3245 4206
rect 3250 4203 3253 4236
rect 3258 4196 3261 4216
rect 3242 4193 3261 4196
rect 3218 4153 3229 4156
rect 3218 4096 3221 4153
rect 3226 4113 3229 4126
rect 3218 4093 3225 4096
rect 3222 3946 3225 4093
rect 3218 3943 3225 3946
rect 3170 3913 3173 3926
rect 3210 3913 3213 3926
rect 3130 3793 3137 3796
rect 3082 3783 3093 3786
rect 3062 3763 3069 3766
rect 3042 3753 3053 3756
rect 3018 3703 3025 3706
rect 3022 3646 3025 3703
rect 3022 3643 3029 3646
rect 3002 3623 3009 3626
rect 2994 3603 2997 3616
rect 3006 3556 3009 3623
rect 3018 3613 3021 3626
rect 2978 3553 2997 3556
rect 2954 3543 2965 3546
rect 2954 3433 2957 3543
rect 2978 3533 2981 3546
rect 2994 3506 2997 3553
rect 2978 3503 2997 3506
rect 3002 3553 3009 3556
rect 2962 3323 2965 3406
rect 2970 3403 2973 3426
rect 2946 3283 2957 3286
rect 2934 3273 2941 3276
rect 2914 3223 2925 3226
rect 2874 3203 2885 3206
rect 2830 3163 2837 3166
rect 2834 3133 2837 3163
rect 2846 3163 2853 3166
rect 2826 3123 2837 3126
rect 2774 3073 2781 3076
rect 2798 3113 2805 3116
rect 2698 3003 2701 3026
rect 2682 2893 2685 2966
rect 2698 2933 2701 2996
rect 2722 2993 2725 3016
rect 2706 2923 2709 2936
rect 2714 2923 2717 2936
rect 2674 2836 2677 2856
rect 2674 2833 2681 2836
rect 2662 2783 2669 2786
rect 2662 2716 2665 2783
rect 2678 2776 2681 2833
rect 2690 2813 2693 2826
rect 2706 2813 2725 2816
rect 2674 2773 2681 2776
rect 2662 2713 2669 2716
rect 2646 2693 2653 2696
rect 2666 2693 2669 2713
rect 2646 2626 2649 2693
rect 2674 2686 2677 2773
rect 2690 2733 2693 2806
rect 2698 2766 2701 2806
rect 2714 2793 2717 2806
rect 2738 2766 2741 2926
rect 2698 2763 2717 2766
rect 2714 2723 2717 2763
rect 2730 2763 2741 2766
rect 2762 2763 2765 3036
rect 2774 2956 2777 3073
rect 2798 3036 2801 3113
rect 2846 3106 2849 3163
rect 2842 3103 2849 3106
rect 2798 3033 2805 3036
rect 2770 2953 2777 2956
rect 2770 2933 2773 2953
rect 2778 2923 2781 2936
rect 2786 2933 2789 3016
rect 2794 2963 2797 3016
rect 2802 2846 2805 3033
rect 2810 3013 2813 3086
rect 2818 2973 2821 3006
rect 2842 2966 2845 3103
rect 2842 2963 2853 2966
rect 2834 2933 2837 2946
rect 2850 2916 2853 2963
rect 2794 2843 2805 2846
rect 2842 2913 2853 2916
rect 2842 2846 2845 2913
rect 2842 2843 2853 2846
rect 2658 2683 2677 2686
rect 2646 2623 2653 2626
rect 2626 2613 2637 2616
rect 2626 2593 2629 2606
rect 2618 2553 2629 2556
rect 2598 2433 2605 2436
rect 2582 2423 2589 2426
rect 2582 2356 2585 2423
rect 2582 2353 2589 2356
rect 2570 2333 2577 2336
rect 2530 2313 2533 2326
rect 2522 2253 2533 2256
rect 2482 2193 2489 2196
rect 2442 2143 2461 2146
rect 2434 2103 2441 2106
rect 2438 2046 2441 2103
rect 2434 2043 2441 2046
rect 2434 2026 2437 2043
rect 2426 2023 2437 2026
rect 2426 1946 2429 2023
rect 2442 1953 2445 2016
rect 2426 1943 2437 1946
rect 2426 1913 2429 1926
rect 2410 1813 2413 1826
rect 2334 1703 2341 1706
rect 2318 1623 2325 1626
rect 2318 1576 2321 1623
rect 2318 1573 2325 1576
rect 2322 1553 2325 1573
rect 2330 1536 2333 1616
rect 2314 1533 2333 1536
rect 2294 1513 2301 1516
rect 2294 1406 2297 1513
rect 2314 1506 2317 1526
rect 2306 1503 2317 1506
rect 2306 1413 2309 1503
rect 2294 1403 2301 1406
rect 2234 1313 2241 1316
rect 2202 1263 2221 1266
rect 2170 1243 2181 1246
rect 2170 1213 2173 1243
rect 2158 1203 2165 1206
rect 2162 966 2165 1203
rect 2186 1156 2189 1206
rect 2178 1153 2189 1156
rect 2178 1103 2181 1153
rect 2186 1013 2189 1146
rect 2194 1056 2197 1176
rect 2218 1173 2221 1263
rect 2234 1236 2237 1313
rect 2226 1233 2237 1236
rect 2226 1156 2229 1233
rect 2234 1213 2237 1226
rect 2250 1166 2253 1316
rect 2266 1256 2269 1333
rect 2282 1303 2285 1326
rect 2290 1303 2293 1326
rect 2298 1313 2301 1403
rect 2306 1273 2309 1336
rect 2314 1283 2317 1416
rect 2338 1363 2341 1703
rect 2354 1603 2357 1656
rect 2386 1626 2389 1716
rect 2394 1703 2397 1726
rect 2402 1713 2405 1786
rect 2418 1766 2421 1816
rect 2414 1763 2421 1766
rect 2414 1666 2417 1763
rect 2414 1663 2421 1666
rect 2386 1623 2397 1626
rect 2354 1413 2357 1436
rect 2362 1396 2365 1536
rect 2378 1533 2381 1616
rect 2394 1546 2397 1623
rect 2418 1583 2421 1663
rect 2426 1603 2429 1756
rect 2386 1543 2397 1546
rect 2386 1523 2389 1543
rect 2410 1516 2413 1556
rect 2418 1533 2421 1546
rect 2426 1526 2429 1536
rect 2434 1526 2437 1943
rect 2442 1753 2445 1816
rect 2450 1803 2453 2136
rect 2458 2096 2461 2143
rect 2482 2113 2485 2193
rect 2530 2176 2533 2253
rect 2554 2213 2557 2306
rect 2562 2213 2565 2326
rect 2574 2226 2577 2333
rect 2586 2316 2589 2353
rect 2594 2323 2597 2416
rect 2602 2353 2605 2433
rect 2610 2423 2613 2526
rect 2602 2333 2613 2336
rect 2618 2333 2621 2546
rect 2626 2413 2629 2553
rect 2634 2543 2637 2613
rect 2642 2526 2645 2596
rect 2650 2553 2653 2623
rect 2638 2523 2645 2526
rect 2638 2376 2641 2523
rect 2650 2383 2653 2506
rect 2658 2396 2661 2683
rect 2698 2613 2701 2626
rect 2674 2523 2677 2606
rect 2666 2403 2669 2506
rect 2674 2413 2677 2516
rect 2698 2503 2701 2526
rect 2658 2393 2669 2396
rect 2638 2373 2645 2376
rect 2586 2313 2597 2316
rect 2610 2313 2613 2326
rect 2570 2223 2577 2226
rect 2570 2196 2573 2223
rect 2526 2173 2533 2176
rect 2562 2193 2573 2196
rect 2514 2113 2517 2126
rect 2498 2103 2509 2106
rect 2458 2093 2469 2096
rect 2466 2036 2469 2093
rect 2514 2063 2517 2106
rect 2526 2036 2529 2173
rect 2546 2116 2549 2136
rect 2546 2113 2553 2116
rect 2458 2033 2469 2036
rect 2522 2033 2529 2036
rect 2458 2013 2461 2033
rect 2482 1936 2485 1956
rect 2498 1953 2501 2016
rect 2478 1933 2485 1936
rect 2506 1933 2509 2006
rect 2514 1933 2517 2016
rect 2522 2013 2525 2033
rect 2530 1943 2533 2016
rect 2538 2003 2541 2096
rect 2466 1813 2469 1926
rect 2478 1886 2481 1933
rect 2490 1896 2493 1916
rect 2490 1893 2501 1896
rect 2478 1883 2485 1886
rect 2450 1653 2453 1796
rect 2474 1616 2477 1816
rect 2482 1703 2485 1883
rect 2498 1776 2501 1893
rect 2514 1843 2517 1926
rect 2530 1826 2533 1926
rect 2538 1913 2541 1956
rect 2550 1946 2553 2113
rect 2546 1943 2553 1946
rect 2546 1923 2549 1943
rect 2562 1923 2565 2193
rect 2578 2143 2581 2206
rect 2594 2203 2597 2313
rect 2626 2213 2629 2336
rect 2634 2313 2637 2326
rect 2642 2256 2645 2373
rect 2638 2253 2645 2256
rect 2638 2176 2641 2253
rect 2638 2173 2645 2176
rect 2578 2133 2589 2136
rect 2570 2083 2573 2126
rect 2514 1823 2533 1826
rect 2514 1813 2517 1823
rect 2522 1803 2525 1816
rect 2490 1773 2501 1776
rect 2442 1533 2445 1616
rect 2458 1613 2477 1616
rect 2490 1613 2493 1773
rect 2498 1676 2501 1726
rect 2514 1723 2533 1726
rect 2498 1673 2505 1676
rect 2450 1553 2453 1606
rect 2426 1523 2437 1526
rect 2450 1523 2453 1536
rect 2410 1513 2421 1516
rect 2418 1436 2421 1513
rect 2418 1433 2429 1436
rect 2358 1393 2365 1396
rect 2322 1333 2325 1346
rect 2222 1153 2229 1156
rect 2246 1163 2253 1166
rect 2258 1253 2269 1256
rect 2202 1076 2205 1126
rect 2210 1093 2213 1136
rect 2202 1073 2213 1076
rect 2194 1053 2201 1056
rect 2162 963 2169 966
rect 2074 896 2077 936
rect 2098 923 2101 936
rect 2122 923 2125 946
rect 2074 893 2085 896
rect 2082 826 2085 893
rect 2074 823 2085 826
rect 2074 796 2077 823
rect 2106 806 2109 876
rect 2050 713 2053 796
rect 2058 793 2077 796
rect 2082 723 2085 806
rect 2090 773 2093 806
rect 2102 803 2109 806
rect 2090 706 2093 756
rect 2102 746 2105 803
rect 2102 743 2109 746
rect 2082 703 2093 706
rect 2058 613 2061 676
rect 2066 613 2069 626
rect 2042 423 2045 536
rect 2050 526 2053 606
rect 2058 533 2061 576
rect 2082 546 2085 703
rect 2098 613 2101 726
rect 2106 573 2109 743
rect 2114 673 2117 796
rect 2122 756 2125 916
rect 2130 773 2133 796
rect 2122 753 2129 756
rect 2126 686 2129 753
rect 2122 683 2129 686
rect 2122 666 2125 683
rect 2114 663 2125 666
rect 2114 566 2117 663
rect 2098 563 2117 566
rect 2066 533 2069 546
rect 2082 543 2093 546
rect 2050 523 2069 526
rect 2090 523 2093 543
rect 2042 413 2053 416
rect 2058 413 2061 446
rect 2098 433 2101 563
rect 2114 533 2117 556
rect 2138 546 2141 956
rect 2166 896 2169 963
rect 2178 923 2181 1006
rect 2162 893 2169 896
rect 2162 873 2165 893
rect 2146 733 2149 816
rect 2154 806 2157 816
rect 2154 803 2173 806
rect 2162 723 2165 736
rect 2170 733 2173 803
rect 2186 753 2189 986
rect 2198 976 2201 1053
rect 2194 973 2201 976
rect 2194 793 2197 973
rect 2210 956 2213 1073
rect 2202 953 2213 956
rect 2202 933 2205 953
rect 2222 936 2225 1153
rect 2234 1123 2237 1146
rect 2222 933 2229 936
rect 2146 696 2149 716
rect 2178 706 2181 736
rect 2202 733 2205 916
rect 2226 913 2229 933
rect 2234 863 2237 1116
rect 2246 1106 2249 1163
rect 2258 1113 2261 1253
rect 2266 1213 2269 1236
rect 2298 1226 2301 1246
rect 2338 1236 2341 1326
rect 2346 1323 2349 1336
rect 2358 1326 2361 1393
rect 2370 1336 2373 1406
rect 2378 1363 2381 1416
rect 2386 1403 2389 1416
rect 2410 1383 2413 1396
rect 2370 1333 2377 1336
rect 2410 1333 2413 1366
rect 2418 1343 2421 1416
rect 2426 1396 2429 1433
rect 2434 1413 2437 1523
rect 2458 1506 2461 1613
rect 2450 1503 2461 1506
rect 2450 1436 2453 1503
rect 2450 1433 2461 1436
rect 2466 1433 2469 1606
rect 2474 1523 2477 1536
rect 2482 1533 2485 1606
rect 2490 1593 2493 1606
rect 2502 1586 2505 1673
rect 2514 1603 2517 1723
rect 2482 1503 2485 1526
rect 2442 1403 2445 1416
rect 2426 1393 2433 1396
rect 2450 1393 2453 1406
rect 2458 1403 2461 1433
rect 2466 1413 2469 1426
rect 2430 1336 2433 1393
rect 2442 1343 2445 1356
rect 2426 1333 2433 1336
rect 2358 1323 2365 1326
rect 2362 1243 2365 1323
rect 2374 1276 2377 1333
rect 2370 1273 2377 1276
rect 2274 1213 2277 1226
rect 2294 1223 2301 1226
rect 2294 1176 2297 1223
rect 2306 1183 2309 1206
rect 2294 1173 2301 1176
rect 2314 1173 2317 1236
rect 2330 1233 2341 1236
rect 2322 1213 2325 1226
rect 2330 1216 2333 1233
rect 2338 1223 2357 1226
rect 2330 1213 2341 1216
rect 2338 1203 2341 1213
rect 2266 1106 2269 1126
rect 2246 1103 2253 1106
rect 2266 1103 2277 1106
rect 2242 923 2245 1006
rect 2250 953 2253 1103
rect 2274 1056 2277 1103
rect 2298 1076 2301 1173
rect 2338 1106 2341 1126
rect 2330 1103 2341 1106
rect 2298 1073 2309 1076
rect 2266 1053 2277 1056
rect 2258 906 2261 1026
rect 2266 1003 2269 1053
rect 2266 926 2269 936
rect 2282 933 2285 1036
rect 2298 1003 2301 1016
rect 2306 966 2309 1073
rect 2330 1036 2333 1103
rect 2330 1033 2341 1036
rect 2298 963 2309 966
rect 2322 966 2325 1016
rect 2338 1003 2341 1033
rect 2346 983 2349 1216
rect 2354 1013 2357 1223
rect 2362 1213 2365 1236
rect 2370 1203 2373 1273
rect 2378 1156 2381 1216
rect 2386 1213 2389 1326
rect 2394 1213 2397 1246
rect 2402 1203 2405 1256
rect 2426 1233 2429 1333
rect 2410 1223 2421 1226
rect 2410 1203 2413 1216
rect 2418 1163 2421 1223
rect 2426 1213 2429 1226
rect 2442 1216 2445 1236
rect 2450 1226 2453 1316
rect 2450 1223 2461 1226
rect 2466 1223 2469 1406
rect 2474 1233 2477 1326
rect 2482 1226 2485 1416
rect 2490 1243 2493 1586
rect 2502 1583 2509 1586
rect 2530 1583 2533 1706
rect 2506 1516 2509 1583
rect 2530 1533 2533 1546
rect 2538 1516 2541 1846
rect 2570 1843 2573 2076
rect 2578 2066 2581 2133
rect 2642 2126 2645 2173
rect 2586 2076 2589 2126
rect 2634 2123 2645 2126
rect 2602 2096 2605 2116
rect 2602 2093 2613 2096
rect 2586 2073 2597 2076
rect 2578 2063 2589 2066
rect 2578 1953 2581 2026
rect 2586 1936 2589 2063
rect 2594 2023 2597 2073
rect 2610 2036 2613 2093
rect 2634 2073 2637 2123
rect 2642 2103 2645 2116
rect 2650 2113 2653 2126
rect 2666 2113 2669 2393
rect 2682 2373 2685 2416
rect 2690 2353 2693 2426
rect 2674 2316 2677 2336
rect 2674 2313 2685 2316
rect 2682 2236 2685 2313
rect 2674 2233 2685 2236
rect 2674 2213 2677 2233
rect 2706 2213 2709 2696
rect 2730 2686 2733 2763
rect 2770 2723 2773 2806
rect 2730 2683 2741 2686
rect 2738 2593 2741 2683
rect 2778 2613 2781 2716
rect 2794 2666 2797 2843
rect 2810 2813 2813 2836
rect 2818 2813 2821 2826
rect 2834 2813 2837 2826
rect 2810 2703 2813 2806
rect 2826 2803 2837 2806
rect 2818 2723 2821 2796
rect 2842 2793 2845 2806
rect 2850 2773 2853 2843
rect 2842 2716 2845 2766
rect 2842 2713 2853 2716
rect 2810 2676 2813 2696
rect 2842 2686 2845 2706
rect 2834 2683 2845 2686
rect 2810 2673 2821 2676
rect 2794 2663 2805 2666
rect 2802 2646 2805 2663
rect 2802 2643 2809 2646
rect 2786 2603 2789 2616
rect 2786 2533 2789 2546
rect 2722 2403 2725 2426
rect 2730 2413 2741 2416
rect 2738 2373 2741 2406
rect 2754 2403 2757 2526
rect 2778 2513 2781 2526
rect 2794 2516 2797 2626
rect 2806 2566 2809 2643
rect 2790 2513 2797 2516
rect 2802 2563 2809 2566
rect 2778 2413 2781 2426
rect 2790 2416 2793 2513
rect 2790 2413 2797 2416
rect 2730 2196 2733 2316
rect 2746 2206 2749 2276
rect 2754 2213 2757 2386
rect 2786 2376 2789 2396
rect 2782 2373 2789 2376
rect 2762 2336 2765 2356
rect 2762 2333 2773 2336
rect 2770 2266 2773 2333
rect 2762 2263 2773 2266
rect 2762 2213 2765 2263
rect 2714 2193 2733 2196
rect 2738 2193 2741 2206
rect 2746 2203 2757 2206
rect 2770 2196 2773 2246
rect 2782 2236 2785 2373
rect 2754 2193 2773 2196
rect 2778 2233 2785 2236
rect 2674 2106 2677 2116
rect 2690 2113 2693 2126
rect 2658 2103 2677 2106
rect 2682 2046 2685 2106
rect 2714 2096 2717 2193
rect 2754 2133 2757 2193
rect 2738 2103 2741 2116
rect 2714 2093 2733 2096
rect 2730 2056 2733 2093
rect 2730 2053 2741 2056
rect 2682 2043 2693 2046
rect 2602 2033 2613 2036
rect 2602 2016 2605 2033
rect 2594 2013 2613 2016
rect 2690 2013 2693 2043
rect 2626 2003 2653 2006
rect 2582 1933 2589 1936
rect 2582 1866 2585 1933
rect 2578 1863 2585 1866
rect 2578 1813 2581 1863
rect 2554 1743 2557 1806
rect 2586 1796 2589 1846
rect 2570 1793 2589 1796
rect 2546 1706 2549 1726
rect 2546 1703 2553 1706
rect 2550 1626 2553 1703
rect 2498 1513 2509 1516
rect 2534 1513 2541 1516
rect 2546 1623 2553 1626
rect 2498 1493 2501 1513
rect 2534 1436 2537 1513
rect 2534 1433 2541 1436
rect 2498 1333 2501 1416
rect 2474 1223 2485 1226
rect 2442 1213 2453 1216
rect 2434 1193 2437 1206
rect 2442 1173 2445 1206
rect 2378 1153 2385 1156
rect 2370 1103 2373 1146
rect 2382 1106 2385 1153
rect 2418 1133 2421 1146
rect 2394 1113 2397 1126
rect 2378 1103 2385 1106
rect 2378 1083 2381 1103
rect 2402 1076 2405 1096
rect 2402 1073 2409 1076
rect 2394 1036 2397 1056
rect 2386 1033 2397 1036
rect 2386 966 2389 1033
rect 2406 1026 2409 1073
rect 2402 1023 2409 1026
rect 2402 976 2405 1023
rect 2402 973 2409 976
rect 2322 963 2333 966
rect 2386 963 2397 966
rect 2266 923 2285 926
rect 2258 903 2281 906
rect 2278 846 2281 903
rect 2298 886 2301 963
rect 2298 883 2313 886
rect 2210 813 2213 826
rect 2170 703 2181 706
rect 2186 723 2205 726
rect 2146 693 2157 696
rect 2154 636 2157 693
rect 2170 646 2173 703
rect 2170 643 2181 646
rect 2146 633 2157 636
rect 2146 613 2149 633
rect 2178 623 2181 643
rect 2186 636 2189 723
rect 2202 643 2205 716
rect 2218 636 2221 736
rect 2186 633 2205 636
rect 2186 616 2189 633
rect 2178 613 2189 616
rect 2138 543 2145 546
rect 2142 496 2145 543
rect 2138 493 2145 496
rect 2130 413 2133 436
rect 2138 413 2141 493
rect 2146 413 2149 426
rect 2154 416 2157 606
rect 2194 603 2197 616
rect 2202 613 2205 633
rect 2214 633 2221 636
rect 2202 586 2205 606
rect 2194 583 2205 586
rect 2162 523 2165 546
rect 2194 476 2197 583
rect 2214 556 2217 633
rect 2214 553 2221 556
rect 2194 473 2205 476
rect 2154 413 2165 416
rect 2170 413 2173 436
rect 2050 393 2053 406
rect 2050 366 2053 386
rect 2098 383 2101 406
rect 2050 363 2061 366
rect 2058 306 2061 363
rect 2106 333 2109 406
rect 2138 333 2141 406
rect 2050 303 2061 306
rect 2050 213 2053 303
rect 2114 213 2117 236
rect 2154 213 2157 336
rect 2162 323 2165 413
rect 2170 323 2173 406
rect 2178 403 2181 456
rect 2194 393 2197 406
rect 2202 383 2205 473
rect 2178 216 2181 376
rect 2210 363 2213 536
rect 2218 373 2221 553
rect 2226 526 2229 626
rect 2234 573 2237 846
rect 2278 843 2285 846
rect 2250 813 2269 816
rect 2250 783 2253 806
rect 2266 803 2269 813
rect 2266 753 2269 796
rect 2242 613 2245 626
rect 2258 623 2261 716
rect 2258 593 2261 616
rect 2266 586 2269 616
rect 2274 603 2277 826
rect 2282 733 2285 843
rect 2290 733 2293 856
rect 2310 826 2313 883
rect 2330 846 2333 963
rect 2346 913 2349 926
rect 2322 843 2333 846
rect 2370 843 2373 936
rect 2386 913 2389 926
rect 2298 813 2301 826
rect 2310 823 2317 826
rect 2290 706 2293 726
rect 2306 723 2309 806
rect 2314 716 2317 823
rect 2322 786 2325 843
rect 2338 823 2365 826
rect 2338 803 2341 823
rect 2346 813 2357 816
rect 2362 813 2365 823
rect 2354 796 2357 806
rect 2362 803 2373 806
rect 2378 796 2381 826
rect 2354 793 2381 796
rect 2322 783 2341 786
rect 2338 766 2341 783
rect 2286 703 2293 706
rect 2298 713 2317 716
rect 2330 763 2341 766
rect 2286 606 2289 703
rect 2298 613 2301 713
rect 2286 603 2293 606
rect 2258 583 2269 586
rect 2234 533 2245 536
rect 2250 533 2253 546
rect 2226 523 2245 526
rect 2226 366 2229 436
rect 2258 433 2261 583
rect 2274 526 2277 536
rect 2270 523 2277 526
rect 2270 466 2273 523
rect 2282 493 2285 526
rect 2290 513 2293 603
rect 2306 593 2309 696
rect 2330 666 2333 763
rect 2370 693 2373 786
rect 2394 783 2397 963
rect 2406 906 2409 973
rect 2418 926 2421 1106
rect 2434 1043 2437 1136
rect 2450 1103 2453 1213
rect 2450 1046 2453 1076
rect 2458 1053 2461 1223
rect 2466 1183 2469 1216
rect 2450 1043 2461 1046
rect 2442 1013 2445 1026
rect 2458 1013 2461 1043
rect 2466 1013 2469 1116
rect 2426 943 2445 946
rect 2426 933 2429 943
rect 2418 923 2429 926
rect 2434 923 2437 936
rect 2442 923 2445 943
rect 2406 903 2413 906
rect 2410 826 2413 903
rect 2402 823 2413 826
rect 2378 713 2381 726
rect 2330 663 2341 666
rect 2314 616 2317 626
rect 2322 616 2325 646
rect 2314 613 2325 616
rect 2314 523 2317 613
rect 2322 563 2325 606
rect 2266 463 2273 466
rect 2266 416 2269 463
rect 2330 423 2333 606
rect 2338 533 2341 663
rect 2346 616 2349 666
rect 2354 616 2357 626
rect 2346 613 2357 616
rect 2346 513 2349 613
rect 2354 593 2357 606
rect 2362 603 2365 656
rect 2402 653 2405 823
rect 2426 813 2429 923
rect 2418 763 2421 806
rect 2442 776 2445 816
rect 2450 803 2453 1006
rect 2474 1003 2477 1223
rect 2482 1183 2485 1206
rect 2466 803 2469 836
rect 2426 773 2445 776
rect 2426 733 2429 773
rect 2418 713 2421 726
rect 2426 696 2429 726
rect 2422 693 2429 696
rect 2402 616 2405 626
rect 2410 623 2413 666
rect 2422 616 2425 693
rect 2434 623 2437 736
rect 2474 733 2477 916
rect 2482 906 2485 1166
rect 2490 1113 2493 1216
rect 2506 1206 2509 1426
rect 2538 1413 2541 1433
rect 2514 1343 2533 1346
rect 2514 1323 2517 1343
rect 2522 1323 2525 1336
rect 2530 1333 2533 1343
rect 2530 1283 2533 1326
rect 2538 1266 2541 1346
rect 2546 1306 2549 1623
rect 2554 1533 2557 1606
rect 2562 1543 2565 1736
rect 2570 1723 2573 1793
rect 2586 1623 2589 1716
rect 2586 1523 2589 1616
rect 2594 1506 2597 1956
rect 2602 1933 2605 1986
rect 2602 1563 2605 1926
rect 2618 1743 2621 1956
rect 2586 1503 2597 1506
rect 2586 1446 2589 1503
rect 2586 1443 2597 1446
rect 2602 1443 2605 1516
rect 2610 1503 2613 1716
rect 2618 1713 2621 1726
rect 2618 1586 2621 1616
rect 2626 1603 2629 1886
rect 2634 1813 2637 1826
rect 2642 1813 2645 1916
rect 2650 1906 2653 2003
rect 2666 1953 2669 2006
rect 2738 1976 2741 2053
rect 2754 1993 2757 2006
rect 2730 1973 2741 1976
rect 2714 1913 2717 1926
rect 2650 1903 2661 1906
rect 2658 1846 2661 1903
rect 2650 1843 2661 1846
rect 2634 1696 2637 1806
rect 2650 1753 2653 1843
rect 2658 1783 2661 1816
rect 2666 1793 2669 1826
rect 2682 1813 2693 1816
rect 2698 1813 2717 1816
rect 2706 1793 2709 1806
rect 2714 1783 2717 1806
rect 2730 1803 2733 1973
rect 2754 1893 2757 1936
rect 2762 1933 2765 2016
rect 2770 1876 2773 2046
rect 2754 1873 2773 1876
rect 2650 1733 2653 1746
rect 2634 1693 2641 1696
rect 2674 1693 2677 1726
rect 2618 1583 2629 1586
rect 2618 1523 2621 1536
rect 2626 1456 2629 1583
rect 2638 1536 2641 1693
rect 2618 1453 2629 1456
rect 2634 1533 2641 1536
rect 2554 1323 2557 1416
rect 2546 1303 2553 1306
rect 2502 1203 2509 1206
rect 2534 1263 2541 1266
rect 2502 1156 2505 1203
rect 2514 1166 2517 1196
rect 2514 1163 2525 1166
rect 2502 1153 2509 1156
rect 2506 1136 2509 1153
rect 2506 1133 2513 1136
rect 2490 1003 2493 1026
rect 2490 923 2493 956
rect 2498 933 2501 1126
rect 2510 1056 2513 1133
rect 2506 1053 2513 1056
rect 2482 903 2493 906
rect 2490 836 2493 903
rect 2482 833 2493 836
rect 2442 723 2461 726
rect 2482 723 2485 833
rect 2490 763 2493 816
rect 2498 793 2501 806
rect 2370 613 2381 616
rect 2386 613 2405 616
rect 2378 586 2381 606
rect 2374 583 2381 586
rect 2218 363 2229 366
rect 2186 323 2205 326
rect 2210 306 2213 336
rect 2202 303 2213 306
rect 2202 256 2205 303
rect 2202 253 2213 256
rect 2210 233 2213 253
rect 2026 133 2029 166
rect 2066 163 2069 206
rect 2146 203 2157 206
rect 2162 203 2165 216
rect 2178 213 2197 216
rect 2034 133 2037 146
rect 2090 133 2093 166
rect 2018 123 2037 126
rect 2138 123 2141 136
rect 2170 133 2173 206
rect 2186 183 2189 206
rect 2194 133 2197 206
rect 2210 203 2213 216
rect 2218 213 2221 363
rect 2226 333 2229 356
rect 2226 306 2229 326
rect 2234 323 2237 386
rect 2250 333 2253 416
rect 2262 413 2269 416
rect 2262 316 2265 413
rect 2282 393 2285 416
rect 2258 313 2265 316
rect 2226 303 2237 306
rect 2234 236 2237 303
rect 2226 233 2237 236
rect 2258 236 2261 313
rect 2258 233 2269 236
rect 2210 123 2213 196
rect 2226 183 2229 233
rect 2266 216 2269 233
rect 2234 203 2237 216
rect 2258 213 2277 216
rect 2250 123 2253 206
rect 2266 183 2269 206
rect 2274 193 2277 206
rect 2282 196 2285 346
rect 2330 343 2333 416
rect 2346 413 2349 426
rect 2362 413 2365 536
rect 2374 516 2377 583
rect 2386 526 2389 576
rect 2386 523 2397 526
rect 2402 523 2405 613
rect 2418 613 2425 616
rect 2442 613 2445 723
rect 2458 663 2461 716
rect 2506 703 2509 1053
rect 2522 1036 2525 1163
rect 2534 1126 2537 1263
rect 2550 1256 2553 1303
rect 2546 1253 2553 1256
rect 2534 1123 2541 1126
rect 2514 1033 2525 1036
rect 2538 1036 2541 1123
rect 2546 1116 2549 1253
rect 2554 1123 2557 1216
rect 2578 1186 2581 1406
rect 2594 1296 2597 1443
rect 2634 1423 2637 1533
rect 2610 1393 2613 1406
rect 2602 1313 2605 1336
rect 2626 1323 2629 1336
rect 2634 1323 2637 1416
rect 2642 1386 2645 1516
rect 2650 1403 2653 1686
rect 2674 1623 2677 1646
rect 2682 1633 2685 1716
rect 2690 1623 2701 1626
rect 2690 1576 2693 1616
rect 2690 1573 2701 1576
rect 2658 1523 2661 1536
rect 2690 1516 2693 1536
rect 2698 1533 2701 1573
rect 2682 1513 2693 1516
rect 2682 1466 2685 1513
rect 2682 1463 2693 1466
rect 2642 1383 2649 1386
rect 2646 1326 2649 1383
rect 2642 1323 2649 1326
rect 2642 1306 2645 1323
rect 2634 1303 2645 1306
rect 2594 1293 2605 1296
rect 2578 1183 2589 1186
rect 2562 1143 2565 1166
rect 2578 1156 2581 1176
rect 2574 1153 2581 1156
rect 2546 1113 2565 1116
rect 2538 1033 2549 1036
rect 2514 923 2517 1033
rect 2530 933 2533 1016
rect 2538 903 2541 936
rect 2546 896 2549 1033
rect 2562 923 2565 1113
rect 2574 976 2577 1153
rect 2586 1053 2589 1183
rect 2602 1146 2605 1293
rect 2634 1196 2637 1303
rect 2658 1226 2661 1446
rect 2690 1333 2693 1463
rect 2698 1413 2701 1526
rect 2706 1493 2709 1506
rect 2714 1416 2717 1756
rect 2722 1703 2725 1746
rect 2730 1723 2733 1786
rect 2754 1756 2757 1873
rect 2778 1823 2781 2233
rect 2794 2216 2797 2413
rect 2802 2393 2805 2563
rect 2818 2546 2821 2673
rect 2810 2543 2821 2546
rect 2834 2546 2837 2683
rect 2834 2543 2845 2546
rect 2810 2516 2813 2543
rect 2818 2523 2837 2526
rect 2810 2513 2821 2516
rect 2818 2456 2821 2513
rect 2842 2506 2845 2543
rect 2838 2503 2845 2506
rect 2818 2453 2829 2456
rect 2786 2213 2797 2216
rect 2786 2106 2789 2213
rect 2794 2123 2797 2206
rect 2802 2143 2805 2216
rect 2810 2203 2813 2376
rect 2826 2206 2829 2453
rect 2838 2396 2841 2503
rect 2850 2473 2853 2713
rect 2858 2676 2861 3196
rect 2882 3156 2885 3203
rect 2874 3153 2885 3156
rect 2866 2723 2869 3016
rect 2874 3006 2877 3153
rect 2882 3103 2885 3136
rect 2890 3033 2893 3126
rect 2906 3123 2909 3146
rect 2914 3123 2917 3216
rect 2874 3003 2893 3006
rect 2874 2976 2877 2996
rect 2874 2973 2881 2976
rect 2878 2836 2881 2973
rect 2874 2833 2881 2836
rect 2874 2693 2877 2833
rect 2882 2803 2885 2816
rect 2882 2713 2885 2736
rect 2890 2676 2893 3003
rect 2898 2933 2901 3006
rect 2906 2973 2909 3026
rect 2914 2943 2917 3096
rect 2898 2813 2901 2846
rect 2906 2833 2909 2936
rect 2914 2903 2917 2916
rect 2922 2856 2925 3223
rect 2938 3206 2941 3273
rect 2938 3203 2945 3206
rect 2930 3113 2933 3196
rect 2942 3106 2945 3203
rect 2954 3193 2957 3283
rect 2970 3206 2973 3236
rect 2966 3203 2973 3206
rect 2966 3146 2969 3203
rect 2966 3143 2973 3146
rect 2970 3126 2973 3143
rect 2954 3123 2973 3126
rect 2938 3103 2945 3106
rect 2930 2963 2933 3036
rect 2930 2923 2933 2946
rect 2918 2853 2925 2856
rect 2918 2806 2921 2853
rect 2930 2813 2933 2846
rect 2918 2803 2925 2806
rect 2914 2733 2917 2756
rect 2858 2673 2869 2676
rect 2866 2556 2869 2673
rect 2858 2553 2869 2556
rect 2882 2673 2893 2676
rect 2882 2556 2885 2673
rect 2882 2553 2893 2556
rect 2858 2426 2861 2553
rect 2866 2513 2869 2526
rect 2874 2503 2877 2536
rect 2882 2513 2885 2536
rect 2890 2496 2893 2553
rect 2886 2493 2893 2496
rect 2850 2423 2861 2426
rect 2850 2406 2853 2423
rect 2858 2413 2869 2416
rect 2850 2403 2861 2406
rect 2838 2393 2845 2396
rect 2818 2203 2829 2206
rect 2786 2103 2797 2106
rect 2794 2036 2797 2103
rect 2790 2033 2797 2036
rect 2790 1946 2793 2033
rect 2786 1943 2793 1946
rect 2786 1896 2789 1943
rect 2802 1936 2805 2016
rect 2818 2013 2821 2203
rect 2842 2156 2845 2393
rect 2850 2313 2853 2326
rect 2858 2313 2861 2403
rect 2874 2336 2877 2456
rect 2886 2346 2889 2493
rect 2898 2453 2901 2726
rect 2914 2426 2917 2716
rect 2922 2706 2925 2803
rect 2930 2723 2933 2736
rect 2922 2703 2929 2706
rect 2926 2476 2929 2703
rect 2898 2423 2917 2426
rect 2922 2473 2929 2476
rect 2886 2343 2893 2346
rect 2870 2333 2877 2336
rect 2870 2246 2873 2333
rect 2870 2243 2877 2246
rect 2866 2203 2869 2226
rect 2842 2153 2861 2156
rect 2834 2106 2837 2126
rect 2830 2103 2837 2106
rect 2830 2026 2833 2103
rect 2830 2023 2837 2026
rect 2834 2003 2837 2023
rect 2842 2013 2845 2146
rect 2850 2103 2853 2126
rect 2858 2106 2861 2153
rect 2874 2123 2877 2243
rect 2882 2213 2885 2326
rect 2890 2196 2893 2343
rect 2898 2223 2901 2423
rect 2914 2333 2917 2416
rect 2906 2213 2909 2316
rect 2890 2193 2901 2196
rect 2898 2116 2901 2193
rect 2922 2146 2925 2473
rect 2930 2423 2933 2456
rect 2930 2333 2933 2416
rect 2938 2386 2941 3103
rect 2946 3013 2949 3056
rect 2946 2833 2949 2966
rect 2954 2943 2957 3016
rect 2962 2926 2965 3046
rect 2970 3023 2973 3036
rect 2958 2923 2965 2926
rect 2946 2803 2949 2826
rect 2958 2786 2961 2923
rect 2970 2793 2973 2966
rect 2958 2783 2965 2786
rect 2962 2626 2965 2783
rect 2978 2776 2981 3503
rect 2994 3413 2997 3426
rect 2986 3116 2989 3196
rect 3002 3186 3005 3553
rect 3010 3516 3013 3536
rect 3010 3513 3017 3516
rect 3014 3426 3017 3513
rect 3010 3423 3017 3426
rect 3010 3403 3013 3423
rect 3010 3323 3013 3346
rect 3026 3286 3029 3643
rect 3034 3603 3037 3716
rect 3042 3613 3045 3753
rect 3066 3743 3069 3763
rect 3058 3713 3061 3736
rect 3066 3733 3077 3736
rect 3090 3733 3093 3783
rect 3098 3763 3101 3793
rect 3122 3746 3125 3766
rect 3118 3743 3125 3746
rect 3042 3573 3045 3606
rect 3034 3413 3037 3426
rect 3050 3413 3053 3616
rect 3074 3613 3077 3626
rect 3082 3533 3085 3696
rect 3090 3583 3093 3726
rect 3098 3723 3101 3736
rect 3058 3523 3077 3526
rect 3050 3333 3053 3356
rect 3074 3346 3077 3516
rect 3082 3403 3085 3526
rect 3090 3503 3093 3536
rect 3098 3493 3101 3616
rect 3106 3576 3109 3736
rect 3118 3626 3121 3743
rect 3134 3736 3137 3793
rect 3130 3733 3137 3736
rect 3130 3676 3133 3733
rect 3130 3673 3141 3676
rect 3118 3623 3125 3626
rect 3114 3593 3117 3606
rect 3106 3573 3113 3576
rect 3110 3486 3113 3573
rect 3106 3483 3113 3486
rect 3090 3393 3093 3406
rect 3074 3343 3081 3346
rect 3050 3296 3053 3326
rect 3050 3293 3057 3296
rect 3026 3283 3045 3286
rect 3010 3203 3013 3226
rect 3026 3213 3029 3256
rect 3002 3183 3013 3186
rect 2986 3113 2997 3116
rect 2994 3046 2997 3113
rect 2986 3043 2997 3046
rect 2986 2853 2989 3043
rect 2974 2773 2981 2776
rect 2974 2636 2977 2773
rect 2974 2633 2981 2636
rect 2954 2623 2965 2626
rect 2954 2496 2957 2623
rect 2970 2596 2973 2616
rect 2966 2593 2973 2596
rect 2966 2516 2969 2593
rect 2978 2526 2981 2633
rect 2986 2613 2989 2816
rect 2978 2523 2985 2526
rect 2966 2513 2973 2516
rect 2954 2493 2965 2496
rect 2946 2403 2949 2446
rect 2938 2383 2945 2386
rect 2942 2326 2945 2383
rect 2938 2323 2945 2326
rect 2938 2276 2941 2323
rect 2954 2293 2957 2476
rect 2934 2273 2941 2276
rect 2934 2156 2937 2273
rect 2934 2153 2941 2156
rect 2890 2113 2901 2116
rect 2914 2143 2925 2146
rect 2858 2103 2869 2106
rect 2866 2036 2869 2103
rect 2890 2096 2893 2113
rect 2858 2033 2869 2036
rect 2882 2093 2893 2096
rect 2882 2036 2885 2093
rect 2882 2033 2893 2036
rect 2802 1933 2821 1936
rect 2794 1913 2797 1926
rect 2786 1893 2793 1896
rect 2778 1793 2781 1816
rect 2790 1786 2793 1893
rect 2802 1803 2805 1933
rect 2786 1783 2793 1786
rect 2754 1753 2773 1756
rect 2730 1713 2741 1716
rect 2738 1693 2741 1706
rect 2746 1676 2749 1726
rect 2738 1673 2749 1676
rect 2730 1646 2733 1666
rect 2726 1643 2733 1646
rect 2726 1546 2729 1643
rect 2726 1543 2733 1546
rect 2730 1523 2733 1543
rect 2738 1513 2741 1673
rect 2746 1623 2749 1636
rect 2754 1633 2757 1706
rect 2762 1703 2765 1716
rect 2746 1523 2749 1536
rect 2754 1503 2757 1626
rect 2762 1613 2765 1626
rect 2770 1596 2773 1753
rect 2786 1736 2789 1783
rect 2766 1593 2773 1596
rect 2778 1733 2789 1736
rect 2714 1413 2725 1416
rect 2666 1293 2669 1326
rect 2682 1313 2685 1326
rect 2698 1303 2701 1326
rect 2706 1263 2709 1406
rect 2722 1366 2725 1413
rect 2738 1403 2741 1416
rect 2714 1363 2725 1366
rect 2714 1276 2717 1363
rect 2754 1346 2757 1406
rect 2766 1366 2769 1593
rect 2766 1363 2773 1366
rect 2754 1343 2761 1346
rect 2730 1323 2733 1336
rect 2758 1296 2761 1343
rect 2754 1293 2761 1296
rect 2754 1276 2757 1293
rect 2714 1273 2725 1276
rect 2654 1223 2661 1226
rect 2634 1193 2645 1196
rect 2642 1173 2645 1193
rect 2594 1143 2605 1146
rect 2626 1143 2645 1146
rect 2594 1086 2597 1143
rect 2626 1133 2629 1143
rect 2602 1103 2605 1126
rect 2634 1113 2637 1136
rect 2642 1123 2645 1143
rect 2594 1083 2605 1086
rect 2602 976 2605 1083
rect 2654 1066 2657 1223
rect 2654 1063 2661 1066
rect 2618 1013 2621 1026
rect 2642 1003 2645 1056
rect 2658 1043 2661 1063
rect 2658 1013 2661 1026
rect 2574 973 2581 976
rect 2538 893 2549 896
rect 2522 746 2525 826
rect 2538 813 2541 893
rect 2514 743 2525 746
rect 2450 613 2453 626
rect 2410 533 2413 606
rect 2418 603 2421 613
rect 2374 513 2381 516
rect 2378 453 2381 513
rect 2354 336 2357 406
rect 2306 323 2309 336
rect 2354 333 2365 336
rect 2394 333 2397 523
rect 2402 413 2405 456
rect 2418 446 2421 576
rect 2442 573 2445 606
rect 2450 583 2453 606
rect 2490 586 2493 606
rect 2482 583 2493 586
rect 2414 443 2421 446
rect 2414 396 2417 443
rect 2414 393 2421 396
rect 2442 393 2445 556
rect 2482 516 2485 583
rect 2498 523 2501 616
rect 2506 593 2509 606
rect 2514 603 2517 743
rect 2522 733 2541 736
rect 2530 546 2533 726
rect 2538 723 2541 733
rect 2538 703 2541 716
rect 2554 686 2557 736
rect 2562 713 2565 826
rect 2570 803 2573 936
rect 2578 916 2581 973
rect 2594 973 2605 976
rect 2578 913 2589 916
rect 2578 893 2581 906
rect 2586 876 2589 913
rect 2582 873 2589 876
rect 2582 816 2585 873
rect 2578 813 2585 816
rect 2578 803 2581 813
rect 2594 756 2597 973
rect 2602 943 2621 946
rect 2602 923 2605 943
rect 2610 923 2613 936
rect 2618 933 2621 943
rect 2642 933 2645 946
rect 2602 893 2605 916
rect 2618 893 2621 926
rect 2610 783 2613 806
rect 2626 803 2629 906
rect 2586 753 2597 756
rect 2586 733 2589 753
rect 2602 723 2605 736
rect 2546 683 2557 686
rect 2546 636 2549 683
rect 2546 633 2557 636
rect 2522 543 2533 546
rect 2482 513 2493 516
rect 2490 413 2493 513
rect 2522 466 2525 543
rect 2546 516 2549 536
rect 2542 513 2549 516
rect 2522 463 2533 466
rect 2530 433 2533 463
rect 2542 436 2545 513
rect 2542 433 2549 436
rect 2546 413 2549 433
rect 2466 393 2469 406
rect 2418 346 2421 393
rect 2490 353 2509 356
rect 2418 343 2429 346
rect 2362 323 2365 333
rect 2426 296 2429 343
rect 2442 313 2445 326
rect 2418 293 2429 296
rect 2418 216 2421 293
rect 2474 276 2477 326
rect 2482 313 2485 326
rect 2474 273 2485 276
rect 2490 273 2493 353
rect 2498 333 2501 346
rect 2506 333 2509 353
rect 2514 343 2517 356
rect 2498 323 2517 326
rect 2282 193 2293 196
rect 2290 176 2293 193
rect 2306 176 2309 206
rect 2354 193 2357 216
rect 2418 213 2437 216
rect 2426 183 2429 206
rect 2442 193 2445 206
rect 2290 173 2309 176
rect 2290 133 2293 173
rect 2330 133 2333 166
rect 2450 146 2453 216
rect 2378 113 2381 126
rect 2418 123 2421 146
rect 2434 143 2453 146
rect 2426 73 2429 136
rect 2434 123 2437 143
rect 2442 113 2445 136
rect 2458 133 2461 186
rect 2474 156 2477 206
rect 2482 203 2485 273
rect 2498 213 2501 256
rect 2514 203 2517 323
rect 2530 246 2533 396
rect 2554 346 2557 633
rect 2562 613 2565 686
rect 2562 523 2565 606
rect 2602 603 2605 716
rect 2634 706 2637 726
rect 2630 703 2637 706
rect 2630 626 2633 703
rect 2630 623 2637 626
rect 2610 603 2613 616
rect 2554 343 2561 346
rect 2558 296 2561 343
rect 2526 243 2533 246
rect 2554 293 2561 296
rect 2526 196 2529 243
rect 2538 223 2541 236
rect 2554 213 2557 293
rect 2570 273 2573 536
rect 2586 523 2589 566
rect 2610 516 2613 536
rect 2602 513 2613 516
rect 2602 466 2605 513
rect 2618 506 2621 616
rect 2634 603 2637 623
rect 2642 613 2645 786
rect 2650 596 2653 986
rect 2658 813 2661 926
rect 2666 906 2669 1216
rect 2674 1106 2677 1136
rect 2682 1123 2685 1236
rect 2698 1213 2701 1246
rect 2722 1186 2725 1273
rect 2746 1273 2757 1276
rect 2746 1226 2749 1273
rect 2770 1266 2773 1363
rect 2778 1343 2781 1733
rect 2786 1613 2789 1726
rect 2810 1663 2813 1926
rect 2826 1923 2829 1996
rect 2842 1893 2845 1926
rect 2818 1813 2821 1826
rect 2834 1803 2837 1826
rect 2818 1783 2821 1796
rect 2834 1733 2837 1766
rect 2818 1723 2845 1726
rect 2810 1623 2813 1656
rect 2818 1613 2821 1723
rect 2850 1716 2853 1876
rect 2858 1813 2861 2033
rect 2866 1933 2869 1956
rect 2874 1923 2877 2016
rect 2882 1916 2885 2016
rect 2890 2013 2893 2033
rect 2890 1923 2893 1966
rect 2874 1913 2885 1916
rect 2834 1713 2853 1716
rect 2834 1696 2837 1713
rect 2830 1693 2837 1696
rect 2830 1556 2833 1693
rect 2858 1683 2861 1736
rect 2866 1703 2869 1856
rect 2874 1733 2877 1913
rect 2882 1813 2885 1836
rect 2890 1803 2893 1896
rect 2898 1796 2901 2066
rect 2914 2026 2917 2143
rect 2914 2023 2925 2026
rect 2930 2023 2933 2136
rect 2938 2096 2941 2153
rect 2946 2113 2949 2266
rect 2954 2203 2957 2246
rect 2962 2186 2965 2493
rect 2970 2213 2973 2513
rect 2982 2236 2985 2523
rect 2978 2233 2985 2236
rect 2958 2183 2965 2186
rect 2958 2116 2961 2183
rect 2970 2123 2973 2166
rect 2958 2113 2965 2116
rect 2938 2093 2949 2096
rect 2906 1993 2909 2006
rect 2906 1813 2909 1926
rect 2890 1793 2901 1796
rect 2890 1726 2893 1793
rect 2914 1736 2917 1896
rect 2922 1813 2925 2023
rect 2946 2016 2949 2093
rect 2938 2013 2949 2016
rect 2938 1936 2941 2013
rect 2962 1996 2965 2113
rect 2978 2106 2981 2233
rect 2974 2103 2981 2106
rect 2974 2006 2977 2103
rect 2986 2013 2989 2216
rect 2994 2166 2997 3026
rect 3010 2996 3013 3183
rect 3002 2993 3013 2996
rect 3034 2993 3037 3216
rect 3042 3193 3045 3283
rect 3054 3226 3057 3293
rect 3066 3283 3069 3336
rect 3078 3256 3081 3343
rect 3074 3253 3081 3256
rect 3074 3233 3077 3253
rect 3050 3223 3057 3226
rect 3050 3203 3053 3223
rect 3074 3213 3077 3226
rect 3042 3003 3045 3036
rect 3058 3023 3061 3206
rect 3074 3163 3077 3206
rect 3090 3123 3093 3326
rect 3098 3323 3101 3416
rect 3106 3256 3109 3483
rect 3114 3423 3117 3436
rect 3114 3323 3117 3416
rect 3122 3366 3125 3623
rect 3130 3603 3133 3666
rect 3138 3526 3141 3673
rect 3146 3603 3149 3726
rect 3130 3523 3141 3526
rect 3130 3386 3133 3523
rect 3138 3493 3141 3516
rect 3146 3513 3149 3526
rect 3154 3466 3157 3746
rect 3162 3716 3165 3796
rect 3178 3743 3181 3896
rect 3186 3736 3189 3876
rect 3194 3803 3197 3906
rect 3218 3893 3221 3943
rect 3226 3823 3229 3926
rect 3234 3873 3237 4086
rect 3242 4013 3245 4076
rect 3250 4033 3253 4146
rect 3266 4133 3269 4206
rect 3274 4176 3277 4216
rect 3298 4213 3301 4276
rect 3306 4203 3309 4416
rect 3314 4403 3317 4433
rect 3330 4423 3333 4616
rect 3338 4433 3341 4526
rect 3346 4506 3349 4526
rect 3346 4503 3357 4506
rect 3354 4456 3357 4503
rect 3346 4453 3357 4456
rect 3314 4293 3317 4356
rect 3314 4196 3317 4216
rect 3322 4203 3325 4336
rect 3330 4273 3333 4416
rect 3346 4413 3349 4453
rect 3362 4413 3365 4436
rect 3370 4413 3373 4606
rect 3386 4506 3389 4526
rect 3394 4523 3397 4616
rect 3402 4523 3405 4566
rect 3410 4543 3429 4546
rect 3410 4533 3413 4543
rect 3418 4523 3421 4536
rect 3426 4523 3429 4543
rect 3450 4533 3453 4616
rect 3474 4613 3493 4616
rect 3386 4503 3397 4506
rect 3394 4446 3397 4503
rect 3386 4443 3397 4446
rect 3442 4443 3445 4526
rect 3466 4473 3469 4526
rect 3386 4423 3389 4443
rect 3474 4436 3477 4536
rect 3490 4533 3493 4613
rect 3482 4463 3485 4526
rect 3474 4433 3493 4436
rect 3426 4413 3429 4426
rect 3338 4306 3341 4336
rect 3354 4333 3357 4406
rect 3474 4373 3477 4416
rect 3458 4333 3461 4366
rect 3474 4333 3477 4346
rect 3346 4323 3357 4326
rect 3338 4303 3345 4306
rect 3330 4213 3333 4256
rect 3330 4196 3333 4206
rect 3274 4173 3281 4176
rect 3266 4113 3269 4126
rect 3278 4106 3281 4173
rect 3274 4103 3281 4106
rect 3274 4033 3277 4103
rect 3242 3836 3245 4006
rect 3250 3946 3253 4006
rect 3258 3996 3261 4016
rect 3266 4003 3269 4016
rect 3274 3996 3277 4006
rect 3258 3993 3277 3996
rect 3282 3956 3285 4016
rect 3290 4013 3293 4126
rect 3298 4113 3301 4196
rect 3314 4193 3333 4196
rect 3342 4166 3345 4303
rect 3354 4296 3357 4323
rect 3362 4313 3365 4326
rect 3354 4293 3365 4296
rect 3362 4236 3365 4293
rect 3354 4233 3365 4236
rect 3354 4213 3357 4233
rect 3306 4143 3325 4146
rect 3306 4133 3309 4143
rect 3314 4103 3317 4136
rect 3322 4123 3325 4143
rect 3298 3983 3301 4086
rect 3330 4046 3333 4166
rect 3338 4163 3345 4166
rect 3338 4133 3341 4163
rect 3354 4133 3357 4146
rect 3338 4113 3341 4126
rect 3306 4043 3333 4046
rect 3274 3953 3285 3956
rect 3250 3943 3261 3946
rect 3234 3833 3245 3836
rect 3202 3743 3205 3816
rect 3234 3766 3237 3833
rect 3242 3803 3245 3826
rect 3226 3763 3237 3766
rect 3178 3733 3189 3736
rect 3162 3713 3169 3716
rect 3166 3656 3169 3713
rect 3162 3653 3169 3656
rect 3162 3593 3165 3653
rect 3178 3636 3181 3733
rect 3174 3633 3181 3636
rect 3174 3586 3177 3633
rect 3186 3593 3189 3616
rect 3170 3583 3177 3586
rect 3170 3516 3173 3583
rect 3178 3523 3181 3536
rect 3186 3533 3189 3546
rect 3170 3513 3181 3516
rect 3154 3463 3161 3466
rect 3138 3403 3141 3436
rect 3146 3413 3149 3456
rect 3158 3406 3161 3463
rect 3178 3456 3181 3513
rect 3178 3453 3185 3456
rect 3154 3403 3161 3406
rect 3130 3383 3141 3386
rect 3122 3363 3129 3366
rect 3126 3316 3129 3363
rect 3102 3253 3109 3256
rect 3122 3313 3129 3316
rect 3102 3146 3105 3253
rect 3102 3143 3109 3146
rect 3098 3083 3101 3126
rect 3106 3056 3109 3143
rect 3114 3123 3117 3246
rect 3102 3053 3109 3056
rect 3058 2993 3061 3006
rect 3002 2416 3005 2993
rect 3026 2936 3029 2976
rect 3010 2853 3013 2936
rect 3018 2933 3029 2936
rect 3074 2923 3077 2936
rect 3090 2923 3093 3016
rect 3102 2976 3105 3053
rect 3102 2973 3109 2976
rect 3082 2856 3085 2886
rect 3066 2853 3085 2856
rect 3010 2576 3013 2846
rect 3026 2813 3029 2836
rect 3042 2803 3045 2816
rect 3026 2746 3029 2786
rect 3026 2743 3045 2746
rect 3018 2716 3021 2736
rect 3018 2713 3029 2716
rect 3026 2656 3029 2713
rect 3018 2653 3029 2656
rect 3018 2596 3021 2653
rect 3042 2636 3045 2743
rect 3026 2633 3045 2636
rect 3026 2613 3029 2633
rect 3066 2626 3069 2853
rect 3098 2803 3101 2816
rect 3106 2736 3109 2973
rect 3122 2966 3125 3313
rect 3138 3266 3141 3383
rect 3154 3326 3157 3403
rect 3182 3376 3185 3453
rect 3178 3373 3185 3376
rect 3178 3336 3181 3373
rect 3178 3333 3185 3336
rect 3154 3323 3173 3326
rect 3130 3263 3141 3266
rect 3130 3243 3133 3263
rect 3130 3223 3133 3236
rect 3154 3233 3157 3316
rect 3138 3136 3141 3226
rect 3162 3216 3165 3256
rect 3158 3213 3165 3216
rect 3158 3146 3161 3213
rect 3130 3133 3141 3136
rect 3146 3133 3149 3146
rect 3158 3143 3165 3146
rect 3130 3093 3133 3133
rect 3154 3106 3157 3126
rect 3150 3103 3157 3106
rect 3130 3066 3133 3086
rect 3130 3063 3141 3066
rect 3138 2996 3141 3063
rect 3118 2963 3125 2966
rect 3130 2993 3141 2996
rect 3150 2996 3153 3103
rect 3150 2993 3157 2996
rect 3118 2796 3121 2963
rect 3130 2883 3133 2993
rect 3146 2803 3149 2976
rect 3154 2933 3157 2993
rect 3162 2986 3165 3143
rect 3170 3006 3173 3323
rect 3182 3266 3185 3333
rect 3178 3263 3185 3266
rect 3178 3223 3181 3263
rect 3178 3203 3181 3216
rect 3186 3203 3189 3246
rect 3178 3013 3181 3136
rect 3186 3133 3189 3146
rect 3186 3103 3189 3126
rect 3194 3086 3197 3606
rect 3202 3513 3205 3606
rect 3226 3583 3229 3763
rect 3250 3753 3253 3806
rect 3258 3763 3261 3943
rect 3274 3926 3277 3953
rect 3282 3943 3301 3946
rect 3282 3933 3285 3943
rect 3274 3923 3285 3926
rect 3266 3793 3269 3816
rect 3274 3783 3277 3806
rect 3266 3733 3269 3746
rect 3282 3726 3285 3923
rect 3290 3903 3293 3936
rect 3298 3923 3301 3943
rect 3306 3933 3309 4043
rect 3314 3936 3317 4036
rect 3322 4003 3325 4016
rect 3330 4013 3341 4016
rect 3346 3996 3349 4106
rect 3362 4003 3365 4016
rect 3342 3993 3349 3996
rect 3342 3936 3345 3993
rect 3314 3933 3333 3936
rect 3342 3933 3349 3936
rect 3290 3813 3293 3836
rect 3234 3523 3237 3616
rect 3242 3613 3245 3726
rect 3282 3723 3293 3726
rect 3282 3693 3285 3716
rect 3290 3686 3293 3723
rect 3274 3683 3293 3686
rect 3258 3626 3261 3646
rect 3254 3623 3261 3626
rect 3254 3536 3257 3623
rect 3266 3563 3269 3616
rect 3274 3613 3277 3683
rect 3274 3596 3277 3606
rect 3282 3603 3285 3626
rect 3290 3596 3293 3616
rect 3298 3603 3301 3766
rect 3306 3613 3309 3726
rect 3314 3643 3317 3926
rect 3330 3756 3333 3933
rect 3346 3916 3349 3933
rect 3354 3923 3357 3966
rect 3370 3963 3373 4066
rect 3386 4046 3389 4276
rect 3410 4213 3413 4326
rect 3426 4276 3429 4306
rect 3426 4273 3437 4276
rect 3434 4206 3437 4273
rect 3458 4236 3461 4326
rect 3474 4303 3477 4326
rect 3490 4323 3493 4433
rect 3498 4403 3501 4526
rect 3498 4324 3501 4356
rect 3426 4203 3437 4206
rect 3450 4233 3461 4236
rect 3402 4113 3405 4126
rect 3418 4046 3421 4146
rect 3382 4043 3389 4046
rect 3410 4043 3421 4046
rect 3382 3976 3385 4043
rect 3382 3973 3389 3976
rect 3386 3956 3389 3973
rect 3386 3953 3405 3956
rect 3370 3943 3389 3946
rect 3370 3923 3373 3943
rect 3346 3913 3357 3916
rect 3354 3836 3357 3913
rect 3378 3903 3381 3936
rect 3386 3933 3389 3943
rect 3386 3913 3389 3926
rect 3370 3856 3373 3876
rect 3370 3853 3381 3856
rect 3354 3833 3365 3836
rect 3338 3793 3341 3806
rect 3330 3753 3337 3756
rect 3314 3596 3317 3616
rect 3274 3593 3293 3596
rect 3298 3593 3317 3596
rect 3274 3566 3277 3586
rect 3274 3563 3281 3566
rect 3254 3533 3261 3536
rect 3202 3413 3205 3426
rect 3226 3403 3229 3466
rect 3242 3413 3245 3426
rect 3210 3233 3213 3336
rect 3210 3213 3213 3226
rect 3190 3083 3197 3086
rect 3170 3003 3181 3006
rect 3162 2983 3169 2986
rect 3166 2926 3169 2983
rect 3162 2923 3169 2926
rect 3118 2793 3125 2796
rect 3090 2693 3093 2736
rect 3106 2733 3113 2736
rect 3066 2623 3085 2626
rect 3018 2593 3029 2596
rect 3074 2593 3077 2606
rect 3010 2573 3017 2576
rect 3014 2466 3017 2573
rect 3010 2463 3017 2466
rect 3010 2423 3013 2463
rect 3026 2446 3029 2593
rect 3050 2523 3053 2536
rect 3058 2533 3061 2546
rect 3018 2443 3029 2446
rect 3002 2413 3013 2416
rect 3010 2326 3013 2413
rect 3018 2376 3021 2443
rect 3034 2403 3037 2416
rect 3074 2413 3077 2526
rect 3050 2393 3053 2406
rect 3018 2373 3037 2376
rect 3010 2323 3021 2326
rect 3002 2223 3005 2316
rect 3018 2276 3021 2323
rect 3010 2273 3021 2276
rect 2994 2163 3005 2166
rect 2974 2003 2981 2006
rect 2958 1993 2965 1996
rect 2958 1936 2961 1993
rect 2930 1933 2941 1936
rect 2930 1796 2933 1933
rect 2938 1903 2941 1926
rect 2946 1916 2949 1936
rect 2958 1933 2965 1936
rect 2970 1933 2973 1986
rect 2978 1933 2981 2003
rect 2946 1913 2957 1916
rect 2946 1853 2949 1906
rect 2938 1813 2941 1836
rect 2930 1793 2941 1796
rect 2930 1773 2933 1786
rect 2882 1723 2893 1726
rect 2842 1586 2845 1666
rect 2850 1613 2853 1626
rect 2842 1583 2849 1586
rect 2830 1553 2837 1556
rect 2786 1393 2789 1406
rect 2794 1396 2797 1516
rect 2802 1413 2805 1436
rect 2794 1393 2801 1396
rect 2778 1313 2781 1326
rect 2798 1296 2801 1393
rect 2794 1293 2801 1296
rect 2770 1263 2781 1266
rect 2746 1223 2757 1226
rect 2754 1203 2757 1223
rect 2762 1213 2765 1256
rect 2778 1216 2781 1263
rect 2770 1213 2781 1216
rect 2794 1213 2797 1293
rect 2802 1213 2805 1276
rect 2770 1193 2773 1213
rect 2810 1193 2813 1536
rect 2818 1523 2821 1536
rect 2826 1506 2829 1536
rect 2822 1503 2829 1506
rect 2822 1426 2825 1503
rect 2834 1446 2837 1553
rect 2846 1456 2849 1583
rect 2858 1523 2861 1636
rect 2874 1546 2877 1616
rect 2866 1543 2877 1546
rect 2846 1453 2853 1456
rect 2834 1443 2845 1446
rect 2822 1423 2829 1426
rect 2826 1403 2829 1423
rect 2842 1403 2845 1443
rect 2818 1313 2821 1326
rect 2842 1316 2845 1336
rect 2834 1313 2845 1316
rect 2818 1213 2821 1296
rect 2834 1236 2837 1313
rect 2834 1233 2845 1236
rect 2842 1216 2845 1233
rect 2834 1213 2845 1216
rect 2714 1183 2725 1186
rect 2714 1166 2717 1183
rect 2698 1163 2717 1166
rect 2674 1103 2681 1106
rect 2678 946 2681 1103
rect 2674 943 2681 946
rect 2674 923 2677 943
rect 2682 913 2685 926
rect 2666 903 2673 906
rect 2670 766 2673 903
rect 2690 856 2693 1046
rect 2698 983 2701 1163
rect 2714 1113 2717 1156
rect 2706 923 2709 1006
rect 2690 853 2697 856
rect 2694 806 2697 853
rect 2714 836 2717 936
rect 2722 933 2725 986
rect 2714 833 2721 836
rect 2706 813 2709 826
rect 2690 803 2697 806
rect 2670 763 2677 766
rect 2674 686 2677 763
rect 2690 713 2693 803
rect 2698 723 2701 786
rect 2718 776 2721 833
rect 2746 803 2749 1116
rect 2762 1113 2765 1126
rect 2794 1123 2797 1156
rect 2802 1113 2805 1126
rect 2818 1086 2821 1206
rect 2842 1193 2845 1206
rect 2842 1106 2845 1176
rect 2810 1083 2821 1086
rect 2834 1103 2845 1106
rect 2786 1023 2805 1026
rect 2786 953 2789 1023
rect 2770 923 2773 936
rect 2794 923 2797 1016
rect 2802 1013 2805 1023
rect 2802 996 2805 1006
rect 2810 1003 2813 1083
rect 2834 1046 2837 1103
rect 2834 1043 2845 1046
rect 2842 1023 2845 1043
rect 2818 996 2821 1016
rect 2850 1006 2853 1453
rect 2866 1423 2869 1543
rect 2874 1523 2877 1536
rect 2882 1506 2885 1723
rect 2906 1686 2909 1736
rect 2914 1733 2925 1736
rect 2898 1683 2909 1686
rect 2898 1576 2901 1683
rect 2914 1653 2917 1726
rect 2922 1716 2925 1733
rect 2922 1713 2929 1716
rect 2926 1576 2929 1713
rect 2898 1573 2909 1576
rect 2878 1503 2885 1506
rect 2878 1426 2881 1503
rect 2874 1423 2881 1426
rect 2874 1416 2877 1423
rect 2866 1413 2877 1416
rect 2866 1396 2869 1413
rect 2862 1393 2869 1396
rect 2862 1266 2865 1393
rect 2874 1276 2877 1406
rect 2882 1293 2885 1416
rect 2890 1403 2893 1536
rect 2898 1413 2901 1526
rect 2906 1513 2909 1573
rect 2922 1573 2929 1576
rect 2922 1436 2925 1573
rect 2938 1533 2941 1793
rect 2946 1763 2949 1816
rect 2954 1793 2957 1913
rect 2962 1803 2965 1933
rect 2986 1926 2989 1996
rect 2978 1923 2989 1926
rect 2970 1813 2973 1916
rect 2994 1913 2997 2006
rect 3002 1986 3005 2163
rect 3010 1993 3013 2273
rect 3034 2256 3037 2373
rect 3082 2366 3085 2623
rect 3098 2613 3101 2726
rect 3110 2606 3113 2733
rect 3090 2533 3093 2606
rect 3106 2603 3113 2606
rect 3106 2533 3109 2603
rect 3090 2483 3093 2526
rect 3122 2516 3125 2793
rect 3138 2706 3141 2726
rect 3134 2703 3141 2706
rect 3134 2636 3137 2703
rect 3134 2633 3141 2636
rect 3130 2563 3133 2616
rect 3138 2603 3141 2633
rect 3130 2523 3133 2546
rect 3074 2363 3085 2366
rect 3074 2266 3077 2363
rect 3090 2276 3093 2396
rect 3098 2326 3101 2516
rect 3122 2513 3133 2516
rect 3122 2476 3125 2496
rect 3118 2473 3125 2476
rect 3118 2356 3121 2473
rect 3118 2353 3125 2356
rect 3106 2333 3117 2336
rect 3098 2323 3109 2326
rect 3090 2273 3097 2276
rect 3074 2263 3085 2266
rect 3022 2253 3037 2256
rect 3022 2146 3025 2253
rect 3034 2203 3037 2226
rect 3050 2213 3053 2236
rect 3058 2223 3069 2226
rect 3074 2223 3077 2246
rect 3082 2206 3085 2263
rect 3042 2163 3045 2206
rect 3074 2203 3085 2206
rect 3018 2143 3025 2146
rect 3018 2006 3021 2143
rect 3026 2023 3029 2126
rect 3050 2096 3053 2146
rect 3074 2136 3077 2203
rect 3094 2196 3097 2273
rect 3090 2193 3097 2196
rect 3090 2143 3093 2193
rect 3074 2133 3085 2136
rect 3050 2093 3061 2096
rect 3058 2076 3061 2093
rect 3050 2073 3061 2076
rect 3050 2006 3053 2073
rect 3018 2003 3025 2006
rect 3050 2003 3061 2006
rect 3002 1983 3013 1986
rect 3002 1866 3005 1886
rect 2998 1863 3005 1866
rect 2986 1813 2989 1846
rect 2970 1773 2973 1806
rect 2946 1643 2949 1726
rect 2978 1716 2981 1796
rect 2998 1756 3001 1863
rect 3010 1813 3013 1983
rect 3022 1906 3025 2003
rect 3034 1913 3037 1926
rect 3058 1923 3061 2003
rect 3074 1966 3077 2096
rect 3082 2066 3085 2133
rect 3082 2063 3093 2066
rect 3090 2046 3093 2063
rect 3090 2043 3097 2046
rect 3094 1976 3097 2043
rect 3106 2013 3109 2323
rect 3114 2203 3117 2316
rect 3122 2233 3125 2353
rect 3130 2306 3133 2513
rect 3138 2413 3141 2536
rect 3146 2496 3149 2796
rect 3162 2733 3165 2923
rect 3178 2866 3181 3003
rect 3190 2886 3193 3083
rect 3202 2896 3205 3196
rect 3218 3136 3221 3296
rect 3242 3136 3245 3216
rect 3218 3133 3229 3136
rect 3210 3106 3213 3126
rect 3210 3103 3217 3106
rect 3214 3046 3217 3103
rect 3210 3043 3217 3046
rect 3210 3013 3213 3043
rect 3226 3026 3229 3133
rect 3238 3133 3245 3136
rect 3238 3036 3241 3133
rect 3250 3116 3253 3516
rect 3258 3476 3261 3533
rect 3278 3486 3281 3563
rect 3274 3483 3281 3486
rect 3258 3473 3265 3476
rect 3262 3376 3265 3473
rect 3258 3373 3265 3376
rect 3258 3353 3261 3373
rect 3258 3333 3261 3346
rect 3266 3313 3269 3336
rect 3258 3163 3261 3206
rect 3266 3183 3269 3206
rect 3274 3176 3277 3483
rect 3290 3466 3293 3566
rect 3298 3523 3301 3593
rect 3290 3463 3301 3466
rect 3322 3463 3325 3746
rect 3334 3626 3337 3753
rect 3346 3633 3349 3826
rect 3362 3776 3365 3833
rect 3358 3773 3365 3776
rect 3358 3636 3361 3773
rect 3378 3756 3381 3853
rect 3402 3776 3405 3953
rect 3410 3943 3413 4043
rect 3426 3996 3429 4203
rect 3450 4186 3453 4233
rect 3450 4183 3461 4186
rect 3434 4003 3437 4126
rect 3442 4113 3445 4126
rect 3458 4026 3461 4183
rect 3474 4143 3477 4206
rect 3482 4143 3501 4146
rect 3482 4133 3485 4143
rect 3482 4113 3485 4126
rect 3490 4103 3493 4136
rect 3498 4123 3501 4143
rect 3506 4086 3509 4556
rect 3514 4383 3517 4526
rect 3522 4516 3525 4566
rect 3530 4533 3533 4616
rect 3554 4593 3557 4606
rect 3570 4553 3573 4616
rect 3650 4613 3653 4636
rect 3682 4633 3685 4663
rect 3522 4513 3533 4516
rect 3546 4513 3549 4526
rect 3530 4436 3533 4513
rect 3554 4476 3557 4536
rect 3562 4486 3565 4546
rect 3578 4543 3581 4606
rect 3674 4583 3677 4606
rect 3690 4603 3693 4616
rect 3706 4606 3709 4673
rect 3762 4613 3765 4626
rect 3786 4623 3789 4740
rect 3818 4626 3821 4740
rect 3810 4623 3821 4626
rect 3698 4603 3709 4606
rect 3698 4586 3701 4603
rect 3682 4583 3701 4586
rect 3570 4523 3573 4536
rect 3594 4513 3597 4536
rect 3562 4483 3573 4486
rect 3554 4473 3565 4476
rect 3522 4433 3533 4436
rect 3522 4353 3525 4433
rect 3538 4396 3541 4416
rect 3546 4403 3549 4436
rect 3554 4413 3557 4446
rect 3554 4396 3557 4406
rect 3538 4393 3557 4396
rect 3514 4343 3533 4346
rect 3514 4323 3517 4343
rect 3522 4303 3525 4336
rect 3530 4333 3533 4343
rect 3538 4326 3541 4386
rect 3562 4343 3565 4473
rect 3570 4466 3573 4483
rect 3570 4463 3577 4466
rect 3574 4376 3577 4463
rect 3586 4413 3589 4426
rect 3594 4413 3597 4436
rect 3570 4373 3577 4376
rect 3530 4323 3541 4326
rect 3530 4253 3533 4323
rect 3546 4313 3549 4326
rect 3554 4303 3557 4326
rect 3562 4246 3565 4336
rect 3570 4286 3573 4373
rect 3586 4313 3589 4326
rect 3602 4313 3605 4526
rect 3682 4523 3685 4583
rect 3626 4413 3629 4426
rect 3610 4286 3613 4306
rect 3570 4283 3589 4286
rect 3562 4243 3573 4246
rect 3522 4213 3525 4236
rect 3554 4176 3557 4216
rect 3562 4213 3565 4236
rect 3570 4196 3573 4243
rect 3586 4226 3589 4283
rect 3546 4173 3557 4176
rect 3566 4193 3573 4196
rect 3578 4223 3589 4226
rect 3602 4283 3613 4286
rect 3602 4226 3605 4283
rect 3602 4223 3613 4226
rect 3498 4083 3509 4086
rect 3514 4083 3517 4136
rect 3530 4133 3533 4166
rect 3522 4113 3525 4126
rect 3458 4023 3465 4026
rect 3426 3993 3445 3996
rect 3426 3926 3429 3956
rect 3418 3923 3429 3926
rect 3418 3826 3421 3923
rect 3434 3906 3437 3936
rect 3442 3913 3445 3993
rect 3450 3933 3453 4016
rect 3462 3966 3465 4023
rect 3474 3973 3477 4026
rect 3482 3993 3485 4026
rect 3462 3963 3473 3966
rect 3450 3913 3453 3926
rect 3430 3903 3437 3906
rect 3430 3846 3433 3903
rect 3430 3843 3437 3846
rect 3418 3823 3429 3826
rect 3418 3783 3421 3806
rect 3402 3773 3421 3776
rect 3354 3633 3361 3636
rect 3370 3753 3381 3756
rect 3330 3623 3337 3626
rect 3330 3583 3333 3623
rect 3338 3576 3341 3606
rect 3338 3573 3345 3576
rect 3342 3506 3345 3573
rect 3354 3543 3357 3633
rect 3362 3603 3365 3616
rect 3338 3503 3345 3506
rect 3298 3356 3301 3463
rect 3306 3396 3309 3406
rect 3314 3403 3317 3456
rect 3338 3426 3341 3503
rect 3330 3423 3341 3426
rect 3346 3423 3349 3436
rect 3322 3396 3325 3416
rect 3306 3393 3325 3396
rect 3282 3333 3285 3346
rect 3290 3226 3293 3356
rect 3298 3353 3309 3356
rect 3298 3303 3301 3326
rect 3306 3323 3309 3353
rect 3322 3313 3325 3326
rect 3282 3213 3285 3226
rect 3290 3223 3305 3226
rect 3266 3173 3277 3176
rect 3266 3123 3269 3173
rect 3274 3116 3277 3136
rect 3282 3123 3285 3186
rect 3290 3133 3293 3216
rect 3302 3176 3305 3223
rect 3322 3213 3325 3226
rect 3302 3173 3309 3176
rect 3290 3116 3293 3126
rect 3250 3113 3269 3116
rect 3274 3113 3293 3116
rect 3238 3033 3245 3036
rect 3218 3023 3229 3026
rect 3202 2893 3209 2896
rect 3190 2883 3197 2886
rect 3178 2863 3185 2866
rect 3170 2823 3173 2856
rect 3182 2816 3185 2863
rect 3178 2813 3185 2816
rect 3178 2793 3181 2813
rect 3154 2713 3157 2726
rect 3162 2723 3173 2726
rect 3154 2613 3157 2686
rect 3154 2513 3157 2596
rect 3146 2493 3153 2496
rect 3150 2406 3153 2493
rect 3146 2403 3153 2406
rect 3138 2323 3141 2336
rect 3130 2303 3137 2306
rect 3134 2236 3137 2303
rect 3130 2233 3137 2236
rect 3130 2216 3133 2233
rect 3146 2216 3149 2403
rect 3154 2346 3157 2386
rect 3162 2366 3165 2706
rect 3170 2623 3173 2696
rect 3170 2586 3173 2616
rect 3178 2603 3181 2646
rect 3194 2613 3197 2883
rect 3206 2846 3209 2893
rect 3202 2843 3209 2846
rect 3202 2813 3205 2843
rect 3218 2826 3221 3023
rect 3242 3006 3245 3033
rect 3234 3003 3245 3006
rect 3234 2986 3237 3003
rect 3230 2983 3237 2986
rect 3230 2836 3233 2983
rect 3230 2833 3237 2836
rect 3210 2823 3221 2826
rect 3202 2713 3205 2726
rect 3210 2703 3213 2823
rect 3234 2816 3237 2833
rect 3218 2813 3237 2816
rect 3194 2593 3197 2606
rect 3170 2583 3189 2586
rect 3170 2513 3173 2566
rect 3186 2526 3189 2583
rect 3202 2533 3205 2546
rect 3186 2523 3197 2526
rect 3170 2383 3173 2456
rect 3186 2413 3189 2426
rect 3194 2396 3197 2523
rect 3218 2493 3221 2806
rect 3234 2773 3237 2813
rect 3226 2586 3229 2676
rect 3242 2636 3245 2996
rect 3250 2923 3253 3106
rect 3258 3023 3261 3036
rect 3266 2956 3269 3113
rect 3258 2953 3269 2956
rect 3258 2803 3261 2953
rect 3266 2916 3269 2936
rect 3282 2933 3285 3016
rect 3290 2976 3293 3113
rect 3298 3103 3301 3126
rect 3298 2983 3301 3006
rect 3290 2973 3301 2976
rect 3290 2923 3293 2946
rect 3298 2933 3301 2973
rect 3266 2913 3277 2916
rect 3274 2836 3277 2913
rect 3298 2846 3301 2926
rect 3306 2863 3309 3173
rect 3314 3073 3317 3126
rect 3330 3023 3333 3423
rect 3354 3246 3357 3536
rect 3362 3413 3365 3586
rect 3370 3396 3373 3753
rect 3378 3733 3389 3736
rect 3378 3583 3381 3676
rect 3394 3673 3397 3726
rect 3410 3723 3413 3736
rect 3386 3596 3389 3606
rect 3394 3603 3397 3616
rect 3402 3596 3405 3616
rect 3386 3593 3405 3596
rect 3410 3593 3413 3606
rect 3410 3566 3413 3586
rect 3418 3573 3421 3773
rect 3426 3703 3429 3823
rect 3426 3603 3429 3616
rect 3378 3523 3381 3546
rect 3386 3426 3389 3566
rect 3402 3563 3413 3566
rect 3402 3436 3405 3563
rect 3434 3546 3437 3843
rect 3442 3803 3445 3906
rect 3442 3696 3445 3746
rect 3450 3716 3453 3906
rect 3458 3903 3461 3926
rect 3470 3836 3473 3963
rect 3490 3913 3493 3926
rect 3470 3833 3477 3836
rect 3458 3736 3461 3816
rect 3466 3743 3469 3816
rect 3474 3743 3477 3833
rect 3482 3813 3485 3876
rect 3498 3836 3501 4083
rect 3506 4003 3509 4016
rect 3514 4003 3517 4036
rect 3530 4003 3533 4016
rect 3546 4003 3549 4173
rect 3566 4136 3569 4193
rect 3562 4133 3569 4136
rect 3490 3833 3501 3836
rect 3458 3733 3477 3736
rect 3474 3723 3477 3733
rect 3482 3716 3485 3806
rect 3490 3753 3493 3833
rect 3498 3796 3501 3816
rect 3506 3803 3509 3816
rect 3514 3796 3517 3806
rect 3498 3793 3517 3796
rect 3522 3746 3525 3886
rect 3514 3743 3525 3746
rect 3450 3713 3461 3716
rect 3442 3693 3449 3696
rect 3446 3606 3449 3693
rect 3418 3526 3421 3546
rect 3414 3523 3421 3526
rect 3426 3543 3437 3546
rect 3442 3603 3449 3606
rect 3414 3456 3417 3523
rect 3414 3453 3421 3456
rect 3402 3433 3413 3436
rect 3366 3393 3373 3396
rect 3378 3423 3389 3426
rect 3366 3316 3369 3393
rect 3378 3323 3381 3423
rect 3394 3353 3397 3406
rect 3410 3376 3413 3433
rect 3402 3373 3413 3376
rect 3386 3323 3389 3346
rect 3366 3313 3373 3316
rect 3370 3293 3373 3313
rect 3402 3306 3405 3373
rect 3418 3366 3421 3453
rect 3394 3303 3405 3306
rect 3410 3363 3421 3366
rect 3346 3243 3357 3246
rect 3394 3246 3397 3303
rect 3394 3243 3405 3246
rect 3346 3146 3349 3243
rect 3370 3166 3373 3206
rect 3342 3143 3349 3146
rect 3366 3163 3373 3166
rect 3342 3036 3345 3143
rect 3342 3033 3349 3036
rect 3314 3013 3341 3016
rect 3314 2956 3317 3006
rect 3330 2973 3333 3006
rect 3314 2953 3325 2956
rect 3314 2933 3317 2946
rect 3322 2926 3325 2953
rect 3314 2923 3325 2926
rect 3298 2843 3305 2846
rect 3266 2833 3277 2836
rect 3266 2813 3269 2833
rect 3302 2776 3305 2843
rect 3266 2756 3269 2776
rect 3298 2773 3305 2776
rect 3266 2753 3277 2756
rect 3258 2693 3261 2746
rect 3274 2696 3277 2753
rect 3266 2693 3277 2696
rect 3266 2673 3269 2693
rect 3234 2633 3245 2636
rect 3234 2593 3237 2633
rect 3242 2613 3245 2626
rect 3258 2613 3277 2616
rect 3282 2613 3285 2626
rect 3226 2583 3237 2586
rect 3226 2513 3229 2526
rect 3234 2506 3237 2583
rect 3226 2503 3237 2506
rect 3186 2393 3197 2396
rect 3162 2363 3173 2366
rect 3154 2343 3161 2346
rect 3158 2236 3161 2343
rect 3122 2213 3133 2216
rect 3142 2213 3149 2216
rect 3154 2233 3161 2236
rect 3114 2133 3117 2166
rect 3122 2116 3125 2213
rect 3130 2133 3133 2206
rect 3142 2136 3145 2213
rect 3154 2146 3157 2233
rect 3170 2216 3173 2363
rect 3186 2236 3189 2393
rect 3186 2233 3197 2236
rect 3170 2213 3181 2216
rect 3154 2143 3165 2146
rect 3138 2133 3145 2136
rect 3118 2113 3125 2116
rect 3118 2036 3121 2113
rect 3118 2033 3125 2036
rect 3114 2003 3117 2016
rect 3090 1973 3097 1976
rect 3074 1963 3085 1966
rect 3074 1913 3077 1926
rect 3018 1903 3025 1906
rect 3018 1883 3021 1903
rect 3082 1873 3085 1963
rect 2998 1753 3005 1756
rect 2970 1713 2981 1716
rect 2986 1713 2989 1726
rect 2970 1666 2973 1713
rect 3002 1666 3005 1753
rect 2970 1663 2981 1666
rect 2978 1633 2981 1663
rect 2998 1663 3005 1666
rect 2946 1523 2949 1616
rect 2970 1593 2973 1606
rect 2986 1586 2989 1616
rect 2978 1583 2989 1586
rect 2962 1533 2965 1546
rect 2922 1433 2933 1436
rect 2906 1403 2909 1426
rect 2914 1346 2917 1406
rect 2930 1366 2933 1433
rect 2890 1313 2893 1336
rect 2898 1296 2901 1346
rect 2894 1293 2901 1296
rect 2906 1343 2917 1346
rect 2922 1363 2933 1366
rect 2922 1343 2925 1363
rect 2954 1346 2957 1526
rect 2970 1506 2973 1526
rect 2966 1503 2973 1506
rect 2966 1436 2969 1503
rect 2966 1433 2973 1436
rect 2970 1413 2973 1433
rect 2978 1406 2981 1583
rect 2998 1566 3001 1663
rect 2994 1563 3001 1566
rect 2986 1423 2989 1536
rect 2994 1516 2997 1563
rect 3002 1533 3005 1546
rect 2994 1513 3001 1516
rect 2998 1416 3001 1513
rect 2970 1403 2981 1406
rect 2994 1413 3001 1416
rect 2930 1343 2957 1346
rect 2874 1273 2885 1276
rect 2862 1263 2869 1266
rect 2866 1236 2869 1263
rect 2866 1233 2873 1236
rect 2858 1013 2861 1226
rect 2870 1186 2873 1233
rect 2866 1183 2873 1186
rect 2802 993 2821 996
rect 2842 1003 2853 1006
rect 2842 936 2845 1003
rect 2842 933 2853 936
rect 2850 846 2853 933
rect 2858 923 2861 1006
rect 2866 906 2869 1183
rect 2882 1166 2885 1273
rect 2894 1246 2897 1293
rect 2906 1256 2909 1343
rect 2914 1273 2917 1336
rect 2922 1303 2925 1326
rect 2906 1253 2917 1256
rect 2894 1243 2901 1246
rect 2898 1173 2901 1243
rect 2874 1163 2885 1166
rect 2874 1126 2877 1163
rect 2882 1143 2901 1146
rect 2882 1133 2885 1143
rect 2890 1126 2893 1136
rect 2874 1123 2893 1126
rect 2898 1123 2901 1143
rect 2874 1013 2877 1066
rect 2882 1003 2885 1016
rect 2890 966 2893 1123
rect 2906 1003 2909 1156
rect 2914 1133 2917 1253
rect 2930 1233 2933 1343
rect 2962 1333 2965 1346
rect 2970 1333 2973 1403
rect 2938 1176 2941 1326
rect 2946 1313 2949 1326
rect 2970 1306 2973 1326
rect 2978 1323 2981 1376
rect 2986 1333 2989 1356
rect 2994 1323 2997 1413
rect 3002 1333 3005 1346
rect 3010 1316 3013 1806
rect 3018 1733 3021 1846
rect 3026 1713 3029 1826
rect 3034 1796 3037 1816
rect 3034 1793 3041 1796
rect 3038 1706 3041 1793
rect 3050 1783 3053 1806
rect 3034 1703 3041 1706
rect 3034 1626 3037 1703
rect 3030 1623 3037 1626
rect 3030 1566 3033 1623
rect 3026 1563 3033 1566
rect 3026 1406 3029 1563
rect 3042 1413 3045 1616
rect 3050 1566 3053 1736
rect 3058 1693 3061 1816
rect 3066 1733 3069 1806
rect 3074 1803 3077 1816
rect 3090 1716 3093 1973
rect 3122 1963 3125 2033
rect 3130 2013 3133 2126
rect 3138 2026 3141 2133
rect 3146 2093 3149 2126
rect 3154 2123 3157 2136
rect 3138 2023 3149 2026
rect 3130 1993 3133 2006
rect 3098 1933 3101 1956
rect 3138 1953 3141 2016
rect 3098 1893 3101 1916
rect 3106 1856 3109 1876
rect 3102 1853 3109 1856
rect 3102 1786 3105 1853
rect 3114 1796 3117 1936
rect 3122 1813 3125 1826
rect 3114 1793 3125 1796
rect 3102 1783 3109 1786
rect 3082 1713 3093 1716
rect 3082 1646 3085 1713
rect 3098 1693 3101 1726
rect 3082 1643 3093 1646
rect 3050 1563 3061 1566
rect 3058 1426 3061 1563
rect 3074 1523 3077 1606
rect 3090 1596 3093 1643
rect 3098 1603 3101 1676
rect 3106 1613 3109 1783
rect 3122 1716 3125 1793
rect 3118 1713 3125 1716
rect 3118 1636 3121 1713
rect 3114 1633 3121 1636
rect 3090 1593 3109 1596
rect 3114 1593 3117 1633
rect 3122 1603 3125 1616
rect 3130 1613 3133 1696
rect 3138 1596 3141 1926
rect 3146 1803 3149 2023
rect 3154 1883 3157 2076
rect 3162 2043 3165 2143
rect 3162 2013 3165 2036
rect 3170 2003 3173 2206
rect 3162 1923 3165 1936
rect 3178 1886 3181 2213
rect 3194 2143 3197 2233
rect 3202 2213 3205 2416
rect 3210 2403 3213 2426
rect 3226 2346 3229 2503
rect 3242 2456 3245 2536
rect 3258 2533 3261 2613
rect 3298 2606 3301 2773
rect 3314 2616 3317 2923
rect 3322 2813 3325 2916
rect 3346 2823 3349 3033
rect 3354 2923 3357 3136
rect 3366 3116 3369 3163
rect 3378 3123 3381 3186
rect 3402 3166 3405 3243
rect 3366 3113 3373 3116
rect 3370 3016 3373 3113
rect 3386 3106 3389 3166
rect 3362 3013 3373 3016
rect 3382 3103 3389 3106
rect 3394 3163 3405 3166
rect 3362 2993 3365 3013
rect 3370 2936 3373 3006
rect 3382 2956 3385 3103
rect 3382 2953 3389 2956
rect 3394 2953 3397 3163
rect 3366 2933 3373 2936
rect 3386 2936 3389 2953
rect 3386 2933 3393 2936
rect 3366 2886 3369 2933
rect 3366 2883 3373 2886
rect 3370 2866 3373 2883
rect 3378 2873 3381 2926
rect 3370 2863 3381 2866
rect 3362 2813 3365 2826
rect 3346 2793 3349 2806
rect 3354 2756 3357 2776
rect 3338 2753 3357 2756
rect 3338 2636 3341 2753
rect 3362 2736 3365 2806
rect 3354 2733 3365 2736
rect 3354 2656 3357 2733
rect 3354 2653 3365 2656
rect 3338 2633 3357 2636
rect 3314 2613 3341 2616
rect 3294 2603 3301 2606
rect 3266 2516 3269 2586
rect 3238 2453 3245 2456
rect 3262 2513 3269 2516
rect 3238 2376 3241 2453
rect 3238 2373 3245 2376
rect 3218 2343 3229 2346
rect 3242 2346 3245 2373
rect 3262 2366 3265 2513
rect 3262 2363 3269 2366
rect 3242 2343 3249 2346
rect 3266 2343 3269 2363
rect 3218 2246 3221 2343
rect 3218 2243 3225 2246
rect 3210 2213 3213 2226
rect 3222 2146 3225 2243
rect 3222 2143 3229 2146
rect 3186 1993 3189 2136
rect 3194 2116 3197 2136
rect 3194 2113 3205 2116
rect 3218 2113 3221 2126
rect 3202 2026 3205 2113
rect 3226 2063 3229 2143
rect 3234 2136 3237 2336
rect 3246 2236 3249 2343
rect 3246 2233 3253 2236
rect 3242 2143 3245 2226
rect 3234 2133 3245 2136
rect 3194 2023 3205 2026
rect 3194 1936 3197 2023
rect 3170 1883 3181 1886
rect 3186 1933 3197 1936
rect 3154 1813 3157 1826
rect 3154 1746 3157 1796
rect 3154 1743 3161 1746
rect 3134 1593 3141 1596
rect 3082 1583 3093 1586
rect 3082 1506 3085 1583
rect 3050 1423 3061 1426
rect 3074 1503 3085 1506
rect 3074 1426 3077 1503
rect 3074 1423 3085 1426
rect 3026 1403 3037 1406
rect 3034 1356 3037 1403
rect 3030 1353 3037 1356
rect 3006 1313 3013 1316
rect 2962 1213 2965 1306
rect 2970 1303 2981 1306
rect 2978 1246 2981 1303
rect 2970 1243 2981 1246
rect 2970 1223 2973 1243
rect 3006 1226 3009 1313
rect 3006 1223 3013 1226
rect 2930 1173 2941 1176
rect 2930 1066 2933 1173
rect 3002 1166 3005 1206
rect 2998 1163 3005 1166
rect 2930 1063 2937 1066
rect 2922 1023 2925 1056
rect 2934 1016 2937 1063
rect 2890 963 2909 966
rect 2866 903 2877 906
rect 2850 843 2861 846
rect 2718 773 2725 776
rect 2646 593 2653 596
rect 2658 683 2677 686
rect 2626 533 2629 546
rect 2634 513 2637 526
rect 2618 503 2625 506
rect 2602 463 2613 466
rect 2586 393 2589 406
rect 2610 403 2613 463
rect 2622 416 2625 503
rect 2646 466 2649 593
rect 2658 476 2661 683
rect 2706 676 2709 726
rect 2698 673 2709 676
rect 2698 626 2701 673
rect 2722 666 2725 773
rect 2746 703 2749 736
rect 2754 723 2757 736
rect 2762 733 2765 756
rect 2770 693 2773 726
rect 2786 723 2789 836
rect 2794 813 2797 826
rect 2818 723 2821 736
rect 2826 733 2829 816
rect 2834 813 2837 826
rect 2842 813 2853 816
rect 2842 733 2845 776
rect 2850 726 2853 736
rect 2842 723 2853 726
rect 2714 663 2725 666
rect 2698 623 2709 626
rect 2682 563 2685 616
rect 2658 473 2665 476
rect 2646 463 2653 466
rect 2622 413 2629 416
rect 2602 333 2621 336
rect 2578 313 2581 326
rect 2526 193 2533 196
rect 2514 166 2517 176
rect 2530 166 2533 193
rect 2474 153 2481 156
rect 2466 133 2469 146
rect 2450 123 2469 126
rect 2478 106 2481 153
rect 2498 123 2501 166
rect 2514 163 2533 166
rect 2562 163 2565 206
rect 2570 203 2573 246
rect 2594 213 2597 246
rect 2514 133 2517 163
rect 2602 153 2605 333
rect 2610 203 2613 286
rect 2618 213 2621 326
rect 2626 283 2629 413
rect 2634 333 2637 416
rect 2562 123 2565 146
rect 2618 143 2621 206
rect 2626 156 2629 216
rect 2634 183 2637 326
rect 2642 323 2645 376
rect 2650 306 2653 463
rect 2662 356 2665 473
rect 2674 393 2677 556
rect 2706 553 2709 623
rect 2698 523 2701 546
rect 2698 406 2701 416
rect 2698 403 2709 406
rect 2698 373 2701 403
rect 2658 353 2665 356
rect 2658 323 2661 353
rect 2650 303 2657 306
rect 2642 203 2645 296
rect 2654 236 2657 303
rect 2650 233 2657 236
rect 2626 153 2637 156
rect 2474 103 2481 106
rect 2474 83 2477 103
rect 2618 0 2621 126
rect 2634 123 2637 153
rect 2642 103 2645 136
rect 2650 123 2653 233
rect 2658 123 2661 216
rect 2666 203 2669 316
rect 2674 303 2677 336
rect 2682 313 2685 326
rect 2698 323 2701 346
rect 2714 333 2717 663
rect 2778 613 2781 626
rect 2730 593 2733 606
rect 2794 536 2797 616
rect 2810 613 2813 706
rect 2842 693 2845 723
rect 2858 716 2861 843
rect 2874 776 2877 903
rect 2882 883 2885 946
rect 2890 813 2893 826
rect 2898 803 2901 816
rect 2874 773 2885 776
rect 2866 723 2869 766
rect 2882 716 2885 773
rect 2898 733 2901 756
rect 2906 733 2909 963
rect 2914 923 2917 1016
rect 2930 1013 2937 1016
rect 2930 943 2933 1013
rect 2946 966 2949 1126
rect 2954 986 2957 1046
rect 2962 1013 2965 1076
rect 2962 996 2965 1006
rect 2970 1003 2973 1046
rect 2978 996 2981 1016
rect 2962 993 2981 996
rect 2954 983 2965 986
rect 2946 963 2953 966
rect 2914 813 2925 816
rect 2922 783 2925 806
rect 2850 713 2861 716
rect 2874 713 2885 716
rect 2786 533 2797 536
rect 2762 423 2765 436
rect 2722 323 2725 336
rect 2730 306 2733 336
rect 2722 303 2733 306
rect 2722 236 2725 303
rect 2722 233 2733 236
rect 2674 213 2693 216
rect 2682 186 2685 206
rect 2698 203 2701 216
rect 2730 213 2733 233
rect 2738 213 2741 416
rect 2762 403 2765 416
rect 2770 403 2773 506
rect 2778 403 2781 416
rect 2746 313 2749 336
rect 2762 243 2773 246
rect 2722 193 2725 206
rect 2754 193 2757 226
rect 2762 223 2765 236
rect 2762 203 2765 216
rect 2770 213 2773 243
rect 2778 233 2781 316
rect 2682 183 2693 186
rect 2674 133 2677 146
rect 2690 133 2693 183
rect 2706 133 2709 176
rect 2682 113 2685 126
rect 2730 123 2733 146
rect 2770 113 2773 206
rect 2786 53 2789 533
rect 2794 513 2797 526
rect 2794 223 2797 436
rect 2802 333 2805 546
rect 2810 543 2813 556
rect 2818 543 2821 616
rect 2826 603 2829 616
rect 2826 593 2837 596
rect 2826 573 2829 593
rect 2842 556 2845 616
rect 2834 553 2845 556
rect 2810 516 2813 536
rect 2834 533 2837 553
rect 2810 513 2817 516
rect 2814 416 2817 513
rect 2810 413 2817 416
rect 2810 266 2813 413
rect 2826 403 2829 526
rect 2834 413 2837 516
rect 2842 396 2845 516
rect 2818 393 2845 396
rect 2818 323 2821 393
rect 2850 376 2853 713
rect 2858 603 2861 636
rect 2866 603 2869 616
rect 2866 583 2869 596
rect 2874 576 2877 713
rect 2914 656 2917 726
rect 2922 703 2925 736
rect 2906 653 2917 656
rect 2890 603 2893 636
rect 2898 613 2901 626
rect 2906 603 2909 653
rect 2914 586 2917 616
rect 2858 573 2877 576
rect 2906 583 2917 586
rect 2858 513 2861 573
rect 2906 506 2909 583
rect 2906 503 2917 506
rect 2842 373 2853 376
rect 2826 313 2829 326
rect 2842 276 2845 373
rect 2842 273 2853 276
rect 2802 263 2813 266
rect 2802 203 2805 236
rect 2810 213 2829 216
rect 2834 213 2837 226
rect 2850 213 2853 273
rect 2858 213 2861 416
rect 2890 413 2893 486
rect 2898 393 2901 406
rect 2906 396 2909 416
rect 2914 403 2917 503
rect 2922 483 2925 616
rect 2930 613 2933 916
rect 2950 886 2953 963
rect 2946 883 2953 886
rect 2938 733 2941 766
rect 2946 723 2949 883
rect 2954 813 2957 826
rect 2962 733 2965 983
rect 2970 906 2973 936
rect 2986 923 2989 1136
rect 2998 1046 3001 1163
rect 3010 1063 3013 1223
rect 3018 1213 3021 1336
rect 3030 1246 3033 1353
rect 3050 1346 3053 1423
rect 3042 1343 3053 1346
rect 3030 1243 3037 1246
rect 3026 1213 3029 1226
rect 3018 1123 3021 1136
rect 2998 1043 3005 1046
rect 2970 903 2981 906
rect 2978 846 2981 903
rect 2970 843 2981 846
rect 2970 813 2973 843
rect 2994 826 2997 1026
rect 3002 903 3005 1043
rect 3010 1036 3013 1056
rect 3026 1053 3029 1126
rect 3034 1053 3037 1243
rect 3042 1096 3045 1343
rect 3050 1323 3053 1336
rect 3058 1303 3061 1326
rect 3050 1116 3053 1216
rect 3066 1203 3069 1406
rect 3074 1213 3077 1326
rect 3082 1286 3085 1423
rect 3090 1413 3093 1536
rect 3098 1423 3101 1526
rect 3106 1516 3109 1593
rect 3134 1546 3137 1593
rect 3146 1553 3149 1736
rect 3158 1646 3161 1743
rect 3154 1643 3161 1646
rect 3134 1543 3141 1546
rect 3114 1523 3117 1536
rect 3106 1513 3113 1516
rect 3110 1436 3113 1513
rect 3110 1433 3117 1436
rect 3098 1363 3101 1416
rect 3106 1383 3109 1406
rect 3114 1373 3117 1433
rect 3122 1403 3125 1526
rect 3138 1436 3141 1543
rect 3138 1433 3145 1436
rect 3130 1403 3133 1426
rect 3142 1386 3145 1433
rect 3138 1383 3145 1386
rect 3098 1303 3101 1326
rect 3122 1303 3125 1366
rect 3138 1363 3141 1383
rect 3154 1353 3157 1643
rect 3162 1613 3165 1626
rect 3170 1596 3173 1883
rect 3186 1813 3189 1933
rect 3194 1916 3197 1926
rect 3202 1923 3205 1936
rect 3210 1916 3213 2006
rect 3218 1933 3221 2016
rect 3226 2003 3229 2016
rect 3234 2013 3237 2126
rect 3242 2013 3245 2133
rect 3250 2076 3253 2233
rect 3258 2216 3261 2326
rect 3274 2223 3277 2536
rect 3282 2523 3285 2566
rect 3294 2556 3297 2603
rect 3294 2553 3301 2556
rect 3298 2533 3301 2553
rect 3282 2376 3285 2416
rect 3306 2403 3309 2596
rect 3314 2523 3317 2606
rect 3322 2436 3325 2556
rect 3330 2513 3333 2606
rect 3338 2596 3341 2613
rect 3338 2593 3345 2596
rect 3342 2506 3345 2593
rect 3338 2503 3345 2506
rect 3322 2433 3333 2436
rect 3322 2413 3325 2426
rect 3330 2406 3333 2433
rect 3322 2403 3333 2406
rect 3282 2373 3293 2376
rect 3290 2323 3293 2373
rect 3298 2323 3301 2336
rect 3306 2306 3309 2396
rect 3314 2313 3317 2326
rect 3298 2303 3309 2306
rect 3258 2213 3269 2216
rect 3258 2096 3261 2136
rect 3274 2113 3277 2206
rect 3282 2193 3285 2236
rect 3298 2156 3301 2303
rect 3314 2286 3317 2306
rect 3310 2283 3317 2286
rect 3310 2196 3313 2283
rect 3322 2203 3325 2403
rect 3338 2393 3341 2503
rect 3354 2486 3357 2633
rect 3350 2483 3357 2486
rect 3310 2193 3317 2196
rect 3298 2153 3309 2156
rect 3282 2123 3285 2136
rect 3290 2116 3293 2136
rect 3282 2113 3293 2116
rect 3258 2093 3269 2096
rect 3250 2073 3257 2076
rect 3254 2016 3257 2073
rect 3250 2013 3257 2016
rect 3250 1996 3253 2013
rect 3242 1993 3253 1996
rect 3194 1913 3213 1916
rect 3186 1686 3189 1756
rect 3210 1746 3213 1876
rect 3226 1863 3229 1936
rect 3242 1926 3245 1993
rect 3266 1986 3269 2093
rect 3282 2046 3285 2113
rect 3306 2106 3309 2153
rect 3258 1983 3269 1986
rect 3278 2043 3285 2046
rect 3298 2103 3309 2106
rect 3258 1933 3261 1983
rect 3278 1946 3281 2043
rect 3298 2036 3301 2103
rect 3290 2033 3301 2036
rect 3278 1943 3285 1946
rect 3242 1923 3253 1926
rect 3218 1793 3221 1806
rect 3210 1743 3217 1746
rect 3186 1683 3205 1686
rect 3166 1593 3173 1596
rect 3166 1466 3169 1593
rect 3166 1463 3173 1466
rect 3170 1443 3173 1463
rect 3178 1426 3181 1676
rect 3202 1603 3205 1683
rect 3214 1656 3217 1743
rect 3226 1723 3229 1816
rect 3250 1813 3253 1923
rect 3274 1833 3277 1926
rect 3234 1733 3237 1806
rect 3242 1793 3245 1806
rect 3258 1753 3261 1796
rect 3234 1713 3237 1726
rect 3258 1723 3269 1726
rect 3274 1713 3277 1726
rect 3214 1653 3237 1656
rect 3234 1596 3237 1653
rect 3226 1593 3237 1596
rect 3174 1423 3181 1426
rect 3082 1283 3093 1286
rect 3082 1203 3085 1276
rect 3090 1213 3093 1283
rect 3098 1276 3101 1296
rect 3146 1276 3149 1336
rect 3098 1273 3117 1276
rect 3114 1176 3117 1273
rect 3098 1173 3117 1176
rect 3138 1273 3149 1276
rect 3138 1176 3141 1273
rect 3138 1173 3149 1176
rect 3058 1123 3061 1136
rect 3050 1113 3061 1116
rect 3042 1093 3049 1096
rect 3046 1046 3049 1093
rect 3042 1043 3049 1046
rect 3010 1033 3021 1036
rect 3018 966 3021 1033
rect 3042 993 3045 1043
rect 3010 963 3021 966
rect 3010 833 3013 963
rect 3058 946 3061 1113
rect 3066 1096 3069 1136
rect 3090 1133 3093 1166
rect 3082 1113 3085 1126
rect 3066 1093 3077 1096
rect 3098 1093 3101 1173
rect 3074 1026 3077 1093
rect 3066 1023 3077 1026
rect 3066 1003 3069 1023
rect 3106 1013 3109 1136
rect 3122 1133 3125 1146
rect 3146 1143 3149 1173
rect 3162 1106 3165 1366
rect 3174 1316 3177 1423
rect 3186 1403 3189 1416
rect 3202 1413 3205 1526
rect 3218 1433 3221 1536
rect 3226 1376 3229 1593
rect 3250 1543 3253 1616
rect 3250 1523 3253 1536
rect 3234 1396 3237 1416
rect 3234 1393 3245 1396
rect 3174 1313 3181 1316
rect 3178 1293 3181 1313
rect 3186 1276 3189 1356
rect 3178 1273 3189 1276
rect 3178 1176 3181 1273
rect 3178 1173 3189 1176
rect 3170 1123 3173 1136
rect 3186 1116 3189 1173
rect 3194 1146 3197 1336
rect 3202 1333 3213 1336
rect 3202 1303 3205 1326
rect 3218 1323 3221 1376
rect 3226 1373 3233 1376
rect 3230 1316 3233 1373
rect 3226 1313 3233 1316
rect 3226 1256 3229 1313
rect 3218 1253 3229 1256
rect 3194 1143 3205 1146
rect 3202 1136 3205 1143
rect 3202 1133 3213 1136
rect 3202 1123 3205 1133
rect 3186 1113 3205 1116
rect 3138 1076 3141 1096
rect 3130 1073 3141 1076
rect 3130 1016 3133 1073
rect 3130 1013 3141 1016
rect 3018 896 3021 926
rect 3018 893 3029 896
rect 2986 823 3005 826
rect 2986 813 2989 823
rect 2994 806 2997 816
rect 2978 803 2997 806
rect 2978 753 2981 803
rect 3002 766 3005 823
rect 3026 813 3029 893
rect 3034 876 3037 946
rect 3058 943 3065 946
rect 3062 896 3065 943
rect 3058 893 3065 896
rect 3034 873 3045 876
rect 3058 873 3061 893
rect 3042 806 3045 873
rect 3034 803 3045 806
rect 2994 763 3005 766
rect 2970 743 2989 746
rect 2954 673 2957 726
rect 2970 723 2973 743
rect 2978 723 2981 736
rect 2986 733 2989 743
rect 2994 723 2997 763
rect 3010 756 3013 766
rect 3002 753 3013 756
rect 3034 753 3037 803
rect 3074 756 3077 926
rect 3082 913 3085 926
rect 3106 916 3109 996
rect 3114 923 3117 996
rect 3106 913 3117 916
rect 3122 913 3125 926
rect 3138 913 3141 1013
rect 3146 933 3149 946
rect 3154 936 3157 1106
rect 3162 1103 3169 1106
rect 3166 1036 3169 1103
rect 3162 1033 3169 1036
rect 3162 973 3165 1033
rect 3170 943 3173 1016
rect 3186 983 3189 1016
rect 3154 933 3165 936
rect 3090 813 3093 836
rect 3090 783 3093 806
rect 3098 803 3109 806
rect 3114 763 3117 913
rect 3122 803 3125 826
rect 3130 813 3133 896
rect 3130 773 3133 806
rect 3146 796 3149 816
rect 3154 803 3157 926
rect 3162 813 3165 933
rect 3162 796 3165 806
rect 3146 793 3165 796
rect 3074 753 3085 756
rect 3002 733 3005 753
rect 3018 723 3021 736
rect 3026 723 3037 726
rect 3058 723 3061 736
rect 2930 533 2933 606
rect 2954 533 2957 616
rect 2962 603 2965 616
rect 2994 603 2997 616
rect 3010 576 3013 656
rect 3010 573 3021 576
rect 3018 516 3021 573
rect 3034 523 3037 616
rect 3018 513 3029 516
rect 2922 413 2925 436
rect 2922 396 2925 406
rect 2906 393 2925 396
rect 2866 333 2869 346
rect 2874 343 2893 346
rect 2874 323 2877 343
rect 2882 226 2885 336
rect 2890 333 2893 343
rect 2898 323 2901 366
rect 2906 313 2909 326
rect 2914 323 2917 346
rect 2930 323 2933 416
rect 2938 413 2941 426
rect 2946 393 2949 416
rect 2978 413 2981 426
rect 2946 313 2949 326
rect 2882 223 2893 226
rect 2810 193 2813 206
rect 2826 203 2829 213
rect 2826 183 2829 196
rect 2842 133 2845 166
rect 2802 113 2805 126
rect 2850 113 2853 126
rect 2858 123 2861 206
rect 2882 163 2885 216
rect 2890 203 2893 223
rect 2898 203 2901 216
rect 2906 213 2909 226
rect 2938 193 2941 206
rect 2946 156 2949 216
rect 2954 203 2957 216
rect 2962 213 2965 246
rect 2970 213 2973 256
rect 2962 193 2965 206
rect 2946 153 2957 156
rect 2938 133 2941 146
rect 2954 133 2957 153
rect 2994 133 2997 346
rect 3026 343 3029 513
rect 3050 413 3053 536
rect 3066 533 3069 556
rect 3058 513 3061 526
rect 3050 336 3053 406
rect 3082 393 3085 753
rect 3106 753 3133 756
rect 3106 733 3109 753
rect 3130 733 3133 753
rect 3090 593 3093 616
rect 3130 593 3133 606
rect 3138 586 3141 686
rect 3130 583 3141 586
rect 3146 583 3149 606
rect 3106 523 3109 536
rect 3114 523 3117 536
rect 3122 496 3125 536
rect 3130 513 3133 583
rect 3154 576 3157 766
rect 3162 613 3165 726
rect 3138 533 3141 576
rect 3146 573 3157 576
rect 3146 523 3149 573
rect 3154 533 3157 546
rect 3162 533 3165 596
rect 3170 573 3173 916
rect 3186 886 3189 976
rect 3202 936 3205 1113
rect 3210 1103 3213 1126
rect 3218 1093 3221 1253
rect 3242 1246 3245 1393
rect 3250 1333 3253 1416
rect 3258 1343 3261 1406
rect 3242 1243 3261 1246
rect 3226 1113 3229 1126
rect 3234 1016 3237 1206
rect 3242 1133 3245 1243
rect 3266 1203 3269 1536
rect 3274 1523 3277 1546
rect 3274 1413 3277 1436
rect 3282 1423 3285 1943
rect 3290 1923 3293 2033
rect 3298 1993 3301 2006
rect 3306 1973 3309 2016
rect 3298 1933 3301 1966
rect 3314 1936 3317 2193
rect 3322 2013 3325 2146
rect 3330 2126 3333 2386
rect 3350 2336 3353 2483
rect 3362 2343 3365 2653
rect 3338 2316 3341 2336
rect 3350 2333 3357 2336
rect 3338 2313 3345 2316
rect 3342 2236 3345 2313
rect 3354 2303 3357 2333
rect 3338 2233 3345 2236
rect 3370 2236 3373 2826
rect 3378 2493 3381 2863
rect 3390 2826 3393 2933
rect 3386 2823 3393 2826
rect 3386 2803 3389 2823
rect 3394 2793 3397 2806
rect 3402 2773 3405 3156
rect 3386 2716 3389 2736
rect 3386 2713 3393 2716
rect 3390 2566 3393 2713
rect 3386 2563 3393 2566
rect 3386 2506 3389 2563
rect 3386 2503 3393 2506
rect 3390 2416 3393 2503
rect 3390 2413 3397 2416
rect 3378 2336 3381 2406
rect 3394 2393 3397 2413
rect 3402 2403 3405 2756
rect 3410 2583 3413 3363
rect 3426 3336 3429 3543
rect 3434 3513 3437 3536
rect 3426 3333 3437 3336
rect 3426 3303 3429 3326
rect 3418 3203 3421 3216
rect 3426 3213 3429 3296
rect 3418 3083 3421 3156
rect 3426 3133 3429 3146
rect 3434 3093 3437 3333
rect 3442 3106 3445 3603
rect 3458 3586 3461 3713
rect 3474 3713 3485 3716
rect 3474 3593 3477 3713
rect 3498 3626 3501 3736
rect 3498 3623 3505 3626
rect 3450 3583 3461 3586
rect 3450 3563 3453 3583
rect 3458 3413 3461 3536
rect 3482 3506 3485 3526
rect 3490 3523 3493 3616
rect 3502 3546 3505 3623
rect 3514 3613 3517 3743
rect 3498 3543 3505 3546
rect 3482 3503 3493 3506
rect 3474 3446 3477 3466
rect 3470 3443 3477 3446
rect 3470 3376 3473 3443
rect 3490 3413 3493 3503
rect 3498 3496 3501 3543
rect 3514 3533 3517 3596
rect 3506 3513 3509 3526
rect 3498 3493 3505 3496
rect 3502 3406 3505 3493
rect 3530 3456 3533 3856
rect 3538 3813 3541 3946
rect 3562 3906 3565 4133
rect 3570 4113 3573 4126
rect 3578 3946 3581 4223
rect 3586 4123 3589 4206
rect 3610 4203 3613 4223
rect 3618 4186 3621 4296
rect 3634 4223 3637 4356
rect 3626 4213 3637 4216
rect 3614 4183 3621 4186
rect 3594 4106 3597 4146
rect 3590 4103 3597 4106
rect 3590 4006 3593 4103
rect 3590 4003 3597 4006
rect 3594 3983 3597 4003
rect 3554 3903 3565 3906
rect 3574 3943 3581 3946
rect 3554 3846 3557 3903
rect 3574 3896 3577 3943
rect 3586 3923 3589 3936
rect 3574 3893 3581 3896
rect 3578 3873 3581 3893
rect 3594 3876 3597 3926
rect 3602 3883 3605 4116
rect 3614 4056 3617 4183
rect 3626 4066 3629 4206
rect 3634 4083 3637 4213
rect 3650 4203 3653 4436
rect 3706 4416 3709 4586
rect 3786 4583 3789 4606
rect 3810 4546 3813 4623
rect 3826 4606 3829 4616
rect 3882 4613 3885 4740
rect 3930 4623 3933 4740
rect 3826 4603 3837 4606
rect 3810 4543 3821 4546
rect 3722 4506 3725 4526
rect 3818 4523 3821 4543
rect 3722 4503 3733 4506
rect 3730 4446 3733 4503
rect 3826 4476 3829 4596
rect 3834 4553 3837 4603
rect 3850 4533 3853 4576
rect 3906 4573 3909 4606
rect 3922 4563 3925 4616
rect 3954 4613 3957 4626
rect 4050 4613 4053 4740
rect 4194 4633 4197 4740
rect 3754 4446 3757 4466
rect 3722 4443 3733 4446
rect 3750 4443 3757 4446
rect 3706 4413 3713 4416
rect 3674 4373 3677 4406
rect 3658 4333 3661 4346
rect 3666 4323 3669 4356
rect 3698 4323 3701 4406
rect 3710 4346 3713 4413
rect 3722 4403 3725 4443
rect 3730 4413 3733 4426
rect 3706 4343 3713 4346
rect 3738 4343 3741 4416
rect 3750 4376 3753 4443
rect 3770 4413 3773 4426
rect 3750 4373 3757 4376
rect 3674 4203 3677 4226
rect 3658 4133 3661 4146
rect 3642 4103 3645 4126
rect 3626 4063 3637 4066
rect 3614 4053 3621 4056
rect 3618 3946 3621 4053
rect 3634 3946 3637 4063
rect 3650 3993 3653 4006
rect 3666 3986 3669 4006
rect 3610 3943 3621 3946
rect 3626 3943 3637 3946
rect 3594 3873 3605 3876
rect 3546 3843 3557 3846
rect 3546 3483 3549 3843
rect 3554 3723 3557 3816
rect 3570 3743 3573 3816
rect 3602 3813 3605 3873
rect 3610 3836 3613 3943
rect 3618 3843 3621 3936
rect 3626 3853 3629 3943
rect 3650 3933 3653 3986
rect 3662 3983 3669 3986
rect 3634 3923 3645 3926
rect 3634 3896 3637 3916
rect 3634 3893 3641 3896
rect 3610 3833 3617 3836
rect 3614 3786 3617 3833
rect 3638 3796 3641 3893
rect 3634 3793 3641 3796
rect 3614 3783 3621 3786
rect 3618 3766 3621 3783
rect 3618 3763 3625 3766
rect 3594 3733 3597 3746
rect 3554 3676 3557 3706
rect 3554 3673 3573 3676
rect 3570 3556 3573 3673
rect 3554 3553 3573 3556
rect 3530 3453 3541 3456
rect 3498 3403 3505 3406
rect 3470 3373 3477 3376
rect 3450 3213 3453 3366
rect 3474 3296 3477 3373
rect 3498 3346 3501 3403
rect 3494 3343 3501 3346
rect 3514 3346 3517 3446
rect 3538 3413 3541 3453
rect 3514 3343 3525 3346
rect 3474 3293 3485 3296
rect 3458 3183 3461 3216
rect 3482 3203 3485 3293
rect 3494 3236 3497 3343
rect 3494 3233 3501 3236
rect 3490 3183 3493 3216
rect 3450 3123 3453 3136
rect 3442 3103 3449 3106
rect 3446 3046 3449 3103
rect 3446 3043 3453 3046
rect 3426 2966 3429 3006
rect 3450 2996 3453 3043
rect 3458 3013 3461 3126
rect 3466 3123 3469 3176
rect 3490 3116 3493 3136
rect 3482 3113 3493 3116
rect 3482 3066 3485 3113
rect 3498 3106 3501 3233
rect 3506 3213 3509 3336
rect 3522 3206 3525 3343
rect 3514 3203 3525 3206
rect 3514 3173 3517 3203
rect 3506 3123 3509 3146
rect 3498 3103 3505 3106
rect 3482 3063 3493 3066
rect 3490 3013 3493 3063
rect 3502 3006 3505 3103
rect 3514 3013 3517 3136
rect 3538 3126 3541 3406
rect 3546 3213 3549 3236
rect 3522 3103 3525 3126
rect 3538 3123 3545 3126
rect 3530 3053 3533 3116
rect 3542 3076 3545 3123
rect 3538 3073 3545 3076
rect 3538 3036 3541 3073
rect 3530 3033 3541 3036
rect 3442 2993 3453 2996
rect 3426 2963 3433 2966
rect 3418 2716 3421 2956
rect 3430 2826 3433 2963
rect 3426 2823 3433 2826
rect 3426 2753 3429 2823
rect 3442 2816 3445 2993
rect 3458 2933 3461 2946
rect 3466 2926 3469 3006
rect 3498 3003 3505 3006
rect 3474 2943 3477 2996
rect 3498 2936 3501 3003
rect 3530 2976 3533 3033
rect 3530 2973 3541 2976
rect 3498 2933 3509 2936
rect 3450 2923 3477 2926
rect 3442 2813 3453 2816
rect 3434 2733 3437 2806
rect 3450 2726 3453 2813
rect 3442 2723 3453 2726
rect 3418 2713 3429 2716
rect 3426 2636 3429 2713
rect 3418 2633 3429 2636
rect 3418 2546 3421 2633
rect 3442 2626 3445 2723
rect 3442 2623 3453 2626
rect 3418 2543 3429 2546
rect 3418 2376 3421 2496
rect 3426 2453 3429 2543
rect 3434 2523 3437 2616
rect 3450 2576 3453 2623
rect 3446 2573 3453 2576
rect 3446 2496 3449 2573
rect 3466 2546 3469 2923
rect 3482 2803 3485 2926
rect 3506 2826 3509 2933
rect 3538 2876 3541 2973
rect 3498 2823 3509 2826
rect 3530 2873 3541 2876
rect 3498 2806 3501 2823
rect 3494 2803 3501 2806
rect 3494 2746 3497 2803
rect 3494 2743 3501 2746
rect 3490 2563 3493 2726
rect 3498 2706 3501 2743
rect 3506 2723 3509 2806
rect 3498 2703 3509 2706
rect 3506 2636 3509 2703
rect 3498 2633 3509 2636
rect 3530 2636 3533 2873
rect 3546 2856 3549 3056
rect 3554 2936 3557 3553
rect 3594 3546 3597 3726
rect 3610 3696 3613 3756
rect 3606 3693 3613 3696
rect 3606 3596 3609 3693
rect 3622 3686 3625 3763
rect 3618 3683 3625 3686
rect 3618 3603 3621 3683
rect 3634 3603 3637 3793
rect 3650 3776 3653 3846
rect 3662 3836 3665 3983
rect 3662 3833 3669 3836
rect 3642 3773 3653 3776
rect 3642 3733 3645 3773
rect 3658 3753 3661 3816
rect 3666 3726 3669 3833
rect 3606 3593 3613 3596
rect 3590 3543 3597 3546
rect 3562 3443 3565 3526
rect 3570 3453 3573 3536
rect 3578 3436 3581 3526
rect 3590 3446 3593 3543
rect 3590 3443 3597 3446
rect 3562 3256 3565 3436
rect 3570 3433 3581 3436
rect 3570 3403 3573 3433
rect 3562 3253 3569 3256
rect 3566 3106 3569 3253
rect 3578 3193 3581 3416
rect 3586 3413 3589 3426
rect 3594 3256 3597 3443
rect 3602 3413 3605 3536
rect 3602 3313 3605 3326
rect 3594 3253 3601 3256
rect 3586 3223 3589 3246
rect 3562 3103 3569 3106
rect 3562 3083 3565 3103
rect 3570 2963 3573 3026
rect 3578 3013 3581 3106
rect 3586 2956 3589 3206
rect 3598 3156 3601 3253
rect 3594 3153 3601 3156
rect 3594 3106 3597 3153
rect 3602 3123 3605 3136
rect 3594 3103 3601 3106
rect 3598 3036 3601 3103
rect 3598 3033 3605 3036
rect 3594 3003 3597 3026
rect 3602 2993 3605 3033
rect 3586 2953 3605 2956
rect 3554 2933 3565 2936
rect 3542 2853 3549 2856
rect 3542 2806 3545 2853
rect 3554 2813 3557 2926
rect 3562 2886 3565 2933
rect 3586 2923 3589 2946
rect 3562 2883 3569 2886
rect 3566 2806 3569 2883
rect 3542 2803 3549 2806
rect 3546 2683 3549 2803
rect 3562 2803 3569 2806
rect 3530 2633 3541 2636
rect 3466 2543 3477 2546
rect 3442 2493 3449 2496
rect 3442 2473 3445 2493
rect 3474 2466 3477 2543
rect 3466 2463 3477 2466
rect 3450 2436 3453 2456
rect 3466 2436 3469 2463
rect 3498 2453 3501 2633
rect 3538 2616 3541 2633
rect 3506 2523 3509 2616
rect 3514 2596 3517 2606
rect 3522 2603 3525 2616
rect 3530 2596 3533 2616
rect 3538 2613 3549 2616
rect 3514 2593 3533 2596
rect 3514 2566 3517 2586
rect 3514 2563 3521 2566
rect 3518 2516 3521 2563
rect 3538 2553 3541 2606
rect 3538 2526 3541 2536
rect 3514 2513 3521 2516
rect 3530 2523 3541 2526
rect 3446 2433 3453 2436
rect 3458 2433 3469 2436
rect 3402 2373 3421 2376
rect 3378 2333 3389 2336
rect 3402 2333 3405 2373
rect 3386 2306 3389 2333
rect 3386 2303 3397 2306
rect 3386 2246 3389 2296
rect 3394 2276 3397 2303
rect 3394 2273 3405 2276
rect 3386 2243 3393 2246
rect 3370 2233 3381 2236
rect 3338 2213 3341 2233
rect 3354 2143 3357 2206
rect 3362 2126 3365 2216
rect 3378 2213 3381 2233
rect 3330 2123 3341 2126
rect 3338 2036 3341 2123
rect 3354 2123 3365 2126
rect 3354 2046 3357 2123
rect 3354 2043 3365 2046
rect 3334 2033 3341 2036
rect 3306 1933 3317 1936
rect 3306 1916 3309 1933
rect 3302 1913 3309 1916
rect 3290 1793 3293 1896
rect 3302 1826 3305 1913
rect 3314 1863 3317 1926
rect 3298 1823 3305 1826
rect 3298 1776 3301 1823
rect 3294 1773 3301 1776
rect 3294 1556 3297 1773
rect 3294 1553 3301 1556
rect 3298 1533 3301 1553
rect 3298 1506 3301 1526
rect 3294 1503 3301 1506
rect 3294 1426 3297 1503
rect 3294 1423 3301 1426
rect 3290 1386 3293 1406
rect 3298 1403 3301 1423
rect 3290 1383 3297 1386
rect 3274 1303 3277 1326
rect 3282 1323 3285 1356
rect 3294 1316 3297 1383
rect 3306 1363 3309 1816
rect 3314 1786 3317 1826
rect 3322 1803 3325 2006
rect 3334 1846 3337 2033
rect 3362 2023 3365 2043
rect 3330 1843 3337 1846
rect 3330 1823 3333 1843
rect 3346 1826 3349 2016
rect 3354 1923 3357 1946
rect 3362 1923 3365 1986
rect 3370 1906 3373 2206
rect 3378 2183 3381 2206
rect 3390 2186 3393 2243
rect 3386 2183 3393 2186
rect 3366 1903 3373 1906
rect 3342 1823 3349 1826
rect 3314 1783 3321 1786
rect 3318 1686 3321 1783
rect 3314 1683 3321 1686
rect 3314 1663 3317 1683
rect 3290 1313 3297 1316
rect 3250 1123 3253 1136
rect 3226 1013 3237 1016
rect 3226 1003 3229 1013
rect 3234 966 3237 1006
rect 3242 996 3245 1016
rect 3250 1003 3253 1016
rect 3258 996 3261 1006
rect 3242 993 3261 996
rect 3234 963 3253 966
rect 3182 883 3189 886
rect 3198 933 3205 936
rect 3182 776 3185 883
rect 3198 836 3201 933
rect 3198 833 3205 836
rect 3178 773 3185 776
rect 3178 683 3181 773
rect 3194 676 3197 816
rect 3202 763 3205 833
rect 3210 813 3213 926
rect 3234 923 3237 936
rect 3226 813 3229 836
rect 3218 736 3221 776
rect 3250 763 3253 963
rect 3266 933 3269 1126
rect 3290 1106 3293 1313
rect 3314 1136 3317 1656
rect 3330 1626 3333 1816
rect 3342 1766 3345 1823
rect 3342 1763 3349 1766
rect 3338 1726 3341 1736
rect 3346 1733 3349 1763
rect 3338 1723 3349 1726
rect 3354 1723 3357 1836
rect 3366 1766 3369 1903
rect 3366 1763 3373 1766
rect 3370 1743 3373 1763
rect 3346 1656 3349 1723
rect 3346 1653 3357 1656
rect 3322 1623 3333 1626
rect 3322 1396 3325 1623
rect 3330 1533 3333 1616
rect 3338 1613 3341 1636
rect 3330 1413 3333 1436
rect 3338 1403 3341 1606
rect 3346 1603 3349 1626
rect 3354 1613 3357 1653
rect 3362 1553 3365 1726
rect 3370 1623 3373 1726
rect 3346 1413 3349 1526
rect 3354 1403 3357 1536
rect 3370 1446 3373 1606
rect 3378 1546 3381 2116
rect 3386 2013 3389 2183
rect 3402 2166 3405 2273
rect 3394 2163 3405 2166
rect 3394 2116 3397 2163
rect 3410 2133 3413 2146
rect 3418 2133 3421 2216
rect 3434 2116 3437 2396
rect 3446 2346 3449 2433
rect 3458 2393 3461 2433
rect 3466 2413 3469 2426
rect 3490 2413 3501 2416
rect 3506 2413 3509 2426
rect 3490 2376 3493 2413
rect 3470 2373 3493 2376
rect 3446 2343 3453 2346
rect 3442 2313 3445 2326
rect 3442 2123 3445 2146
rect 3394 2113 3405 2116
rect 3402 2036 3405 2113
rect 3394 2033 3405 2036
rect 3426 2113 3437 2116
rect 3426 2036 3429 2113
rect 3426 2033 3437 2036
rect 3394 2013 3397 2033
rect 3402 1953 3405 2006
rect 3410 2003 3413 2016
rect 3418 1936 3421 2006
rect 3426 1993 3429 2006
rect 3386 1916 3389 1936
rect 3386 1913 3393 1916
rect 3390 1856 3393 1913
rect 3386 1853 3393 1856
rect 3386 1813 3389 1853
rect 3402 1836 3405 1936
rect 3418 1933 3425 1936
rect 3410 1903 3413 1926
rect 3422 1876 3425 1933
rect 3418 1873 3425 1876
rect 3418 1853 3421 1873
rect 3394 1833 3405 1836
rect 3394 1793 3397 1833
rect 3434 1823 3437 2033
rect 3450 2013 3453 2343
rect 3470 2286 3473 2373
rect 3482 2323 3485 2336
rect 3490 2313 3493 2326
rect 3466 2283 3473 2286
rect 3458 2143 3461 2196
rect 3466 2186 3469 2283
rect 3474 2213 3477 2226
rect 3482 2203 3485 2306
rect 3466 2183 3477 2186
rect 3474 2133 3477 2183
rect 3490 2156 3493 2216
rect 3498 2193 3501 2206
rect 3506 2203 3509 2216
rect 3514 2203 3517 2513
rect 3530 2496 3533 2523
rect 3546 2516 3549 2613
rect 3554 2603 3557 2736
rect 3562 2686 3565 2803
rect 3570 2703 3573 2726
rect 3562 2683 3569 2686
rect 3566 2596 3569 2683
rect 3562 2593 3569 2596
rect 3526 2493 3533 2496
rect 3538 2513 3549 2516
rect 3554 2513 3557 2526
rect 3526 2406 3529 2493
rect 3538 2416 3541 2513
rect 3538 2413 3545 2416
rect 3526 2403 3533 2406
rect 3530 2383 3533 2403
rect 3542 2356 3545 2413
rect 3554 2393 3557 2416
rect 3530 2333 3533 2356
rect 3538 2353 3545 2356
rect 3482 2153 3493 2156
rect 3474 2106 3477 2126
rect 3466 2103 3477 2106
rect 3466 1976 3469 2103
rect 3482 1983 3485 2153
rect 3522 2146 3525 2236
rect 3530 2223 3533 2326
rect 3510 2143 3525 2146
rect 3490 1993 3493 2006
rect 3466 1973 3477 1976
rect 3410 1793 3413 1806
rect 3386 1603 3389 1736
rect 3394 1726 3397 1746
rect 3394 1723 3405 1726
rect 3402 1646 3405 1723
rect 3394 1643 3405 1646
rect 3394 1563 3397 1643
rect 3402 1613 3405 1626
rect 3378 1543 3389 1546
rect 3362 1443 3373 1446
rect 3362 1413 3365 1443
rect 3322 1393 3329 1396
rect 3326 1336 3329 1393
rect 3326 1333 3333 1336
rect 3322 1303 3325 1326
rect 3330 1323 3333 1333
rect 3338 1226 3341 1366
rect 3362 1333 3365 1406
rect 3370 1403 3373 1426
rect 3386 1396 3389 1543
rect 3410 1526 3413 1546
rect 3402 1523 3413 1526
rect 3402 1446 3405 1523
rect 3418 1456 3421 1736
rect 3426 1713 3429 1736
rect 3434 1723 3437 1816
rect 3442 1676 3445 1906
rect 3434 1673 3445 1676
rect 3426 1573 3429 1596
rect 3434 1526 3437 1673
rect 3450 1656 3453 1926
rect 3474 1856 3477 1973
rect 3446 1653 3453 1656
rect 3446 1556 3449 1653
rect 3446 1553 3453 1556
rect 3426 1523 3437 1526
rect 3418 1453 3429 1456
rect 3402 1443 3413 1446
rect 3410 1426 3413 1443
rect 3378 1393 3389 1396
rect 3378 1356 3381 1393
rect 3378 1353 3385 1356
rect 3330 1223 3341 1226
rect 3330 1156 3333 1223
rect 3330 1153 3341 1156
rect 3298 1113 3301 1136
rect 3314 1133 3325 1136
rect 3290 1103 3301 1106
rect 3274 926 3277 1016
rect 3298 1006 3301 1103
rect 3306 1033 3309 1126
rect 3322 1036 3325 1133
rect 3314 1033 3325 1036
rect 3306 1013 3309 1026
rect 3298 1003 3309 1006
rect 3266 923 3277 926
rect 3282 943 3301 946
rect 3282 923 3285 943
rect 3290 923 3293 936
rect 3298 933 3301 943
rect 3202 733 3221 736
rect 3202 716 3205 733
rect 3202 713 3209 716
rect 3190 673 3197 676
rect 3178 583 3181 606
rect 3190 546 3193 673
rect 3206 666 3209 713
rect 3202 663 3209 666
rect 3202 583 3205 663
rect 3190 543 3197 546
rect 3122 493 3133 496
rect 3098 413 3101 426
rect 3002 223 3005 236
rect 3010 203 3013 326
rect 3026 316 3029 336
rect 3050 333 3061 336
rect 3074 333 3077 346
rect 3026 313 3037 316
rect 3034 246 3037 313
rect 3026 243 3037 246
rect 2890 113 2893 126
rect 2978 113 2981 126
rect 3018 113 3021 126
rect 3026 33 3029 243
rect 3058 173 3061 333
rect 3082 323 3085 336
rect 3098 333 3101 356
rect 3090 283 3093 326
rect 3106 293 3109 326
rect 3114 313 3117 416
rect 3130 413 3133 493
rect 3138 413 3141 426
rect 3106 213 3109 226
rect 3138 213 3141 326
rect 3146 303 3149 416
rect 3154 413 3157 526
rect 3194 523 3197 543
rect 3202 506 3205 576
rect 3210 523 3213 606
rect 3218 593 3221 726
rect 3226 723 3229 756
rect 3242 633 3245 756
rect 3258 746 3261 816
rect 3266 783 3269 806
rect 3258 743 3269 746
rect 3266 733 3269 743
rect 3266 613 3269 726
rect 3194 503 3205 506
rect 3194 436 3197 503
rect 3154 396 3157 406
rect 3162 403 3165 436
rect 3194 433 3205 436
rect 3170 396 3173 416
rect 3154 393 3173 396
rect 3170 306 3173 326
rect 3162 303 3173 306
rect 3162 236 3165 303
rect 3162 233 3173 236
rect 3146 213 3149 226
rect 3154 203 3157 216
rect 3170 203 3173 233
rect 3178 203 3181 406
rect 3186 363 3189 416
rect 3186 323 3189 346
rect 3194 323 3197 406
rect 3202 293 3205 433
rect 3218 403 3221 586
rect 3226 533 3229 606
rect 3266 516 3269 536
rect 3258 513 3269 516
rect 3258 436 3261 513
rect 3258 433 3269 436
rect 3266 416 3269 433
rect 3274 423 3277 923
rect 3306 876 3309 1003
rect 3314 996 3317 1033
rect 3322 1013 3333 1016
rect 3338 1006 3341 1153
rect 3346 1133 3349 1216
rect 3362 1133 3365 1326
rect 3382 1306 3385 1353
rect 3378 1303 3385 1306
rect 3370 1113 3373 1126
rect 3378 1046 3381 1303
rect 3394 1226 3397 1346
rect 3402 1343 3405 1426
rect 3410 1423 3417 1426
rect 3414 1366 3417 1423
rect 3410 1363 3417 1366
rect 3410 1316 3413 1363
rect 3426 1346 3429 1453
rect 3442 1423 3445 1536
rect 3450 1523 3453 1553
rect 3458 1456 3461 1856
rect 3474 1853 3481 1856
rect 3478 1776 3481 1853
rect 3474 1773 3481 1776
rect 3466 1513 3469 1756
rect 3474 1733 3477 1773
rect 3490 1756 3493 1936
rect 3498 1933 3501 2106
rect 3510 2046 3513 2143
rect 3506 2043 3513 2046
rect 3482 1753 3493 1756
rect 3482 1733 3485 1753
rect 3474 1623 3477 1726
rect 3490 1713 3493 1726
rect 3498 1693 3501 1736
rect 3506 1733 3509 2043
rect 3514 1996 3517 2026
rect 3522 2003 3525 2136
rect 3530 2023 3533 2206
rect 3538 2086 3541 2353
rect 3546 2103 3549 2336
rect 3554 2113 3557 2386
rect 3562 2296 3565 2593
rect 3578 2533 3581 2836
rect 3586 2736 3589 2816
rect 3594 2753 3597 2826
rect 3602 2763 3605 2953
rect 3610 2753 3613 3593
rect 3618 3323 3621 3536
rect 3634 3413 3637 3426
rect 3634 3333 3637 3346
rect 3642 3333 3645 3726
rect 3658 3723 3669 3726
rect 3658 3713 3669 3716
rect 3674 3706 3677 4086
rect 3682 4013 3685 4126
rect 3698 4116 3701 4316
rect 3706 4173 3709 4343
rect 3714 4253 3717 4326
rect 3722 4213 3725 4236
rect 3738 4196 3741 4326
rect 3754 4323 3757 4373
rect 3770 4346 3773 4406
rect 3766 4343 3773 4346
rect 3766 4256 3769 4343
rect 3766 4253 3773 4256
rect 3746 4213 3757 4216
rect 3762 4213 3765 4236
rect 3738 4193 3749 4196
rect 3770 4193 3773 4253
rect 3698 4113 3705 4116
rect 3690 3936 3693 4106
rect 3702 4036 3705 4113
rect 3698 4033 3705 4036
rect 3698 4013 3701 4033
rect 3706 3983 3709 4006
rect 3714 3993 3717 4016
rect 3722 3943 3725 4006
rect 3738 4003 3741 4126
rect 3746 4076 3749 4193
rect 3778 4146 3781 4336
rect 3786 4306 3789 4476
rect 3818 4473 3829 4476
rect 3818 4403 3821 4473
rect 3834 4413 3837 4446
rect 3794 4326 3797 4386
rect 3834 4383 3837 4406
rect 3874 4363 3877 4416
rect 3882 4403 3885 4416
rect 3890 4353 3893 4556
rect 3930 4533 3933 4596
rect 4002 4573 4005 4606
rect 4026 4573 4029 4606
rect 3898 4413 3901 4446
rect 3938 4386 3941 4406
rect 3930 4383 3941 4386
rect 3794 4323 3805 4326
rect 3786 4303 3793 4306
rect 3790 4156 3793 4303
rect 3802 4213 3805 4256
rect 3810 4196 3813 4206
rect 3818 4203 3821 4216
rect 3826 4196 3829 4216
rect 3834 4203 3837 4346
rect 3858 4313 3861 4326
rect 3882 4323 3885 4336
rect 3898 4333 3901 4366
rect 3930 4326 3933 4383
rect 3946 4333 3949 4416
rect 3954 4403 3957 4416
rect 3898 4313 3901 4326
rect 3930 4323 3941 4326
rect 3842 4213 3845 4246
rect 3874 4203 3877 4216
rect 3882 4213 3885 4236
rect 3810 4193 3829 4196
rect 3890 4183 3893 4226
rect 3898 4166 3901 4206
rect 3890 4163 3901 4166
rect 3790 4153 3805 4156
rect 3762 4133 3765 4146
rect 3778 4143 3789 4146
rect 3746 4073 3757 4076
rect 3754 3996 3757 4073
rect 3746 3993 3757 3996
rect 3778 3993 3781 4016
rect 3690 3933 3697 3936
rect 3658 3703 3677 3706
rect 3650 3543 3653 3606
rect 3658 3583 3661 3703
rect 3682 3693 3685 3926
rect 3694 3856 3697 3933
rect 3706 3913 3709 3936
rect 3714 3903 3717 3926
rect 3690 3853 3697 3856
rect 3690 3626 3693 3853
rect 3698 3796 3701 3836
rect 3706 3813 3709 3876
rect 3722 3833 3725 3936
rect 3730 3923 3733 3936
rect 3746 3933 3749 3993
rect 3786 3976 3789 4143
rect 3794 4013 3797 4126
rect 3802 4076 3805 4153
rect 3802 4073 3813 4076
rect 3810 4006 3813 4073
rect 3778 3973 3789 3976
rect 3802 4003 3813 4006
rect 3698 3793 3705 3796
rect 3702 3716 3705 3793
rect 3714 3786 3717 3806
rect 3722 3793 3725 3816
rect 3730 3803 3733 3916
rect 3738 3873 3741 3926
rect 3778 3896 3781 3973
rect 3802 3903 3805 4003
rect 3818 3933 3821 3946
rect 3778 3893 3789 3896
rect 3746 3793 3749 3806
rect 3754 3786 3757 3816
rect 3714 3783 3725 3786
rect 3714 3733 3717 3746
rect 3722 3733 3725 3783
rect 3746 3783 3757 3786
rect 3702 3713 3709 3716
rect 3686 3623 3693 3626
rect 3666 3513 3669 3526
rect 3674 3523 3677 3606
rect 3650 3333 3653 3456
rect 3634 3323 3645 3326
rect 3634 3236 3637 3323
rect 3626 3233 3637 3236
rect 3618 3143 3621 3206
rect 3626 3196 3629 3233
rect 3626 3193 3637 3196
rect 3618 3053 3621 3126
rect 3586 2733 3593 2736
rect 3590 2606 3593 2733
rect 3586 2603 3593 2606
rect 3586 2583 3589 2603
rect 3586 2523 3589 2536
rect 3594 2533 3597 2566
rect 3570 2503 3573 2516
rect 3570 2413 3597 2416
rect 3570 2403 3573 2413
rect 3570 2316 3573 2396
rect 3578 2323 3581 2406
rect 3586 2323 3589 2356
rect 3570 2313 3581 2316
rect 3562 2293 3569 2296
rect 3566 2196 3569 2293
rect 3578 2213 3581 2313
rect 3594 2233 3597 2406
rect 3602 2393 3605 2746
rect 3618 2733 3621 3016
rect 3626 3003 3629 3136
rect 3634 3133 3637 3193
rect 3626 2906 3629 2996
rect 3634 2923 3637 3086
rect 3626 2903 3633 2906
rect 3630 2826 3633 2903
rect 3626 2823 3633 2826
rect 3626 2743 3629 2823
rect 3634 2773 3637 2806
rect 3642 2783 3645 3286
rect 3650 3123 3653 3326
rect 3658 3283 3661 3476
rect 3686 3456 3689 3623
rect 3706 3616 3709 3713
rect 3698 3613 3709 3616
rect 3730 3613 3733 3726
rect 3746 3703 3749 3783
rect 3754 3726 3757 3736
rect 3754 3723 3765 3726
rect 3754 3623 3757 3723
rect 3686 3453 3693 3456
rect 3690 3433 3693 3453
rect 3682 3393 3685 3406
rect 3666 3203 3669 3346
rect 3674 3323 3677 3356
rect 3690 3306 3693 3336
rect 3682 3303 3693 3306
rect 3682 3226 3685 3303
rect 3682 3223 3693 3226
rect 3658 3156 3661 3176
rect 3658 3153 3665 3156
rect 3650 2966 3653 3096
rect 3662 2996 3665 3153
rect 3674 3093 3677 3126
rect 3682 3123 3685 3206
rect 3690 3106 3693 3223
rect 3698 3133 3701 3613
rect 3786 3596 3789 3893
rect 3826 3856 3829 3986
rect 3834 3923 3837 4006
rect 3842 3933 3845 4126
rect 3850 3933 3853 3996
rect 3866 3993 3869 4146
rect 3890 4066 3893 4163
rect 3906 4153 3909 4266
rect 3938 4213 3941 4323
rect 3962 4233 3965 4566
rect 4106 4563 4109 4616
rect 4194 4613 4197 4626
rect 4146 4556 4149 4606
rect 4122 4553 4149 4556
rect 3978 4413 3981 4526
rect 4018 4456 4021 4546
rect 4002 4453 4021 4456
rect 3978 4256 3981 4366
rect 4002 4356 4005 4453
rect 4026 4413 4029 4446
rect 4034 4403 4037 4426
rect 4042 4403 4045 4526
rect 4098 4513 4101 4526
rect 4002 4353 4021 4356
rect 4018 4333 4021 4353
rect 3978 4253 3985 4256
rect 3982 4176 3985 4253
rect 3994 4213 3997 4326
rect 4026 4186 4029 4376
rect 4042 4323 4045 4396
rect 4026 4183 4045 4186
rect 3978 4173 3985 4176
rect 3890 4063 3897 4066
rect 3894 3966 3897 4063
rect 3858 3933 3861 3966
rect 3890 3963 3897 3966
rect 3802 3813 3805 3836
rect 3810 3813 3813 3856
rect 3822 3853 3829 3856
rect 3822 3766 3825 3853
rect 3842 3813 3845 3836
rect 3810 3763 3825 3766
rect 3810 3676 3813 3763
rect 3802 3673 3813 3676
rect 3802 3626 3805 3673
rect 3834 3666 3837 3726
rect 3842 3713 3845 3796
rect 3818 3663 3837 3666
rect 3802 3623 3813 3626
rect 3706 3523 3709 3536
rect 3714 3533 3717 3596
rect 3770 3593 3789 3596
rect 3706 3203 3709 3436
rect 3714 3346 3717 3526
rect 3730 3456 3733 3536
rect 3738 3526 3741 3586
rect 3738 3523 3757 3526
rect 3746 3476 3749 3496
rect 3722 3453 3733 3456
rect 3742 3473 3749 3476
rect 3722 3366 3725 3453
rect 3742 3366 3745 3473
rect 3722 3363 3733 3366
rect 3742 3363 3749 3366
rect 3714 3343 3721 3346
rect 3718 3246 3721 3343
rect 3714 3243 3721 3246
rect 3714 3153 3717 3243
rect 3730 3226 3733 3363
rect 3746 3343 3749 3363
rect 3754 3336 3757 3523
rect 3762 3413 3765 3506
rect 3770 3493 3773 3593
rect 3778 3533 3781 3546
rect 3786 3533 3789 3556
rect 3794 3433 3797 3536
rect 3802 3513 3805 3526
rect 3810 3496 3813 3623
rect 3818 3613 3821 3663
rect 3842 3636 3845 3696
rect 3834 3633 3845 3636
rect 3806 3493 3813 3496
rect 3806 3426 3809 3493
rect 3806 3423 3813 3426
rect 3786 3356 3789 3416
rect 3722 3223 3733 3226
rect 3746 3333 3757 3336
rect 3778 3353 3789 3356
rect 3686 3103 3693 3106
rect 3686 3026 3689 3103
rect 3658 2993 3665 2996
rect 3674 3023 3689 3026
rect 3658 2973 3661 2993
rect 3650 2963 3661 2966
rect 3650 2923 3653 2946
rect 3650 2736 3653 2826
rect 3658 2813 3661 2963
rect 3674 2946 3677 3023
rect 3682 2953 3685 3016
rect 3698 3013 3701 3106
rect 3714 3093 3717 3126
rect 3690 2993 3693 3006
rect 3706 3003 3709 3016
rect 3714 3013 3717 3086
rect 3722 3033 3725 3223
rect 3746 3213 3749 3333
rect 3778 3316 3781 3353
rect 3786 3333 3789 3346
rect 3770 3313 3781 3316
rect 3770 3206 3773 3313
rect 3794 3213 3797 3336
rect 3802 3323 3805 3406
rect 3810 3363 3813 3423
rect 3810 3313 3813 3356
rect 3818 3256 3821 3576
rect 3826 3563 3829 3616
rect 3826 3503 3829 3526
rect 3834 3486 3837 3633
rect 3842 3613 3845 3626
rect 3850 3576 3853 3856
rect 3858 3646 3861 3926
rect 3866 3793 3869 3926
rect 3890 3876 3893 3963
rect 3890 3873 3901 3876
rect 3898 3853 3901 3873
rect 3890 3766 3893 3806
rect 3882 3763 3893 3766
rect 3882 3733 3885 3763
rect 3898 3733 3901 3756
rect 3898 3713 3901 3726
rect 3906 3696 3909 4146
rect 3914 4013 3917 4126
rect 3930 4116 3933 4136
rect 3930 4113 3941 4116
rect 3938 4066 3941 4113
rect 3978 4073 3981 4173
rect 4002 4133 4005 4146
rect 4026 4133 4029 4166
rect 4042 4133 4045 4183
rect 4050 4166 4053 4336
rect 4058 4313 4061 4456
rect 4074 4333 4077 4406
rect 4082 4353 4085 4416
rect 4098 4413 4101 4506
rect 4106 4333 4109 4416
rect 4114 4363 4117 4406
rect 4122 4373 4125 4553
rect 4138 4513 4141 4526
rect 4146 4503 4149 4536
rect 4162 4533 4165 4546
rect 4194 4536 4197 4546
rect 4186 4533 4197 4536
rect 4162 4523 4173 4526
rect 4130 4413 4133 4436
rect 4138 4403 4141 4456
rect 4162 4413 4165 4516
rect 4170 4416 4173 4523
rect 4178 4423 4181 4526
rect 4170 4413 4181 4416
rect 4098 4303 4101 4326
rect 4050 4163 4061 4166
rect 4058 4146 4061 4163
rect 4058 4143 4069 4146
rect 3986 4123 4013 4126
rect 3930 4063 3941 4066
rect 3914 3776 3917 3936
rect 3922 3923 3925 3936
rect 3930 3923 3933 4063
rect 3946 4006 3949 4016
rect 3954 4013 3957 4046
rect 3938 4003 3949 4006
rect 3938 3866 3941 4003
rect 3946 3933 3949 3956
rect 3954 3916 3957 3936
rect 3954 3913 3961 3916
rect 3922 3863 3941 3866
rect 3922 3803 3925 3863
rect 3914 3773 3925 3776
rect 3898 3693 3909 3696
rect 3858 3643 3869 3646
rect 3858 3593 3861 3606
rect 3830 3483 3837 3486
rect 3830 3426 3833 3483
rect 3806 3253 3821 3256
rect 3826 3423 3833 3426
rect 3806 3206 3809 3253
rect 3730 3203 3741 3206
rect 3770 3203 3781 3206
rect 3730 3163 3733 3203
rect 3730 3056 3733 3156
rect 3738 3076 3741 3186
rect 3778 3173 3781 3203
rect 3802 3203 3809 3206
rect 3802 3136 3805 3203
rect 3826 3166 3829 3423
rect 3834 3213 3837 3416
rect 3842 3376 3845 3576
rect 3850 3573 3857 3576
rect 3854 3496 3857 3573
rect 3866 3553 3869 3643
rect 3882 3576 3885 3636
rect 3890 3603 3893 3626
rect 3882 3573 3889 3576
rect 3866 3513 3869 3536
rect 3874 3523 3877 3566
rect 3886 3516 3889 3573
rect 3882 3513 3889 3516
rect 3854 3493 3861 3496
rect 3842 3373 3849 3376
rect 3846 3286 3849 3373
rect 3842 3283 3849 3286
rect 3842 3183 3845 3283
rect 3858 3266 3861 3493
rect 3850 3263 3861 3266
rect 3850 3196 3853 3263
rect 3850 3193 3861 3196
rect 3826 3163 3837 3166
rect 3762 3093 3765 3136
rect 3778 3103 3781 3136
rect 3794 3133 3805 3136
rect 3738 3073 3749 3076
rect 3730 3053 3737 3056
rect 3722 2993 3725 3016
rect 3734 2996 3737 3053
rect 3730 2993 3737 2996
rect 3730 2976 3733 2993
rect 3722 2973 3733 2976
rect 3674 2943 3685 2946
rect 3666 2823 3669 2926
rect 3674 2886 3677 2936
rect 3682 2916 3685 2943
rect 3698 2933 3701 2946
rect 3682 2913 3701 2916
rect 3674 2883 3685 2886
rect 3682 2826 3685 2883
rect 3674 2823 3685 2826
rect 3610 2693 3613 2726
rect 3626 2706 3629 2726
rect 3622 2703 3629 2706
rect 3622 2636 3625 2703
rect 3622 2633 3629 2636
rect 3626 2613 3629 2633
rect 3634 2606 3637 2736
rect 3642 2733 3653 2736
rect 3642 2713 3645 2733
rect 3658 2706 3661 2806
rect 3666 2793 3669 2816
rect 3674 2803 3677 2823
rect 3698 2796 3701 2913
rect 3722 2816 3725 2973
rect 3746 2966 3749 3073
rect 3794 3066 3797 3133
rect 3794 3063 3801 3066
rect 3738 2963 3749 2966
rect 3722 2813 3733 2816
rect 3682 2793 3701 2796
rect 3730 2793 3733 2813
rect 3650 2703 3661 2706
rect 3650 2616 3653 2703
rect 3618 2603 3637 2606
rect 3642 2613 3653 2616
rect 3610 2523 3613 2536
rect 3618 2533 3621 2603
rect 3642 2566 3645 2613
rect 3666 2606 3669 2756
rect 3682 2723 3685 2793
rect 3722 2646 3725 2726
rect 3714 2643 3725 2646
rect 3714 2613 3717 2643
rect 3666 2603 3677 2606
rect 3638 2563 3645 2566
rect 3610 2473 3613 2516
rect 3626 2493 3629 2526
rect 3638 2496 3641 2563
rect 3638 2493 3645 2496
rect 3642 2476 3645 2493
rect 3610 2403 3613 2416
rect 3602 2333 3621 2336
rect 3626 2333 3629 2346
rect 3602 2316 3605 2333
rect 3634 2323 3637 2476
rect 3642 2473 3649 2476
rect 3646 2336 3649 2473
rect 3642 2333 3649 2336
rect 3602 2313 3613 2316
rect 3610 2236 3613 2313
rect 3642 2306 3645 2333
rect 3602 2233 3613 2236
rect 3634 2303 3645 2306
rect 3566 2193 3573 2196
rect 3570 2106 3573 2193
rect 3586 2143 3589 2226
rect 3602 2216 3605 2233
rect 3594 2213 3605 2216
rect 3602 2133 3605 2206
rect 3610 2203 3613 2216
rect 3634 2166 3637 2303
rect 3650 2286 3653 2316
rect 3646 2283 3653 2286
rect 3646 2226 3649 2283
rect 3658 2273 3661 2596
rect 3674 2556 3677 2603
rect 3670 2553 3677 2556
rect 3670 2406 3673 2553
rect 3722 2543 3725 2616
rect 3730 2536 3733 2746
rect 3682 2413 3685 2526
rect 3666 2403 3673 2406
rect 3666 2383 3669 2403
rect 3666 2333 3685 2336
rect 3666 2323 3669 2333
rect 3666 2266 3669 2296
rect 3674 2286 3677 2326
rect 3690 2303 3693 2496
rect 3706 2483 3709 2536
rect 3722 2533 3733 2536
rect 3722 2506 3725 2533
rect 3718 2503 3725 2506
rect 3698 2323 3701 2406
rect 3706 2323 3709 2456
rect 3718 2346 3721 2503
rect 3714 2343 3721 2346
rect 3674 2283 3693 2286
rect 3666 2263 3673 2266
rect 3646 2223 3653 2226
rect 3634 2163 3645 2166
rect 3610 2133 3613 2146
rect 3618 2143 3637 2146
rect 3562 2103 3573 2106
rect 3538 2083 3549 2086
rect 3514 1993 3525 1996
rect 3514 1893 3517 1936
rect 3522 1903 3525 1993
rect 3530 1876 3533 2016
rect 3546 1966 3549 2083
rect 3522 1873 3533 1876
rect 3538 1963 3549 1966
rect 3474 1463 3477 1616
rect 3458 1453 3465 1456
rect 3406 1313 3413 1316
rect 3418 1343 3429 1346
rect 3442 1343 3445 1406
rect 3450 1343 3453 1446
rect 3462 1356 3465 1453
rect 3458 1353 3465 1356
rect 3406 1256 3409 1313
rect 3418 1256 3421 1343
rect 3458 1333 3461 1353
rect 3406 1253 3413 1256
rect 3418 1253 3429 1256
rect 3410 1233 3413 1253
rect 3394 1223 3405 1226
rect 3374 1043 3381 1046
rect 3354 1013 3357 1026
rect 3330 1003 3341 1006
rect 3314 993 3321 996
rect 3298 873 3309 876
rect 3298 833 3301 873
rect 3318 866 3321 993
rect 3330 883 3333 1003
rect 3362 966 3365 1036
rect 3374 986 3377 1043
rect 3374 983 3381 986
rect 3358 963 3365 966
rect 3378 963 3381 983
rect 3402 973 3405 1223
rect 3418 1133 3421 1166
rect 3426 1046 3429 1253
rect 3434 1116 3437 1326
rect 3442 1123 3445 1216
rect 3474 1146 3477 1456
rect 3482 1393 3485 1536
rect 3490 1533 3493 1556
rect 3498 1536 3501 1576
rect 3506 1543 3509 1726
rect 3498 1533 3509 1536
rect 3490 1523 3501 1526
rect 3514 1523 3517 1536
rect 3490 1483 3493 1523
rect 3490 1376 3493 1466
rect 3486 1373 3493 1376
rect 3486 1246 3489 1373
rect 3498 1266 3501 1516
rect 3506 1273 3509 1416
rect 3514 1413 3517 1436
rect 3522 1326 3525 1873
rect 3538 1856 3541 1963
rect 3562 1956 3565 2103
rect 3578 2013 3581 2026
rect 3570 1993 3573 2006
rect 3594 2003 3597 2126
rect 3618 2123 3621 2143
rect 3626 2036 3629 2136
rect 3634 2133 3637 2143
rect 3642 2123 3645 2163
rect 3650 2123 3653 2223
rect 3658 2056 3661 2236
rect 3670 2166 3673 2263
rect 3690 2213 3693 2283
rect 3706 2246 3709 2306
rect 3714 2293 3717 2343
rect 3730 2303 3733 2526
rect 3738 2496 3741 2963
rect 3746 2923 3749 2936
rect 3754 2903 3757 2926
rect 3746 2686 3749 2806
rect 3762 2803 3765 3036
rect 3798 3006 3801 3063
rect 3810 3013 3813 3126
rect 3818 3123 3821 3146
rect 3834 3106 3837 3163
rect 3858 3143 3861 3193
rect 3874 3136 3877 3376
rect 3882 3333 3885 3513
rect 3898 3496 3901 3693
rect 3914 3626 3917 3766
rect 3922 3633 3925 3773
rect 3938 3763 3941 3806
rect 3946 3766 3949 3906
rect 3958 3826 3961 3913
rect 3954 3823 3961 3826
rect 3954 3803 3957 3823
rect 3946 3763 3957 3766
rect 3906 3613 3909 3626
rect 3914 3623 3925 3626
rect 3914 3593 3917 3616
rect 3922 3576 3925 3623
rect 3918 3573 3925 3576
rect 3894 3493 3901 3496
rect 3894 3436 3897 3493
rect 3906 3446 3909 3526
rect 3918 3506 3921 3573
rect 3930 3513 3933 3756
rect 3938 3743 3957 3746
rect 3938 3723 3941 3743
rect 3946 3723 3949 3736
rect 3954 3733 3957 3743
rect 3946 3613 3949 3626
rect 3918 3503 3925 3506
rect 3906 3443 3913 3446
rect 3894 3433 3901 3436
rect 3890 3343 3893 3416
rect 3898 3316 3901 3433
rect 3890 3313 3901 3316
rect 3890 3246 3893 3313
rect 3910 3306 3913 3443
rect 3906 3303 3913 3306
rect 3890 3243 3897 3246
rect 3858 3116 3861 3136
rect 3874 3133 3885 3136
rect 3826 3103 3837 3106
rect 3850 3113 3861 3116
rect 3826 3083 3829 3103
rect 3850 3046 3853 3113
rect 3850 3043 3861 3046
rect 3798 3003 3805 3006
rect 3770 2876 3773 2926
rect 3786 2923 3789 2936
rect 3802 2916 3805 3003
rect 3842 2956 3845 3006
rect 3858 2986 3861 3043
rect 3866 3003 3869 3126
rect 3882 3026 3885 3133
rect 3874 3023 3885 3026
rect 3834 2953 3845 2956
rect 3850 2983 3861 2986
rect 3834 2923 3837 2953
rect 3794 2913 3805 2916
rect 3770 2873 3777 2876
rect 3774 2796 3777 2873
rect 3794 2816 3797 2913
rect 3770 2793 3777 2796
rect 3786 2813 3797 2816
rect 3770 2733 3773 2793
rect 3786 2743 3789 2813
rect 3746 2683 3753 2686
rect 3750 2536 3753 2683
rect 3770 2616 3773 2726
rect 3786 2643 3789 2726
rect 3770 2613 3777 2616
rect 3746 2533 3753 2536
rect 3746 2513 3749 2533
rect 3762 2516 3765 2606
rect 3774 2536 3777 2613
rect 3794 2593 3797 2806
rect 3802 2793 3805 2806
rect 3810 2796 3813 2816
rect 3818 2803 3821 2816
rect 3834 2813 3837 2836
rect 3826 2796 3829 2806
rect 3810 2793 3829 2796
rect 3802 2716 3805 2736
rect 3802 2713 3813 2716
rect 3810 2636 3813 2713
rect 3802 2633 3813 2636
rect 3802 2613 3805 2633
rect 3826 2626 3829 2766
rect 3842 2743 3845 2906
rect 3850 2726 3853 2983
rect 3874 2946 3877 3023
rect 3894 2976 3897 3243
rect 3894 2973 3901 2976
rect 3874 2943 3881 2946
rect 3858 2813 3861 2926
rect 3842 2723 3853 2726
rect 3858 2723 3861 2736
rect 3842 2646 3845 2723
rect 3842 2643 3853 2646
rect 3826 2623 3837 2626
rect 3810 2593 3813 2606
rect 3818 2573 3821 2616
rect 3834 2566 3837 2623
rect 3850 2613 3853 2643
rect 3858 2613 3861 2706
rect 3866 2596 3869 2936
rect 3878 2776 3881 2943
rect 3890 2793 3893 2806
rect 3898 2803 3901 2973
rect 3906 2823 3909 3303
rect 3922 3286 3925 3503
rect 3938 3413 3941 3496
rect 3918 3283 3925 3286
rect 3918 3196 3921 3283
rect 3930 3203 3933 3406
rect 3946 3396 3949 3566
rect 3954 3556 3957 3726
rect 3962 3723 3965 3806
rect 3962 3563 3965 3646
rect 3970 3593 3973 3996
rect 3986 3913 3989 3926
rect 3978 3746 3981 3766
rect 3978 3743 3985 3746
rect 3982 3666 3985 3743
rect 3994 3716 3997 4123
rect 4066 4096 4069 4143
rect 4074 4123 4077 4216
rect 4090 4166 4093 4236
rect 4086 4163 4093 4166
rect 4106 4166 4109 4226
rect 4114 4213 4117 4326
rect 4122 4306 4125 4336
rect 4130 4323 4133 4356
rect 4146 4343 4149 4406
rect 4170 4376 4173 4406
rect 4154 4373 4173 4376
rect 4138 4323 4141 4336
rect 4154 4333 4157 4373
rect 4178 4336 4181 4413
rect 4186 4343 4189 4533
rect 4194 4433 4197 4526
rect 4202 4513 4205 4536
rect 4210 4456 4213 4606
rect 4226 4533 4229 4616
rect 4234 4613 4237 4626
rect 4306 4613 4309 4636
rect 4206 4453 4213 4456
rect 4206 4376 4209 4453
rect 4226 4413 4229 4526
rect 4206 4373 4213 4376
rect 4122 4303 4129 4306
rect 4126 4226 4129 4303
rect 4138 4236 4141 4316
rect 4138 4233 4145 4236
rect 4126 4223 4133 4226
rect 4106 4163 4113 4166
rect 4086 4106 4089 4163
rect 4110 4106 4113 4163
rect 4130 4126 4133 4223
rect 4142 4156 4145 4233
rect 4122 4123 4133 4126
rect 4138 4153 4145 4156
rect 4086 4103 4093 4106
rect 4110 4103 4117 4106
rect 4058 4093 4069 4096
rect 4002 3933 4005 3946
rect 4010 3943 4029 3946
rect 4010 3923 4013 3943
rect 4018 3923 4021 3936
rect 4026 3933 4029 3943
rect 4034 3926 4037 4006
rect 4042 3943 4045 4016
rect 4058 3993 4061 4093
rect 4090 4086 4093 4103
rect 4090 4083 4101 4086
rect 4098 3966 4101 4083
rect 4114 4036 4117 4103
rect 4138 4063 4141 4153
rect 4146 4043 4149 4136
rect 4090 3963 4101 3966
rect 4106 4033 4117 4036
rect 4154 4036 4157 4326
rect 4170 4266 4173 4336
rect 4178 4333 4189 4336
rect 4178 4313 4181 4326
rect 4170 4263 4177 4266
rect 4162 4213 4165 4256
rect 4162 4133 4165 4206
rect 4174 4176 4177 4263
rect 4186 4253 4189 4333
rect 4194 4223 4197 4326
rect 4170 4173 4177 4176
rect 4170 4153 4173 4173
rect 4170 4133 4173 4146
rect 4178 4113 4181 4126
rect 4186 4123 4189 4206
rect 4194 4143 4197 4216
rect 4202 4193 4205 4346
rect 4210 4183 4213 4373
rect 4234 4353 4237 4526
rect 4242 4333 4245 4536
rect 4250 4523 4253 4606
rect 4282 4573 4285 4606
rect 4362 4603 4365 4616
rect 4258 4446 4261 4536
rect 4266 4533 4269 4546
rect 4266 4453 4269 4526
rect 4274 4503 4277 4526
rect 4282 4476 4285 4556
rect 4298 4533 4301 4556
rect 4274 4473 4285 4476
rect 4250 4443 4261 4446
rect 4250 4413 4253 4443
rect 4274 4306 4277 4473
rect 4298 4436 4301 4526
rect 4298 4433 4309 4436
rect 4306 4386 4309 4433
rect 4298 4383 4309 4386
rect 4298 4333 4301 4383
rect 4306 4313 4309 4326
rect 4266 4303 4277 4306
rect 4266 4246 4269 4303
rect 4262 4243 4269 4246
rect 4226 4163 4229 4206
rect 4262 4186 4265 4243
rect 4274 4213 4277 4236
rect 4178 4046 4181 4066
rect 4178 4043 4185 4046
rect 4154 4033 4173 4036
rect 4002 3733 4005 3776
rect 4026 3763 4029 3926
rect 4034 3923 4045 3926
rect 4042 3856 4045 3923
rect 4034 3853 4045 3856
rect 4034 3746 4037 3853
rect 4090 3846 4093 3963
rect 4106 3856 4109 4033
rect 4114 3923 4117 4016
rect 4146 3993 4149 4016
rect 4162 4013 4165 4026
rect 4170 3976 4173 4033
rect 4162 3973 4173 3976
rect 4154 3933 4157 3946
rect 4106 3853 4117 3856
rect 4090 3843 4101 3846
rect 4026 3743 4037 3746
rect 3994 3713 4005 3716
rect 3978 3663 3985 3666
rect 3978 3643 3981 3663
rect 4002 3636 4005 3713
rect 4026 3696 4029 3743
rect 4042 3723 4045 3816
rect 4074 3793 4077 3806
rect 4050 3703 4053 3726
rect 4058 3713 4061 3736
rect 4066 3723 4069 3776
rect 4090 3773 4093 3806
rect 4074 3733 4077 3756
rect 4082 3706 4085 3766
rect 4098 3733 4101 3843
rect 4074 3703 4085 3706
rect 4026 3693 4037 3696
rect 4034 3636 4037 3693
rect 4002 3633 4013 3636
rect 3954 3553 3973 3556
rect 3962 3533 3965 3546
rect 3954 3423 3957 3526
rect 3942 3393 3949 3396
rect 3954 3393 3957 3416
rect 3942 3286 3945 3393
rect 3962 3353 3965 3516
rect 3970 3493 3973 3553
rect 3970 3403 3973 3486
rect 3978 3393 3981 3406
rect 3942 3283 3949 3286
rect 3918 3193 3925 3196
rect 3922 3146 3925 3193
rect 3918 3143 3925 3146
rect 3918 3036 3921 3143
rect 3946 3136 3949 3283
rect 3954 3153 3957 3206
rect 3930 3133 3949 3136
rect 3930 3043 3933 3133
rect 3918 3033 3925 3036
rect 3914 2813 3917 2926
rect 3878 2773 3893 2776
rect 3890 2733 3893 2773
rect 3922 2733 3925 3033
rect 3938 3013 3941 3126
rect 3954 3086 3957 3146
rect 3962 3143 3965 3336
rect 3970 3306 3973 3386
rect 3986 3323 3989 3416
rect 3994 3413 3997 3606
rect 4010 3383 4013 3633
rect 4026 3633 4037 3636
rect 3970 3303 3981 3306
rect 3978 3236 3981 3303
rect 4002 3266 4005 3286
rect 3970 3233 3981 3236
rect 3994 3263 4005 3266
rect 3970 3186 3973 3233
rect 3978 3203 3981 3216
rect 3970 3183 3981 3186
rect 3950 3083 3957 3086
rect 3950 3006 3953 3083
rect 3946 3003 3953 3006
rect 3946 2933 3949 3003
rect 3962 2933 3965 3136
rect 3978 2986 3981 3183
rect 3994 3166 3997 3263
rect 3994 3163 4005 3166
rect 3994 3076 3997 3146
rect 4002 3123 4005 3163
rect 4010 3143 4013 3366
rect 4026 3356 4029 3633
rect 4074 3606 4077 3703
rect 4090 3613 4093 3726
rect 4042 3593 4045 3606
rect 4074 3603 4085 3606
rect 4058 3536 4061 3586
rect 4082 3546 4085 3603
rect 4106 3576 4109 3796
rect 4114 3786 4117 3853
rect 4114 3783 4121 3786
rect 4118 3576 4121 3783
rect 4054 3533 4061 3536
rect 4074 3543 4085 3546
rect 4098 3573 4109 3576
rect 4114 3573 4121 3576
rect 4034 3403 4037 3426
rect 4054 3406 4057 3533
rect 4066 3413 4069 3526
rect 4074 3476 4077 3543
rect 4074 3473 4085 3476
rect 4082 3406 4085 3473
rect 4098 3466 4101 3573
rect 4114 3553 4117 3573
rect 4130 3556 4133 3926
rect 4162 3883 4165 3973
rect 4182 3956 4185 4043
rect 4178 3953 4185 3956
rect 4170 3826 4173 3936
rect 4126 3553 4133 3556
rect 4114 3523 4117 3536
rect 4114 3473 4117 3516
rect 4098 3463 4109 3466
rect 4026 3353 4033 3356
rect 4030 3306 4033 3353
rect 4026 3303 4033 3306
rect 4026 3283 4029 3303
rect 4026 3203 4029 3226
rect 4018 3113 4021 3126
rect 4034 3123 4037 3206
rect 4042 3196 4045 3406
rect 4054 3403 4061 3406
rect 4050 3213 4053 3226
rect 4042 3193 4049 3196
rect 4058 3193 4061 3403
rect 4074 3403 4085 3406
rect 4046 3116 4049 3193
rect 4074 3156 4077 3403
rect 4106 3373 4109 3463
rect 4126 3456 4129 3553
rect 4126 3453 4133 3456
rect 4082 3333 4085 3346
rect 4090 3343 4109 3346
rect 4130 3343 4133 3453
rect 4090 3323 4093 3343
rect 4098 3256 4101 3336
rect 4106 3333 4109 3343
rect 4130 3313 4133 3326
rect 4138 3296 4141 3806
rect 4146 3803 4149 3816
rect 4154 3813 4157 3826
rect 4162 3823 4173 3826
rect 4162 3746 4165 3823
rect 4146 3743 4165 3746
rect 4170 3743 4173 3816
rect 4146 3696 4149 3743
rect 4154 3713 4157 3726
rect 4162 3723 4165 3736
rect 4170 3706 4173 3736
rect 4166 3703 4173 3706
rect 4146 3693 4153 3696
rect 4150 3576 4153 3693
rect 4166 3636 4169 3703
rect 4166 3633 4173 3636
rect 4162 3593 4165 3616
rect 4146 3573 4153 3576
rect 4146 3383 4149 3573
rect 4170 3556 4173 3633
rect 4178 3573 4181 3953
rect 4186 3896 4189 3936
rect 4194 3933 4197 4016
rect 4202 3993 4205 4156
rect 4242 4146 4245 4186
rect 4262 4183 4269 4186
rect 4234 4143 4245 4146
rect 4218 4113 4221 4126
rect 4234 4096 4237 4143
rect 4266 4133 4269 4183
rect 4290 4156 4293 4266
rect 4314 4246 4317 4336
rect 4330 4333 4333 4406
rect 4338 4333 4341 4416
rect 4346 4413 4349 4526
rect 4378 4413 4381 4526
rect 4386 4523 4389 4616
rect 4442 4556 4445 4616
rect 4442 4553 4453 4556
rect 4466 4553 4469 4606
rect 4426 4543 4445 4546
rect 4394 4413 4397 4526
rect 4426 4523 4429 4543
rect 4434 4506 4437 4536
rect 4442 4533 4445 4543
rect 4426 4503 4437 4506
rect 4426 4436 4429 4503
rect 4442 4486 4445 4526
rect 4450 4523 4453 4553
rect 4474 4523 4485 4526
rect 4442 4483 4453 4486
rect 4426 4433 4437 4436
rect 4322 4263 4325 4326
rect 4338 4313 4341 4326
rect 4314 4243 4325 4246
rect 4298 4213 4309 4216
rect 4314 4213 4317 4236
rect 4286 4153 4293 4156
rect 4286 4106 4289 4153
rect 4306 4133 4309 4166
rect 4322 4143 4325 4243
rect 4286 4103 4293 4106
rect 4234 4093 4245 4096
rect 4242 4056 4245 4093
rect 4238 4053 4245 4056
rect 4218 4016 4221 4046
rect 4218 4013 4229 4016
rect 4210 3933 4213 4006
rect 4226 3966 4229 4013
rect 4238 3996 4241 4053
rect 4290 4046 4293 4103
rect 4266 4043 4293 4046
rect 4238 3993 4245 3996
rect 4242 3976 4245 3993
rect 4242 3973 4253 3976
rect 4218 3963 4229 3966
rect 4194 3913 4197 3926
rect 4186 3893 4197 3896
rect 4194 3846 4197 3893
rect 4186 3843 4197 3846
rect 4186 3823 4189 3843
rect 4186 3613 4189 3726
rect 4202 3723 4205 3806
rect 4210 3716 4213 3926
rect 4218 3906 4221 3963
rect 4226 3943 4245 3946
rect 4226 3923 4229 3943
rect 4234 3923 4237 3936
rect 4242 3933 4245 3943
rect 4250 3926 4253 3973
rect 4266 3956 4269 4043
rect 4266 3953 4277 3956
rect 4242 3923 4253 3926
rect 4218 3903 4229 3906
rect 4226 3816 4229 3903
rect 4242 3833 4245 3923
rect 4266 3906 4269 3936
rect 4258 3903 4269 3906
rect 4218 3813 4229 3816
rect 4218 3793 4221 3813
rect 4258 3766 4261 3903
rect 4258 3763 4269 3766
rect 4202 3713 4213 3716
rect 4202 3613 4205 3713
rect 4154 3553 4173 3556
rect 4154 3523 4157 3553
rect 4162 3533 4165 3546
rect 4170 3543 4189 3546
rect 4170 3523 4173 3543
rect 4154 3413 4157 3506
rect 4178 3456 4181 3536
rect 4186 3533 4189 3543
rect 4194 3536 4197 3606
rect 4194 3533 4205 3536
rect 4186 3493 4189 3526
rect 4194 3503 4197 3526
rect 4178 3453 4189 3456
rect 4186 3393 4189 3453
rect 4202 3403 4205 3533
rect 4218 3363 4221 3726
rect 4250 3723 4253 3746
rect 4250 3613 4253 3716
rect 4266 3656 4269 3763
rect 4274 3733 4277 3953
rect 4282 3923 4285 4016
rect 4306 4003 4309 4016
rect 4298 3906 4301 3976
rect 4290 3903 4301 3906
rect 4290 3836 4293 3903
rect 4290 3833 4301 3836
rect 4282 3766 4285 3806
rect 4290 3783 4293 3816
rect 4282 3763 4289 3766
rect 4274 3713 4277 3726
rect 4286 3706 4289 3763
rect 4262 3653 4269 3656
rect 4282 3703 4289 3706
rect 4262 3576 4265 3653
rect 4262 3573 4269 3576
rect 4234 3506 4237 3556
rect 4258 3523 4261 3536
rect 4266 3506 4269 3573
rect 4234 3503 4245 3506
rect 4242 3446 4245 3503
rect 4234 3443 4245 3446
rect 4258 3503 4269 3506
rect 4090 3253 4101 3256
rect 4130 3293 4141 3296
rect 4090 3213 4093 3253
rect 4130 3206 4133 3293
rect 4146 3213 4149 3326
rect 4130 3203 4141 3206
rect 4042 3113 4049 3116
rect 4058 3153 4077 3156
rect 4042 3096 4045 3113
rect 4034 3093 4045 3096
rect 3994 3073 4013 3076
rect 3970 2983 3981 2986
rect 3930 2796 3933 2816
rect 3962 2813 3965 2926
rect 3970 2796 3973 2983
rect 3978 2946 3981 2966
rect 3978 2943 3985 2946
rect 3982 2826 3985 2943
rect 3930 2793 3937 2796
rect 3874 2703 3877 2726
rect 3914 2703 3917 2726
rect 3826 2563 3837 2566
rect 3850 2593 3869 2596
rect 3758 2513 3765 2516
rect 3770 2533 3777 2536
rect 3738 2493 3749 2496
rect 3746 2356 3749 2493
rect 3758 2436 3761 2513
rect 3758 2433 3765 2436
rect 3762 2413 3765 2433
rect 3742 2353 3749 2356
rect 3742 2296 3745 2353
rect 3738 2293 3745 2296
rect 3702 2243 3709 2246
rect 3702 2166 3705 2243
rect 3670 2163 3677 2166
rect 3674 2116 3677 2163
rect 3666 2113 3677 2116
rect 3690 2163 3705 2166
rect 3666 2093 3669 2113
rect 3658 2053 3665 2056
rect 3626 2033 3637 2036
rect 3618 2013 3621 2026
rect 3562 1953 3573 1956
rect 3534 1853 3541 1856
rect 3534 1746 3537 1853
rect 3546 1756 3549 1946
rect 3554 1913 3557 1926
rect 3570 1836 3573 1953
rect 3602 1933 3605 1966
rect 3610 1933 3613 1946
rect 3562 1833 3573 1836
rect 3562 1776 3565 1833
rect 3570 1796 3573 1816
rect 3578 1803 3581 1816
rect 3586 1796 3589 1806
rect 3570 1793 3589 1796
rect 3594 1776 3597 1816
rect 3562 1773 3573 1776
rect 3546 1753 3557 1756
rect 3534 1743 3541 1746
rect 3538 1686 3541 1743
rect 3534 1683 3541 1686
rect 3534 1636 3537 1683
rect 3554 1676 3557 1753
rect 3546 1673 3557 1676
rect 3534 1633 3541 1636
rect 3530 1523 3533 1606
rect 3538 1566 3541 1633
rect 3546 1583 3549 1673
rect 3570 1656 3573 1773
rect 3586 1773 3597 1776
rect 3586 1716 3589 1773
rect 3602 1723 3605 1926
rect 3618 1923 3621 1996
rect 3634 1986 3637 2033
rect 3626 1983 3637 1986
rect 3626 1963 3629 1983
rect 3634 1906 3637 1926
rect 3626 1903 3637 1906
rect 3626 1836 3629 1903
rect 3626 1833 3637 1836
rect 3610 1723 3613 1816
rect 3634 1813 3637 1833
rect 3642 1796 3645 1926
rect 3634 1793 3645 1796
rect 3586 1713 3597 1716
rect 3562 1653 3573 1656
rect 3562 1636 3565 1653
rect 3594 1636 3597 1713
rect 3558 1633 3565 1636
rect 3578 1633 3597 1636
rect 3538 1563 3545 1566
rect 3542 1516 3545 1563
rect 3558 1546 3561 1633
rect 3558 1543 3565 1546
rect 3538 1513 3545 1516
rect 3538 1453 3541 1513
rect 3554 1496 3557 1526
rect 3562 1503 3565 1543
rect 3550 1493 3557 1496
rect 3550 1436 3553 1493
rect 3570 1466 3573 1616
rect 3578 1613 3581 1633
rect 3594 1613 3605 1616
rect 3610 1613 3613 1636
rect 3578 1533 3581 1606
rect 3562 1463 3573 1466
rect 3550 1433 3557 1436
rect 3554 1416 3557 1433
rect 3546 1413 3557 1416
rect 3562 1413 3565 1463
rect 3578 1423 3581 1526
rect 3586 1513 3589 1526
rect 3594 1523 3605 1526
rect 3586 1486 3589 1506
rect 3586 1483 3597 1486
rect 3594 1406 3597 1483
rect 3538 1383 3541 1406
rect 3554 1393 3557 1406
rect 3562 1403 3597 1406
rect 3530 1333 3533 1346
rect 3514 1323 3525 1326
rect 3498 1263 3509 1266
rect 3486 1243 3493 1246
rect 3474 1143 3485 1146
rect 3434 1113 3445 1116
rect 3426 1043 3437 1046
rect 3418 966 3421 1006
rect 3402 963 3421 966
rect 3338 913 3341 926
rect 3346 923 3349 946
rect 3358 916 3361 963
rect 3358 913 3365 916
rect 3386 913 3389 926
rect 3362 893 3365 913
rect 3318 863 3325 866
rect 3282 783 3285 816
rect 3322 786 3325 863
rect 3314 783 3325 786
rect 3290 603 3293 626
rect 3298 583 3301 686
rect 3290 513 3293 526
rect 3298 466 3301 536
rect 3290 463 3301 466
rect 3266 413 3285 416
rect 3266 363 3269 406
rect 3274 396 3277 406
rect 3290 403 3293 463
rect 3306 456 3309 766
rect 3298 453 3309 456
rect 3298 396 3301 453
rect 3274 393 3301 396
rect 3210 343 3229 346
rect 3210 323 3213 343
rect 3218 313 3221 336
rect 3226 333 3229 343
rect 3186 213 3189 236
rect 3074 123 3077 196
rect 3194 193 3197 206
rect 3202 186 3205 216
rect 3226 213 3229 326
rect 3266 313 3269 326
rect 3282 296 3285 336
rect 3306 313 3309 326
rect 3274 293 3285 296
rect 3202 183 3213 186
rect 3122 133 3125 176
rect 3170 113 3173 126
rect 3202 123 3205 176
rect 3210 133 3213 183
rect 3218 173 3221 206
rect 3234 203 3237 216
rect 3242 133 3245 216
rect 3258 213 3261 246
rect 3274 226 3277 293
rect 3266 223 3277 226
rect 3250 193 3253 206
rect 3258 173 3261 206
rect 3266 133 3269 223
rect 3274 203 3277 216
rect 3290 213 3293 286
rect 3314 283 3317 783
rect 3330 733 3333 766
rect 3338 756 3341 816
rect 3338 753 3357 756
rect 3338 733 3349 736
rect 3322 683 3325 726
rect 3330 703 3333 726
rect 3354 723 3357 753
rect 3362 706 3365 856
rect 3354 703 3365 706
rect 3354 636 3357 703
rect 3378 693 3381 876
rect 3386 766 3389 896
rect 3394 776 3397 946
rect 3402 783 3405 963
rect 3426 943 3429 1026
rect 3434 983 3437 1043
rect 3442 1003 3445 1113
rect 3418 866 3421 886
rect 3414 863 3421 866
rect 3414 796 3417 863
rect 3426 853 3429 936
rect 3442 923 3445 976
rect 3450 896 3453 1116
rect 3458 1023 3461 1126
rect 3466 1123 3469 1136
rect 3474 1056 3477 1136
rect 3466 1053 3477 1056
rect 3458 993 3461 1006
rect 3466 943 3469 1053
rect 3482 1036 3485 1143
rect 3490 1133 3493 1243
rect 3498 1203 3501 1256
rect 3506 1213 3509 1263
rect 3514 1206 3517 1323
rect 3530 1306 3533 1326
rect 3530 1303 3541 1306
rect 3506 1203 3517 1206
rect 3498 1113 3501 1126
rect 3506 1096 3509 1203
rect 3522 1133 3525 1276
rect 3538 1256 3541 1303
rect 3530 1253 3541 1256
rect 3562 1253 3565 1403
rect 3610 1383 3613 1606
rect 3634 1576 3637 1793
rect 3650 1776 3653 1976
rect 3646 1773 3653 1776
rect 3646 1656 3649 1773
rect 3662 1766 3665 2053
rect 3690 2036 3693 2163
rect 3714 2046 3717 2236
rect 3738 2233 3741 2293
rect 3754 2223 3757 2336
rect 3738 2193 3741 2206
rect 3762 2203 3765 2236
rect 3722 2113 3725 2126
rect 3730 2103 3733 2126
rect 3762 2113 3765 2126
rect 3770 2086 3773 2533
rect 3778 2436 3781 2516
rect 3786 2453 3789 2546
rect 3794 2543 3813 2546
rect 3794 2523 3797 2543
rect 3778 2433 3789 2436
rect 3786 2246 3789 2433
rect 3802 2423 3805 2536
rect 3810 2533 3813 2543
rect 3810 2473 3813 2526
rect 3810 2413 3813 2466
rect 3826 2413 3829 2563
rect 3850 2446 3853 2593
rect 3850 2443 3865 2446
rect 3834 2413 3837 2426
rect 3802 2353 3805 2406
rect 3842 2393 3845 2406
rect 3778 2243 3789 2246
rect 3778 2206 3781 2243
rect 3802 2233 3805 2326
rect 3818 2313 3821 2326
rect 3826 2323 3829 2336
rect 3834 2333 3837 2356
rect 3786 2213 3789 2226
rect 3826 2213 3829 2226
rect 3778 2203 3789 2206
rect 3786 2146 3789 2203
rect 3802 2176 3805 2206
rect 3802 2173 3813 2176
rect 3782 2143 3789 2146
rect 3782 2096 3785 2143
rect 3810 2133 3813 2173
rect 3834 2136 3837 2326
rect 3850 2256 3853 2406
rect 3862 2376 3865 2443
rect 3874 2383 3877 2616
rect 3882 2533 3885 2546
rect 3862 2373 3869 2376
rect 3846 2253 3853 2256
rect 3866 2256 3869 2373
rect 3890 2333 3893 2606
rect 3898 2406 3901 2626
rect 3922 2613 3925 2726
rect 3934 2646 3937 2793
rect 3930 2643 3937 2646
rect 3962 2793 3973 2796
rect 3978 2823 3985 2826
rect 3930 2623 3933 2643
rect 3914 2533 3917 2606
rect 3930 2536 3933 2616
rect 3938 2593 3941 2606
rect 3946 2586 3949 2616
rect 3962 2606 3965 2793
rect 3978 2733 3981 2823
rect 3994 2813 3997 2826
rect 3986 2793 3989 2806
rect 4002 2776 4005 2816
rect 3994 2773 4005 2776
rect 3978 2613 3981 2726
rect 3962 2603 3973 2606
rect 3922 2533 3933 2536
rect 3938 2583 3949 2586
rect 3906 2413 3909 2526
rect 3914 2503 3917 2526
rect 3922 2486 3925 2533
rect 3938 2513 3941 2583
rect 3970 2556 3973 2603
rect 3970 2553 3981 2556
rect 3946 2543 3965 2546
rect 3946 2523 3949 2543
rect 3914 2483 3925 2486
rect 3898 2403 3909 2406
rect 3890 2306 3893 2326
rect 3886 2303 3893 2306
rect 3866 2253 3877 2256
rect 3846 2196 3849 2253
rect 3846 2193 3853 2196
rect 3850 2176 3853 2193
rect 3850 2173 3861 2176
rect 3830 2133 3837 2136
rect 3782 2093 3789 2096
rect 3754 2083 3773 2086
rect 3714 2043 3725 2046
rect 3690 2033 3709 2036
rect 3674 1916 3677 2016
rect 3706 1973 3709 2033
rect 3722 1976 3725 2043
rect 3754 2013 3757 2083
rect 3770 2013 3773 2056
rect 3786 2013 3789 2093
rect 3830 2076 3833 2133
rect 3818 2073 3833 2076
rect 3714 1973 3725 1976
rect 3682 1933 3685 1956
rect 3714 1923 3717 1973
rect 3730 1943 3733 1956
rect 3746 1926 3749 1946
rect 3742 1923 3749 1926
rect 3674 1913 3685 1916
rect 3682 1846 3685 1913
rect 3674 1843 3685 1846
rect 3674 1813 3677 1843
rect 3658 1763 3665 1766
rect 3658 1663 3661 1763
rect 3682 1723 3685 1816
rect 3690 1813 3693 1826
rect 3690 1776 3693 1796
rect 3690 1773 3697 1776
rect 3694 1716 3697 1773
rect 3690 1713 3697 1716
rect 3646 1653 3653 1656
rect 3634 1573 3641 1576
rect 3626 1513 3629 1526
rect 3638 1446 3641 1573
rect 3638 1443 3645 1446
rect 3634 1413 3637 1426
rect 3642 1366 3645 1443
rect 3650 1433 3653 1653
rect 3674 1636 3677 1686
rect 3666 1633 3677 1636
rect 3666 1586 3669 1633
rect 3690 1603 3693 1713
rect 3706 1646 3709 1806
rect 3714 1803 3717 1816
rect 3730 1813 3733 1856
rect 3742 1826 3745 1923
rect 3742 1823 3749 1826
rect 3746 1803 3749 1823
rect 3754 1813 3757 1986
rect 3762 1933 3765 2006
rect 3818 1946 3821 2073
rect 3818 1943 3837 1946
rect 3818 1846 3821 1926
rect 3826 1863 3829 1926
rect 3818 1843 3825 1846
rect 3762 1793 3765 1806
rect 3786 1753 3789 1806
rect 3730 1683 3733 1736
rect 3802 1713 3805 1736
rect 3810 1723 3813 1816
rect 3822 1746 3825 1843
rect 3818 1743 3825 1746
rect 3706 1643 3717 1646
rect 3714 1606 3717 1643
rect 3714 1603 3725 1606
rect 3666 1583 3677 1586
rect 3674 1496 3677 1583
rect 3690 1543 3693 1556
rect 3698 1533 3701 1566
rect 3706 1516 3709 1586
rect 3698 1513 3709 1516
rect 3674 1493 3685 1496
rect 3682 1393 3685 1493
rect 3698 1446 3701 1513
rect 3698 1443 3709 1446
rect 3698 1383 3701 1406
rect 3706 1376 3709 1443
rect 3714 1403 3717 1596
rect 3626 1363 3645 1366
rect 3682 1373 3709 1376
rect 3578 1313 3581 1326
rect 3530 1203 3533 1253
rect 3586 1236 3589 1326
rect 3546 1173 3549 1216
rect 3530 1133 3533 1146
rect 3538 1133 3541 1156
rect 3478 1033 3485 1036
rect 3502 1093 3509 1096
rect 3478 976 3481 1033
rect 3478 973 3485 976
rect 3442 893 3453 896
rect 3442 806 3445 893
rect 3458 813 3461 926
rect 3442 803 3461 806
rect 3482 803 3485 973
rect 3502 946 3505 1093
rect 3514 1086 3517 1126
rect 3538 1123 3549 1126
rect 3514 1083 3525 1086
rect 3514 996 3517 1083
rect 3522 1013 3525 1026
rect 3546 1003 3549 1106
rect 3554 1033 3557 1236
rect 3578 1233 3589 1236
rect 3562 1193 3565 1206
rect 3570 1203 3573 1216
rect 3562 1133 3565 1176
rect 3578 1163 3581 1233
rect 3586 1203 3597 1206
rect 3562 1013 3565 1026
rect 3570 1006 3573 1136
rect 3578 1123 3581 1136
rect 3586 1113 3589 1126
rect 3562 1003 3573 1006
rect 3514 993 3533 996
rect 3498 943 3505 946
rect 3498 866 3501 943
rect 3498 863 3509 866
rect 3498 813 3501 846
rect 3414 793 3421 796
rect 3394 773 3413 776
rect 3386 763 3397 766
rect 3394 733 3397 763
rect 3402 656 3405 766
rect 3410 723 3413 773
rect 3418 733 3421 793
rect 3378 653 3405 656
rect 3354 633 3365 636
rect 3322 613 3325 626
rect 3330 603 3333 616
rect 3330 513 3333 526
rect 3338 443 3341 606
rect 3346 586 3349 616
rect 3346 583 3353 586
rect 3350 436 3353 583
rect 3362 566 3365 633
rect 3370 613 3373 626
rect 3378 613 3381 653
rect 3426 623 3429 726
rect 3442 696 3445 726
rect 3450 723 3453 736
rect 3458 703 3461 803
rect 3498 783 3501 806
rect 3466 723 3469 756
rect 3482 733 3485 746
rect 3482 706 3485 726
rect 3474 703 3485 706
rect 3434 693 3445 696
rect 3434 613 3437 693
rect 3474 646 3477 703
rect 3474 643 3485 646
rect 3362 563 3381 566
rect 3378 483 3381 563
rect 3418 533 3421 546
rect 3346 433 3353 436
rect 3322 413 3325 426
rect 3346 366 3349 433
rect 3362 383 3365 416
rect 3346 363 3353 366
rect 3282 183 3285 206
rect 3306 193 3309 206
rect 3314 143 3317 216
rect 3322 203 3325 296
rect 3330 203 3333 336
rect 3338 213 3341 286
rect 3350 276 3353 363
rect 3362 303 3365 326
rect 3370 323 3373 346
rect 3346 273 3353 276
rect 3346 253 3349 273
rect 3362 213 3365 226
rect 3346 183 3349 206
rect 3354 193 3357 206
rect 3210 113 3213 126
rect 3250 113 3253 126
rect 3290 113 3293 126
rect 3346 123 3349 146
rect 3370 123 3373 206
rect 3378 196 3381 216
rect 3386 203 3389 406
rect 3394 396 3397 416
rect 3402 403 3405 526
rect 3410 416 3413 426
rect 3410 413 3421 416
rect 3442 413 3445 426
rect 3450 413 3453 436
rect 3410 396 3413 406
rect 3394 393 3413 396
rect 3394 343 3413 346
rect 3394 323 3397 343
rect 3402 323 3405 336
rect 3410 333 3413 343
rect 3394 216 3397 236
rect 3394 213 3405 216
rect 3394 196 3397 206
rect 3402 203 3405 213
rect 3378 193 3397 196
rect 3410 123 3413 216
rect 3418 213 3421 413
rect 3458 333 3461 616
rect 3474 566 3477 616
rect 3466 563 3477 566
rect 3466 523 3469 563
rect 3482 533 3485 643
rect 3490 586 3493 736
rect 3506 733 3509 863
rect 3514 813 3517 936
rect 3522 933 3525 946
rect 3522 843 3525 926
rect 3530 923 3533 993
rect 3522 803 3525 836
rect 3530 813 3533 826
rect 3514 686 3517 726
rect 3506 683 3517 686
rect 3506 616 3509 683
rect 3506 613 3517 616
rect 3522 613 3525 776
rect 3530 763 3533 806
rect 3498 586 3501 596
rect 3490 583 3501 586
rect 3498 523 3501 583
rect 3514 573 3517 613
rect 3522 596 3525 606
rect 3530 603 3533 756
rect 3538 633 3541 816
rect 3538 596 3541 616
rect 3522 593 3541 596
rect 3546 586 3549 986
rect 3554 773 3557 846
rect 3554 703 3557 736
rect 3562 733 3565 1003
rect 3578 986 3581 1036
rect 3586 1013 3589 1056
rect 3594 1046 3597 1146
rect 3602 1053 3605 1216
rect 3626 1176 3629 1363
rect 3674 1306 3677 1326
rect 3666 1303 3677 1306
rect 3666 1236 3669 1303
rect 3666 1233 3677 1236
rect 3650 1213 3661 1216
rect 3674 1213 3677 1233
rect 3682 1213 3685 1373
rect 3706 1333 3709 1346
rect 3722 1296 3725 1603
rect 3730 1516 3733 1666
rect 3738 1533 3741 1616
rect 3762 1533 3765 1566
rect 3778 1563 3781 1616
rect 3786 1583 3789 1616
rect 3794 1603 3797 1696
rect 3818 1626 3821 1743
rect 3826 1703 3829 1726
rect 3802 1623 3821 1626
rect 3778 1533 3781 1556
rect 3730 1513 3741 1516
rect 3754 1513 3757 1526
rect 3762 1523 3773 1526
rect 3786 1523 3789 1576
rect 3802 1546 3805 1623
rect 3802 1543 3821 1546
rect 3738 1436 3741 1513
rect 3762 1483 3765 1523
rect 3734 1433 3741 1436
rect 3734 1356 3737 1433
rect 3746 1396 3749 1416
rect 3754 1403 3757 1436
rect 3762 1413 3765 1466
rect 3770 1436 3773 1456
rect 3770 1433 3777 1436
rect 3762 1396 3765 1406
rect 3746 1393 3765 1396
rect 3774 1386 3777 1433
rect 3714 1293 3725 1296
rect 3730 1353 3737 1356
rect 3770 1383 3777 1386
rect 3730 1336 3733 1353
rect 3730 1333 3741 1336
rect 3698 1226 3701 1286
rect 3714 1246 3717 1293
rect 3714 1243 3725 1246
rect 3694 1223 3701 1226
rect 3722 1223 3725 1243
rect 3626 1173 3645 1176
rect 3594 1043 3605 1046
rect 3574 983 3581 986
rect 3574 916 3577 983
rect 3586 923 3589 1006
rect 3602 1003 3605 1043
rect 3610 1013 3613 1126
rect 3626 1113 3629 1126
rect 3642 1093 3645 1173
rect 3650 1076 3653 1196
rect 3666 1193 3669 1206
rect 3694 1176 3697 1223
rect 3730 1216 3733 1333
rect 3746 1236 3749 1336
rect 3694 1173 3701 1176
rect 3650 1073 3661 1076
rect 3674 1073 3677 1136
rect 3574 913 3581 916
rect 3578 843 3581 913
rect 3594 906 3597 966
rect 3626 963 3629 1016
rect 3590 903 3597 906
rect 3590 836 3593 903
rect 3590 833 3597 836
rect 3570 743 3573 816
rect 3594 813 3597 833
rect 3602 823 3605 926
rect 3610 916 3613 936
rect 3610 913 3621 916
rect 3618 856 3621 913
rect 3610 853 3621 856
rect 3578 753 3581 806
rect 3578 743 3597 746
rect 3562 683 3565 726
rect 3554 616 3557 636
rect 3554 613 3565 616
rect 3554 593 3557 606
rect 3538 583 3549 586
rect 3506 446 3509 536
rect 3514 523 3517 536
rect 3538 533 3541 583
rect 3546 503 3549 576
rect 3562 546 3565 613
rect 3570 603 3573 736
rect 3578 723 3581 743
rect 3586 723 3589 736
rect 3594 733 3597 743
rect 3602 716 3605 816
rect 3610 793 3613 853
rect 3618 813 3621 836
rect 3634 823 3637 1016
rect 3642 923 3645 1066
rect 3658 1026 3661 1073
rect 3650 1023 3661 1026
rect 3594 713 3605 716
rect 3594 683 3597 713
rect 3578 613 3581 626
rect 3558 543 3565 546
rect 3558 496 3561 543
rect 3570 533 3573 546
rect 3578 533 3581 606
rect 3594 556 3597 616
rect 3602 603 3605 706
rect 3594 553 3605 556
rect 3554 493 3561 496
rect 3570 493 3573 526
rect 3498 443 3509 446
rect 3482 413 3485 426
rect 3498 396 3501 443
rect 3498 393 3509 396
rect 3506 336 3509 393
rect 3530 366 3533 486
rect 3554 396 3557 493
rect 3562 403 3565 416
rect 3570 413 3573 426
rect 3578 413 3581 436
rect 3586 413 3589 526
rect 3594 433 3597 546
rect 3602 533 3605 553
rect 3610 476 3613 726
rect 3618 706 3621 726
rect 3618 703 3625 706
rect 3622 636 3625 703
rect 3634 673 3637 816
rect 3650 766 3653 1023
rect 3666 906 3669 936
rect 3658 903 3669 906
rect 3658 813 3661 903
rect 3666 803 3669 826
rect 3674 786 3677 1056
rect 3682 976 3685 1096
rect 3690 1063 3693 1156
rect 3682 973 3689 976
rect 3686 826 3689 973
rect 3686 823 3693 826
rect 3670 783 3677 786
rect 3650 763 3661 766
rect 3618 633 3625 636
rect 3618 613 3621 633
rect 3626 603 3637 606
rect 3626 513 3629 526
rect 3634 523 3637 603
rect 3642 516 3645 756
rect 3658 676 3661 763
rect 3650 673 3661 676
rect 3670 676 3673 783
rect 3682 753 3685 806
rect 3690 786 3693 823
rect 3698 803 3701 1173
rect 3706 896 3709 1216
rect 3718 1213 3733 1216
rect 3738 1233 3749 1236
rect 3738 1213 3741 1233
rect 3746 1213 3757 1216
rect 3718 1036 3721 1213
rect 3770 1196 3773 1383
rect 3762 1193 3773 1196
rect 3730 1143 3749 1146
rect 3730 1123 3733 1143
rect 3738 1093 3741 1136
rect 3746 1133 3749 1143
rect 3746 1083 3749 1126
rect 3762 1116 3765 1193
rect 3762 1113 3773 1116
rect 3714 1033 3721 1036
rect 3714 973 3717 1033
rect 3714 913 3717 926
rect 3722 923 3725 1016
rect 3738 906 3741 976
rect 3730 903 3741 906
rect 3706 893 3717 896
rect 3690 783 3697 786
rect 3670 673 3677 676
rect 3650 543 3653 673
rect 3638 513 3645 516
rect 3610 473 3621 476
rect 3610 413 3613 426
rect 3554 393 3573 396
rect 3530 363 3549 366
rect 3506 333 3517 336
rect 3458 313 3461 326
rect 3466 323 3477 326
rect 3498 313 3501 326
rect 3514 266 3517 333
rect 3498 263 3517 266
rect 3418 183 3421 206
rect 3434 196 3437 216
rect 3442 203 3445 216
rect 3450 213 3453 246
rect 3450 196 3453 206
rect 3434 193 3453 196
rect 3458 133 3461 156
rect 3474 123 3477 186
rect 3490 143 3493 216
rect 3498 213 3501 263
rect 3546 153 3549 363
rect 3562 243 3565 336
rect 3570 313 3573 393
rect 3554 213 3557 236
rect 3578 193 3581 336
rect 3586 246 3589 326
rect 3618 303 3621 473
rect 3626 323 3629 496
rect 3638 456 3641 513
rect 3650 493 3653 536
rect 3666 533 3669 656
rect 3666 513 3669 526
rect 3674 523 3677 673
rect 3682 613 3685 726
rect 3694 656 3697 783
rect 3714 766 3717 893
rect 3690 653 3697 656
rect 3706 763 3717 766
rect 3730 766 3733 903
rect 3746 773 3749 1076
rect 3762 1013 3765 1096
rect 3770 996 3773 1113
rect 3766 993 3773 996
rect 3754 923 3757 936
rect 3766 916 3769 993
rect 3778 923 3781 1226
rect 3786 1186 3789 1446
rect 3794 1433 3797 1536
rect 3802 1523 3805 1536
rect 3810 1496 3813 1516
rect 3806 1493 3813 1496
rect 3806 1416 3809 1493
rect 3818 1443 3821 1543
rect 3826 1533 3829 1616
rect 3834 1613 3837 1943
rect 3842 1853 3845 2126
rect 3850 1933 3853 2006
rect 3858 2003 3861 2173
rect 3874 2046 3877 2253
rect 3886 2236 3889 2303
rect 3886 2233 3893 2236
rect 3890 2196 3893 2233
rect 3886 2193 3893 2196
rect 3886 2106 3889 2193
rect 3898 2116 3901 2396
rect 3906 2323 3909 2403
rect 3914 2346 3917 2483
rect 3938 2403 3941 2486
rect 3922 2366 3925 2386
rect 3922 2363 3933 2366
rect 3914 2343 3921 2346
rect 3906 2203 3909 2306
rect 3918 2276 3921 2343
rect 3914 2273 3921 2276
rect 3914 2133 3917 2273
rect 3930 2256 3933 2363
rect 3954 2333 3957 2536
rect 3962 2533 3965 2543
rect 3962 2513 3965 2526
rect 3978 2466 3981 2553
rect 3970 2463 3981 2466
rect 3994 2466 3997 2773
rect 4010 2756 4013 3073
rect 4034 2986 4037 3093
rect 4058 3056 4061 3153
rect 4066 3126 4069 3146
rect 4066 3123 4077 3126
rect 4050 3053 4061 3056
rect 4050 3006 4053 3053
rect 4074 3046 4077 3123
rect 4106 3053 4109 3146
rect 4066 3043 4077 3046
rect 4050 3003 4061 3006
rect 4034 2983 4045 2986
rect 4058 2983 4061 3003
rect 4042 2963 4045 2983
rect 4050 2933 4053 2946
rect 4018 2813 4021 2836
rect 4026 2813 4029 2926
rect 4006 2753 4013 2756
rect 4006 2706 4009 2753
rect 4006 2703 4013 2706
rect 4010 2636 4013 2703
rect 4010 2633 4017 2636
rect 4002 2593 4005 2616
rect 4014 2576 4017 2633
rect 4010 2573 4017 2576
rect 4010 2536 4013 2573
rect 4006 2533 4013 2536
rect 4006 2486 4009 2533
rect 4006 2483 4013 2486
rect 3994 2463 4001 2466
rect 3962 2343 3965 2356
rect 3922 2253 3933 2256
rect 3922 2176 3925 2253
rect 3938 2196 3941 2216
rect 3946 2203 3949 2236
rect 3954 2213 3957 2316
rect 3954 2196 3957 2206
rect 3938 2193 3957 2196
rect 3962 2176 3965 2326
rect 3970 2296 3973 2463
rect 3998 2356 4001 2463
rect 3986 2333 3989 2356
rect 3998 2353 4005 2356
rect 4002 2333 4005 2353
rect 3978 2313 3981 2326
rect 3994 2306 3997 2326
rect 3990 2303 3997 2306
rect 3970 2293 3981 2296
rect 3978 2216 3981 2293
rect 3922 2173 3933 2176
rect 3930 2126 3933 2173
rect 3922 2123 3933 2126
rect 3946 2173 3965 2176
rect 3970 2213 3981 2216
rect 3898 2113 3909 2116
rect 3886 2103 3893 2106
rect 3866 2043 3877 2046
rect 3842 1613 3845 1706
rect 3850 1633 3853 1736
rect 3858 1733 3861 1796
rect 3866 1643 3869 2043
rect 3874 1953 3877 2006
rect 3882 1983 3885 2026
rect 3890 2003 3893 2103
rect 3906 2036 3909 2113
rect 3898 2033 3909 2036
rect 3898 1986 3901 2033
rect 3894 1983 3901 1986
rect 3874 1793 3877 1816
rect 3882 1743 3885 1926
rect 3894 1826 3897 1983
rect 3906 1943 3909 2016
rect 3906 1923 3909 1936
rect 3922 1906 3925 2123
rect 3946 1996 3949 2173
rect 3970 2133 3973 2213
rect 3990 2196 3993 2303
rect 3986 2193 3993 2196
rect 3970 2003 3973 2046
rect 3978 2013 3981 2136
rect 3986 2023 3989 2193
rect 3946 1993 3965 1996
rect 3906 1903 3925 1906
rect 3894 1823 3901 1826
rect 3874 1713 3877 1726
rect 3882 1693 3885 1736
rect 3890 1733 3893 1806
rect 3834 1563 3837 1606
rect 3842 1456 3845 1606
rect 3850 1573 3853 1626
rect 3866 1593 3869 1636
rect 3838 1453 3845 1456
rect 3802 1413 3809 1416
rect 3818 1413 3821 1426
rect 3826 1413 3829 1436
rect 3802 1346 3805 1413
rect 3802 1343 3813 1346
rect 3794 1313 3797 1326
rect 3802 1296 3805 1326
rect 3798 1293 3805 1296
rect 3798 1226 3801 1293
rect 3794 1223 3801 1226
rect 3794 1203 3797 1223
rect 3786 1183 3793 1186
rect 3790 916 3793 1183
rect 3766 913 3773 916
rect 3762 813 3765 826
rect 3730 763 3741 766
rect 3706 653 3709 763
rect 3714 733 3717 746
rect 3714 706 3717 726
rect 3722 723 3725 736
rect 3714 703 3721 706
rect 3634 453 3641 456
rect 3634 333 3637 453
rect 3658 403 3661 416
rect 3674 366 3677 406
rect 3682 393 3685 506
rect 3690 403 3693 653
rect 3718 646 3721 703
rect 3714 643 3721 646
rect 3674 363 3685 366
rect 3642 333 3653 336
rect 3674 333 3677 356
rect 3634 283 3637 326
rect 3650 246 3653 326
rect 3666 313 3669 326
rect 3674 303 3677 326
rect 3682 276 3685 363
rect 3706 356 3709 406
rect 3714 373 3717 643
rect 3730 583 3733 696
rect 3738 613 3741 763
rect 3762 753 3765 806
rect 3762 723 3765 736
rect 3762 586 3765 606
rect 3754 583 3765 586
rect 3754 466 3757 583
rect 3770 566 3773 913
rect 3786 913 3793 916
rect 3778 743 3781 816
rect 3786 686 3789 913
rect 3794 803 3797 816
rect 3802 706 3805 1216
rect 3810 1203 3813 1343
rect 3818 1186 3821 1406
rect 3838 1376 3841 1453
rect 3890 1446 3893 1726
rect 3898 1533 3901 1823
rect 3906 1733 3909 1903
rect 3914 1793 3917 1806
rect 3906 1613 3909 1726
rect 3914 1546 3917 1746
rect 3922 1673 3925 1836
rect 3930 1813 3933 1936
rect 3938 1923 3941 1936
rect 3938 1783 3941 1806
rect 3946 1746 3949 1816
rect 3930 1743 3949 1746
rect 3930 1696 3933 1743
rect 3938 1713 3941 1736
rect 3930 1693 3937 1696
rect 3934 1576 3937 1693
rect 3910 1543 3917 1546
rect 3930 1573 3937 1576
rect 3910 1476 3913 1543
rect 3930 1536 3933 1573
rect 3922 1533 3933 1536
rect 3910 1473 3917 1476
rect 3914 1453 3917 1473
rect 3882 1443 3893 1446
rect 3858 1413 3861 1426
rect 3838 1373 3845 1376
rect 3834 1313 3837 1326
rect 3814 1183 3821 1186
rect 3814 1086 3817 1183
rect 3826 1093 3829 1206
rect 3834 1193 3837 1206
rect 3814 1083 3821 1086
rect 3818 1056 3821 1083
rect 3814 1053 3821 1056
rect 3814 976 3817 1053
rect 3834 1013 3837 1126
rect 3842 993 3845 1373
rect 3882 1363 3885 1443
rect 3906 1393 3909 1406
rect 3914 1346 3917 1366
rect 3882 1333 3885 1346
rect 3906 1343 3917 1346
rect 3814 973 3821 976
rect 3818 953 3821 973
rect 3810 723 3813 946
rect 3834 933 3837 956
rect 3818 896 3821 916
rect 3842 913 3845 936
rect 3818 893 3829 896
rect 3826 846 3829 893
rect 3842 886 3845 906
rect 3818 843 3829 846
rect 3838 883 3845 886
rect 3818 723 3821 843
rect 3826 813 3829 826
rect 3826 783 3829 806
rect 3838 786 3841 883
rect 3850 823 3853 1246
rect 3858 923 3861 1216
rect 3866 1133 3869 1216
rect 3874 1213 3877 1246
rect 3874 1123 3877 1206
rect 3882 1133 3885 1316
rect 3906 1246 3909 1343
rect 3922 1256 3925 1533
rect 3930 1506 3933 1526
rect 3930 1503 3937 1506
rect 3934 1426 3937 1503
rect 3930 1423 3937 1426
rect 3930 1313 3933 1423
rect 3938 1383 3941 1406
rect 3938 1333 3941 1346
rect 3922 1253 3929 1256
rect 3906 1243 3917 1246
rect 3890 1196 3893 1216
rect 3898 1203 3901 1216
rect 3906 1213 3909 1226
rect 3906 1196 3909 1206
rect 3890 1193 3909 1196
rect 3890 1123 3893 1186
rect 3882 1003 3885 1016
rect 3898 1013 3901 1136
rect 3906 1113 3909 1126
rect 3914 1096 3917 1243
rect 3910 1093 3917 1096
rect 3910 1006 3913 1093
rect 3926 1056 3929 1253
rect 3946 1243 3949 1736
rect 3954 1693 3957 1746
rect 3962 1733 3965 1993
rect 3994 1933 3997 2136
rect 4002 2096 4005 2326
rect 4010 2196 4013 2483
rect 4018 2413 4021 2526
rect 4026 2483 4029 2806
rect 4034 2803 4037 2826
rect 4058 2793 4061 2806
rect 4066 2803 4069 3043
rect 4074 2943 4077 3006
rect 4082 2916 4085 2986
rect 4090 2953 4093 3006
rect 4090 2923 4093 2936
rect 4114 2923 4117 3016
rect 4082 2913 4093 2916
rect 4090 2826 4093 2913
rect 4130 2906 4133 3126
rect 4138 3123 4141 3203
rect 4170 3143 4173 3336
rect 4210 3323 4213 3336
rect 4218 3306 4221 3356
rect 4210 3303 4221 3306
rect 4186 3193 4189 3216
rect 4210 3146 4213 3303
rect 4210 3143 4221 3146
rect 4170 3026 4173 3136
rect 4202 3063 4205 3126
rect 4162 3023 4173 3026
rect 4122 2903 4133 2906
rect 4138 2906 4141 2926
rect 4162 2906 4165 3023
rect 4178 2916 4181 3016
rect 4186 3013 4189 3026
rect 4218 3016 4221 3143
rect 4226 3123 4229 3206
rect 4234 3143 4237 3443
rect 4258 3436 4261 3503
rect 4258 3433 4269 3436
rect 4242 3396 4245 3406
rect 4250 3403 4253 3416
rect 4242 3393 4253 3396
rect 4258 3393 4261 3406
rect 4242 3193 4245 3386
rect 4250 3376 4253 3393
rect 4250 3373 4257 3376
rect 4254 3186 4257 3373
rect 4250 3183 4257 3186
rect 4250 3136 4253 3183
rect 4234 3106 4237 3136
rect 4250 3133 4257 3136
rect 4230 3103 4237 3106
rect 4230 3036 4233 3103
rect 4230 3033 4237 3036
rect 4218 3013 4225 3016
rect 4202 2933 4205 2946
rect 4210 2916 4213 3006
rect 4178 2913 4189 2916
rect 4138 2903 4149 2906
rect 4162 2903 4173 2906
rect 4122 2846 4125 2903
rect 4146 2856 4149 2903
rect 4138 2853 4149 2856
rect 4122 2843 4133 2846
rect 4090 2823 4101 2826
rect 4130 2823 4133 2843
rect 4074 2766 4077 2816
rect 4070 2763 4077 2766
rect 4034 2513 4037 2526
rect 4042 2413 4045 2616
rect 4058 2613 4061 2726
rect 4018 2323 4021 2406
rect 4042 2393 4045 2406
rect 4058 2376 4061 2536
rect 4070 2486 4073 2763
rect 4098 2746 4101 2823
rect 4130 2803 4133 2816
rect 4138 2813 4141 2853
rect 4154 2813 4157 2836
rect 4090 2743 4101 2746
rect 4090 2686 4093 2743
rect 4082 2683 4093 2686
rect 4082 2493 4085 2683
rect 4098 2603 4101 2626
rect 4106 2603 4109 2726
rect 4090 2576 4093 2596
rect 4114 2593 4117 2616
rect 4122 2603 4125 2616
rect 4130 2613 4133 2646
rect 4138 2606 4141 2806
rect 4130 2603 4141 2606
rect 4146 2603 4149 2806
rect 4154 2623 4157 2726
rect 4162 2723 4165 2796
rect 4170 2736 4173 2903
rect 4186 2836 4189 2913
rect 4178 2833 4189 2836
rect 4202 2913 4213 2916
rect 4202 2836 4205 2913
rect 4222 2906 4225 3013
rect 4234 2933 4237 3033
rect 4242 3013 4245 3126
rect 4254 3036 4257 3133
rect 4250 3033 4257 3036
rect 4250 2946 4253 3033
rect 4258 2993 4261 3016
rect 4266 2986 4269 3433
rect 4274 3276 4277 3536
rect 4282 3296 4285 3703
rect 4290 3313 4293 3626
rect 4298 3543 4301 3833
rect 4306 3793 4309 3996
rect 4322 3966 4325 4016
rect 4330 3993 4333 4236
rect 4338 4003 4341 4216
rect 4346 4213 4349 4256
rect 4362 4233 4365 4336
rect 4370 4303 4373 4326
rect 4394 4226 4397 4356
rect 4402 4333 4405 4426
rect 4410 4396 4413 4406
rect 4418 4403 4421 4416
rect 4426 4396 4429 4416
rect 4410 4393 4429 4396
rect 4434 4346 4437 4433
rect 4426 4343 4437 4346
rect 4394 4223 4401 4226
rect 4346 4196 4349 4206
rect 4354 4203 4357 4216
rect 4362 4196 4365 4216
rect 4346 4193 4365 4196
rect 4370 4193 4373 4206
rect 4346 3973 4349 4146
rect 4354 4113 4357 4126
rect 4322 3963 4341 3966
rect 4298 3513 4301 3526
rect 4298 3413 4301 3426
rect 4298 3333 4301 3406
rect 4306 3403 4309 3736
rect 4314 3513 4317 3946
rect 4322 3813 4325 3963
rect 4338 3933 4341 3963
rect 4354 3943 4357 4096
rect 4362 3933 4365 4006
rect 4330 3813 4333 3826
rect 4322 3423 4325 3806
rect 4338 3793 4341 3926
rect 4330 3523 4333 3726
rect 4346 3716 4349 3736
rect 4342 3713 4349 3716
rect 4342 3636 4345 3713
rect 4342 3633 4349 3636
rect 4346 3613 4349 3633
rect 4338 3526 4341 3606
rect 4354 3543 4357 3736
rect 4362 3733 4365 3816
rect 4362 3596 4365 3696
rect 4370 3633 4373 4056
rect 4378 3983 4381 4216
rect 4386 4133 4389 4216
rect 4398 4176 4401 4223
rect 4394 4173 4401 4176
rect 4386 4013 4389 4116
rect 4394 4113 4397 4173
rect 4410 4156 4413 4336
rect 4426 4326 4429 4343
rect 4422 4323 4429 4326
rect 4422 4246 4425 4323
rect 4422 4243 4429 4246
rect 4418 4213 4421 4226
rect 4402 4153 4413 4156
rect 4402 4096 4405 4153
rect 4410 4123 4413 4146
rect 4398 4093 4405 4096
rect 4398 4026 4401 4093
rect 4398 4023 4405 4026
rect 4394 3993 4397 4006
rect 4402 3966 4405 4023
rect 4410 3986 4413 4116
rect 4418 4103 4421 4156
rect 4426 4133 4429 4243
rect 4434 4213 4437 4336
rect 4442 4333 4445 4406
rect 4450 4353 4453 4483
rect 4458 4403 4461 4446
rect 4466 4396 4469 4416
rect 4474 4403 4477 4523
rect 4490 4513 4493 4616
rect 4562 4613 4565 4626
rect 4642 4623 4645 4740
rect 4586 4573 4589 4606
rect 4482 4413 4485 4436
rect 4482 4396 4485 4406
rect 4466 4393 4485 4396
rect 4458 4333 4461 4346
rect 4442 4313 4445 4326
rect 4482 4313 4485 4326
rect 4538 4306 4541 4326
rect 4546 4316 4549 4446
rect 4554 4413 4557 4526
rect 4562 4393 4565 4456
rect 4586 4446 4589 4536
rect 4602 4453 4605 4526
rect 4610 4456 4613 4616
rect 4754 4613 4757 4626
rect 4778 4576 4781 4606
rect 4682 4533 4685 4576
rect 4778 4573 4789 4576
rect 4610 4453 4625 4456
rect 4586 4443 4613 4446
rect 4570 4343 4573 4406
rect 4578 4396 4581 4416
rect 4586 4403 4589 4426
rect 4594 4416 4597 4436
rect 4594 4413 4605 4416
rect 4594 4396 4597 4406
rect 4578 4393 4597 4396
rect 4602 4336 4605 4413
rect 4554 4333 4573 4336
rect 4546 4313 4553 4316
rect 4530 4303 4541 4306
rect 4442 4133 4445 4146
rect 4434 4056 4437 4126
rect 4450 4123 4453 4256
rect 4530 4236 4533 4303
rect 4550 4256 4553 4313
rect 4550 4253 4565 4256
rect 4530 4233 4541 4236
rect 4490 4203 4493 4216
rect 4418 4053 4437 4056
rect 4418 4003 4421 4053
rect 4458 4043 4461 4126
rect 4474 4106 4477 4126
rect 4498 4123 4501 4216
rect 4514 4213 4533 4216
rect 4538 4213 4541 4233
rect 4546 4213 4549 4226
rect 4506 4186 4509 4206
rect 4506 4183 4513 4186
rect 4510 4116 4513 4183
rect 4506 4113 4513 4116
rect 4474 4103 4485 4106
rect 4482 4036 4485 4103
rect 4426 4003 4429 4016
rect 4442 4013 4445 4036
rect 4474 4033 4485 4036
rect 4450 3993 4453 4026
rect 4410 3983 4429 3986
rect 4402 3963 4413 3966
rect 4386 3913 4389 3926
rect 4410 3886 4413 3963
rect 4402 3883 4413 3886
rect 4378 3693 4381 3846
rect 4402 3843 4405 3883
rect 4426 3866 4429 3983
rect 4458 3946 4461 4006
rect 4474 3993 4477 4033
rect 4506 4023 4509 4113
rect 4522 4096 4525 4136
rect 4518 4093 4525 4096
rect 4518 4026 4521 4093
rect 4530 4053 4533 4213
rect 4546 4193 4549 4206
rect 4562 4183 4565 4253
rect 4570 4213 4573 4333
rect 4586 4333 4605 4336
rect 4578 4313 4581 4326
rect 4578 4193 4581 4206
rect 4518 4023 4525 4026
rect 4410 3863 4429 3866
rect 4450 3943 4461 3946
rect 4450 3866 4453 3943
rect 4450 3863 4461 3866
rect 4386 3733 4397 3736
rect 4386 3723 4397 3726
rect 4370 3613 4373 3626
rect 4402 3606 4405 3836
rect 4410 3793 4413 3863
rect 4410 3723 4413 3736
rect 4418 3723 4421 3816
rect 4426 3646 4429 3796
rect 4442 3743 4445 3806
rect 4458 3776 4461 3863
rect 4454 3773 4461 3776
rect 4454 3726 4457 3773
rect 4418 3643 4429 3646
rect 4450 3723 4457 3726
rect 4450 3646 4453 3723
rect 4450 3643 4461 3646
rect 4402 3603 4409 3606
rect 4362 3593 4369 3596
rect 4366 3536 4369 3593
rect 4362 3533 4369 3536
rect 4338 3523 4349 3526
rect 4330 3416 4333 3436
rect 4322 3413 4333 3416
rect 4306 3323 4309 3396
rect 4314 3333 4317 3366
rect 4322 3333 4325 3413
rect 4322 3306 4325 3326
rect 4314 3303 4325 3306
rect 4282 3293 4301 3296
rect 4274 3273 4285 3276
rect 4282 3196 4285 3273
rect 4242 2943 4253 2946
rect 4258 2983 4269 2986
rect 4274 3193 4285 3196
rect 4274 2983 4277 3193
rect 4298 3176 4301 3293
rect 4282 3173 4301 3176
rect 4314 3176 4317 3303
rect 4330 3286 4333 3406
rect 4338 3396 4341 3416
rect 4346 3403 4349 3523
rect 4362 3433 4365 3533
rect 4378 3503 4381 3536
rect 4394 3533 4397 3596
rect 4406 3556 4409 3603
rect 4418 3573 4421 3643
rect 4458 3626 4461 3643
rect 4434 3613 4437 3626
rect 4450 3623 4461 3626
rect 4466 3623 4469 3926
rect 4474 3803 4477 3936
rect 4482 3933 4485 4006
rect 4498 3993 4501 4006
rect 4522 4003 4525 4023
rect 4554 3966 4557 4156
rect 4586 4123 4589 4333
rect 4594 4306 4597 4326
rect 4610 4323 4613 4443
rect 4622 4406 4625 4453
rect 4634 4413 4637 4426
rect 4642 4413 4645 4436
rect 4622 4403 4629 4406
rect 4626 4336 4629 4403
rect 4626 4333 4641 4336
rect 4626 4313 4629 4326
rect 4594 4303 4605 4306
rect 4602 4226 4605 4303
rect 4638 4266 4641 4333
rect 4650 4276 4653 4496
rect 4658 4413 4661 4526
rect 4698 4493 4701 4526
rect 4754 4513 4757 4526
rect 4674 4413 4677 4426
rect 4674 4323 4677 4376
rect 4722 4373 4725 4406
rect 4786 4386 4789 4573
rect 4778 4383 4789 4386
rect 4650 4273 4661 4276
rect 4638 4263 4645 4266
rect 4594 4223 4605 4226
rect 4594 4203 4597 4223
rect 4642 4216 4645 4263
rect 4602 4146 4605 4206
rect 4594 4143 4605 4146
rect 4594 4133 4597 4143
rect 4610 4136 4613 4186
rect 4618 4146 4621 4216
rect 4642 4213 4649 4216
rect 4626 4183 4629 4206
rect 4634 4153 4637 4206
rect 4646 4146 4649 4213
rect 4618 4143 4629 4146
rect 4602 4123 4605 4136
rect 4610 4133 4621 4136
rect 4626 4133 4629 4143
rect 4642 4143 4649 4146
rect 4562 4013 4565 4026
rect 4586 4003 4589 4016
rect 4602 4013 4605 4026
rect 4610 4003 4613 4126
rect 4550 3963 4557 3966
rect 4626 3966 4629 4126
rect 4626 3963 4637 3966
rect 4482 3823 4485 3926
rect 4490 3923 4493 3936
rect 4490 3816 4493 3886
rect 4482 3813 4493 3816
rect 4482 3796 4485 3813
rect 4474 3793 4485 3796
rect 4474 3723 4477 3793
rect 4490 3756 4493 3806
rect 4498 3786 4501 3906
rect 4506 3863 4509 3926
rect 4530 3923 4533 3936
rect 4506 3793 4509 3806
rect 4514 3803 4517 3826
rect 4522 3813 4525 3916
rect 4538 3826 4541 3936
rect 4550 3886 4553 3963
rect 4618 3933 4621 3946
rect 4550 3883 4557 3886
rect 4534 3823 4541 3826
rect 4554 3826 4557 3883
rect 4586 3826 4589 3926
rect 4634 3923 4637 3963
rect 4554 3823 4561 3826
rect 4498 3783 4517 3786
rect 4482 3753 4493 3756
rect 4450 3606 4453 3623
rect 4458 3613 4469 3616
rect 4426 3603 4445 3606
rect 4450 3603 4461 3606
rect 4402 3553 4409 3556
rect 4386 3523 4397 3526
rect 4338 3393 4349 3396
rect 4354 3393 4357 3406
rect 4326 3283 4333 3286
rect 4326 3196 4329 3283
rect 4326 3193 4333 3196
rect 4314 3173 4325 3176
rect 4218 2903 4225 2906
rect 4202 2833 4213 2836
rect 4178 2803 4181 2833
rect 4178 2743 4181 2786
rect 4202 2763 4205 2816
rect 4210 2793 4213 2833
rect 4170 2733 4181 2736
rect 4194 2733 4197 2746
rect 4178 2716 4181 2733
rect 4162 2713 4181 2716
rect 4090 2573 4097 2576
rect 4094 2486 4097 2573
rect 4106 2503 4109 2526
rect 4070 2483 4077 2486
rect 4074 2456 4077 2483
rect 4070 2453 4077 2456
rect 4090 2483 4097 2486
rect 4090 2456 4093 2483
rect 4090 2453 4097 2456
rect 4070 2386 4073 2453
rect 4070 2383 4077 2386
rect 4054 2373 4061 2376
rect 4026 2293 4029 2326
rect 4018 2213 4021 2226
rect 4010 2193 4017 2196
rect 4014 2116 4017 2193
rect 4026 2133 4029 2236
rect 4034 2133 4037 2336
rect 4054 2316 4057 2373
rect 4066 2323 4069 2366
rect 4054 2313 4061 2316
rect 4014 2113 4021 2116
rect 4002 2093 4009 2096
rect 4006 1986 4009 2093
rect 4002 1983 4009 1986
rect 3978 1836 3981 1856
rect 3974 1833 3981 1836
rect 3974 1786 3977 1833
rect 3986 1793 3989 1926
rect 4002 1853 4005 1983
rect 4018 1966 4021 2113
rect 4042 2106 4045 2296
rect 4058 2246 4061 2313
rect 4058 2243 4069 2246
rect 4058 2213 4061 2226
rect 4014 1963 4021 1966
rect 4034 2103 4045 2106
rect 4014 1856 4017 1963
rect 4026 1883 4029 1936
rect 4010 1853 4017 1856
rect 4010 1833 4013 1853
rect 3974 1783 3981 1786
rect 3978 1736 3981 1783
rect 3962 1713 3965 1726
rect 3954 1596 3957 1656
rect 3970 1613 3973 1736
rect 3978 1733 3989 1736
rect 3978 1703 3981 1726
rect 3954 1593 3965 1596
rect 3962 1436 3965 1593
rect 3978 1483 3981 1636
rect 3986 1606 3989 1733
rect 3994 1723 3997 1826
rect 4002 1813 4021 1816
rect 3994 1613 3997 1636
rect 4002 1616 4005 1813
rect 4010 1756 4013 1806
rect 4018 1773 4021 1806
rect 4010 1753 4021 1756
rect 4018 1676 4021 1753
rect 4010 1673 4021 1676
rect 4010 1653 4013 1673
rect 4034 1653 4037 2103
rect 4050 2086 4053 2136
rect 4066 2133 4069 2243
rect 4046 2083 4053 2086
rect 4046 1986 4049 2083
rect 4058 1993 4061 2126
rect 4046 1983 4053 1986
rect 4050 1936 4053 1983
rect 4042 1923 4045 1936
rect 4050 1933 4061 1936
rect 4066 1933 4069 2126
rect 4074 2083 4077 2383
rect 4082 2166 4085 2376
rect 4094 2366 4097 2453
rect 4106 2396 4109 2496
rect 4122 2443 4125 2526
rect 4130 2503 4133 2603
rect 4138 2533 4141 2546
rect 4138 2493 4141 2526
rect 4114 2413 4117 2426
rect 4154 2413 4157 2426
rect 4106 2393 4125 2396
rect 4138 2393 4141 2406
rect 4090 2363 4097 2366
rect 4090 2313 4093 2363
rect 4098 2343 4117 2346
rect 4098 2323 4101 2343
rect 4106 2303 4109 2336
rect 4114 2333 4117 2343
rect 4122 2323 4125 2393
rect 4130 2306 4133 2336
rect 4122 2303 4133 2306
rect 4122 2246 4125 2303
rect 4122 2243 4133 2246
rect 4106 2193 4109 2206
rect 4122 2203 4125 2216
rect 4122 2176 4125 2196
rect 4118 2173 4125 2176
rect 4082 2163 4093 2166
rect 4074 1976 4077 2076
rect 4090 2056 4093 2163
rect 4118 2096 4121 2173
rect 4118 2093 4125 2096
rect 4082 2053 4093 2056
rect 4082 1996 4085 2053
rect 4090 2013 4093 2036
rect 4106 2013 4109 2026
rect 4122 2013 4125 2093
rect 4130 1996 4133 2243
rect 4138 2193 4141 2326
rect 4162 2153 4165 2713
rect 4170 2613 4173 2686
rect 4186 2613 4189 2636
rect 4170 2403 4173 2446
rect 4178 2426 4181 2606
rect 4194 2543 4197 2726
rect 4218 2686 4221 2903
rect 4214 2683 4221 2686
rect 4214 2606 4217 2683
rect 4226 2613 4229 2796
rect 4234 2676 4237 2926
rect 4242 2903 4245 2943
rect 4242 2753 4245 2816
rect 4250 2766 4253 2936
rect 4258 2923 4261 2983
rect 4274 2913 4277 2926
rect 4282 2896 4285 3173
rect 4290 3113 4293 3136
rect 4290 2993 4293 3016
rect 4306 3013 4309 3136
rect 4314 3123 4317 3156
rect 4322 3106 4325 3173
rect 4318 3103 4325 3106
rect 4318 3036 4321 3103
rect 4318 3033 4325 3036
rect 4322 3013 4325 3033
rect 4330 3006 4333 3193
rect 4274 2893 4285 2896
rect 4258 2803 4261 2846
rect 4274 2826 4277 2893
rect 4274 2823 4285 2826
rect 4266 2776 4269 2806
rect 4266 2773 4277 2776
rect 4250 2763 4261 2766
rect 4258 2746 4261 2763
rect 4258 2743 4265 2746
rect 4242 2713 4245 2726
rect 4262 2686 4265 2743
rect 4258 2683 4265 2686
rect 4234 2673 4245 2676
rect 4202 2533 4205 2606
rect 4214 2603 4221 2606
rect 4178 2423 4185 2426
rect 4182 2366 4185 2423
rect 4194 2373 4197 2526
rect 4202 2496 4205 2526
rect 4218 2513 4221 2603
rect 4234 2593 4237 2616
rect 4226 2533 4229 2546
rect 4234 2496 4237 2536
rect 4242 2523 4245 2673
rect 4258 2666 4261 2683
rect 4254 2663 4261 2666
rect 4254 2596 4257 2663
rect 4274 2656 4277 2773
rect 4266 2653 4277 2656
rect 4266 2603 4269 2653
rect 4282 2613 4285 2823
rect 4290 2803 4293 2936
rect 4298 2906 4301 3006
rect 4306 2923 4309 3006
rect 4314 3003 4333 3006
rect 4314 2993 4317 3003
rect 4298 2903 4305 2906
rect 4302 2826 4305 2903
rect 4302 2823 4309 2826
rect 4290 2733 4293 2756
rect 4290 2713 4293 2726
rect 4274 2603 4285 2606
rect 4254 2593 4261 2596
rect 4250 2543 4253 2556
rect 4258 2526 4261 2593
rect 4274 2553 4277 2603
rect 4266 2533 4269 2546
rect 4254 2523 4261 2526
rect 4202 2493 4213 2496
rect 4210 2436 4213 2493
rect 4202 2433 4213 2436
rect 4226 2493 4237 2496
rect 4202 2413 4205 2433
rect 4182 2363 4189 2366
rect 4186 2276 4189 2363
rect 4194 2296 4197 2316
rect 4218 2313 4221 2326
rect 4226 2323 4229 2493
rect 4242 2393 4245 2516
rect 4254 2356 4257 2523
rect 4266 2366 4269 2526
rect 4274 2503 4277 2526
rect 4266 2363 4273 2366
rect 4234 2333 4237 2356
rect 4254 2353 4261 2356
rect 4194 2293 4213 2296
rect 4138 2013 4141 2126
rect 4082 1993 4093 1996
rect 4074 1973 4081 1976
rect 4058 1876 4061 1933
rect 4078 1926 4081 1973
rect 4050 1873 4061 1876
rect 4074 1923 4081 1926
rect 4050 1816 4053 1873
rect 4050 1813 4061 1816
rect 4066 1813 4069 1866
rect 4058 1793 4061 1813
rect 4042 1733 4045 1756
rect 4074 1726 4077 1923
rect 4090 1846 4093 1993
rect 4122 1993 4133 1996
rect 4122 1916 4125 1993
rect 4146 1983 4149 2006
rect 4154 1966 4157 2086
rect 4162 2043 4165 2136
rect 4178 2096 4181 2276
rect 4186 2273 4197 2276
rect 4194 2196 4197 2273
rect 4174 2093 4181 2096
rect 4186 2193 4197 2196
rect 4174 2036 4177 2093
rect 4186 2046 4189 2193
rect 4210 2176 4213 2293
rect 4242 2283 4245 2326
rect 4250 2323 4253 2336
rect 4250 2213 4253 2316
rect 4258 2196 4261 2353
rect 4270 2256 4273 2363
rect 4282 2323 4285 2596
rect 4290 2483 4293 2646
rect 4298 2416 4301 2816
rect 4306 2636 4309 2823
rect 4314 2683 4317 2986
rect 4322 2976 4325 2996
rect 4338 2993 4341 3386
rect 4346 3356 4349 3393
rect 4346 3353 4357 3356
rect 4346 3276 4349 3346
rect 4354 3296 4357 3353
rect 4362 3333 4365 3416
rect 4386 3406 4389 3426
rect 4378 3403 4389 3406
rect 4378 3356 4381 3403
rect 4378 3353 4389 3356
rect 4370 3313 4373 3336
rect 4386 3296 4389 3353
rect 4394 3343 4397 3506
rect 4402 3403 4405 3553
rect 4410 3523 4413 3536
rect 4402 3333 4405 3366
rect 4354 3293 4365 3296
rect 4346 3273 4353 3276
rect 4350 3196 4353 3273
rect 4346 3193 4353 3196
rect 4346 3133 4349 3193
rect 4362 3176 4365 3293
rect 4354 3173 4365 3176
rect 4378 3293 4389 3296
rect 4378 3176 4381 3293
rect 4378 3173 4389 3176
rect 4354 3153 4357 3173
rect 4362 3133 4365 3146
rect 4346 2976 4349 3126
rect 4386 3123 4389 3173
rect 4394 3123 4397 3326
rect 4354 3086 4357 3106
rect 4410 3103 4413 3516
rect 4418 3383 4421 3556
rect 4426 3516 4429 3603
rect 4434 3523 4437 3576
rect 4458 3526 4461 3603
rect 4474 3543 4477 3616
rect 4482 3583 4485 3753
rect 4490 3733 4493 3746
rect 4490 3613 4493 3626
rect 4490 3533 4493 3606
rect 4498 3533 4501 3726
rect 4506 3553 4509 3736
rect 4514 3723 4517 3783
rect 4534 3766 4537 3823
rect 4534 3763 4541 3766
rect 4522 3723 4525 3736
rect 4530 3733 4533 3746
rect 4530 3713 4533 3726
rect 4538 3696 4541 3763
rect 4546 3733 4549 3816
rect 4558 3766 4561 3823
rect 4554 3763 4561 3766
rect 4582 3823 4589 3826
rect 4582 3766 4585 3823
rect 4582 3763 4589 3766
rect 4530 3693 4541 3696
rect 4426 3513 4437 3516
rect 4434 3456 4437 3513
rect 4434 3453 4441 3456
rect 4438 3386 4441 3453
rect 4450 3413 4453 3526
rect 4458 3523 4469 3526
rect 4466 3466 4469 3523
rect 4498 3513 4501 3526
rect 4506 3496 4509 3536
rect 4514 3526 4517 3636
rect 4530 3576 4533 3693
rect 4546 3676 4549 3706
rect 4542 3673 4549 3676
rect 4542 3596 4545 3673
rect 4542 3593 4549 3596
rect 4530 3573 4541 3576
rect 4522 3533 4525 3556
rect 4530 3533 4533 3546
rect 4514 3523 4533 3526
rect 4458 3463 4469 3466
rect 4502 3493 4509 3496
rect 4434 3383 4441 3386
rect 4434 3363 4437 3383
rect 4418 3323 4421 3336
rect 4426 3313 4429 3326
rect 4434 3246 4437 3336
rect 4442 3303 4445 3326
rect 4434 3243 4445 3246
rect 4434 3156 4437 3236
rect 4442 3216 4445 3243
rect 4450 3233 4453 3406
rect 4458 3366 4461 3463
rect 4482 3403 4485 3436
rect 4502 3426 4505 3493
rect 4498 3423 4505 3426
rect 4458 3363 4469 3366
rect 4466 3236 4469 3363
rect 4482 3316 4485 3336
rect 4478 3313 4485 3316
rect 4478 3246 4481 3313
rect 4478 3243 4485 3246
rect 4458 3233 4469 3236
rect 4442 3213 4449 3216
rect 4430 3153 4437 3156
rect 4430 3106 4433 3153
rect 4446 3146 4449 3213
rect 4442 3143 4449 3146
rect 4442 3113 4445 3143
rect 4430 3103 4437 3106
rect 4354 3083 4361 3086
rect 4322 2973 4333 2976
rect 4330 2856 4333 2973
rect 4322 2853 4333 2856
rect 4342 2973 4349 2976
rect 4322 2653 4325 2853
rect 4342 2836 4345 2973
rect 4358 2966 4361 3083
rect 4354 2963 4361 2966
rect 4330 2813 4333 2836
rect 4342 2833 4349 2836
rect 4306 2633 4317 2636
rect 4314 2566 4317 2633
rect 4330 2613 4333 2726
rect 4338 2613 4341 2816
rect 4346 2603 4349 2833
rect 4354 2763 4357 2963
rect 4370 2933 4373 3016
rect 4378 2993 4381 3006
rect 4386 2983 4389 3006
rect 4394 2996 4397 3016
rect 4402 3003 4405 3016
rect 4410 2996 4413 3006
rect 4394 2993 4413 2996
rect 4418 2936 4421 3026
rect 4378 2933 4389 2936
rect 4418 2933 4425 2936
rect 4362 2886 4365 2906
rect 4362 2883 4369 2886
rect 4366 2756 4369 2883
rect 4362 2753 4369 2756
rect 4306 2563 4317 2566
rect 4306 2533 4309 2563
rect 4314 2533 4317 2546
rect 4322 2543 4341 2546
rect 4290 2413 4301 2416
rect 4306 2413 4309 2526
rect 4314 2506 4317 2526
rect 4322 2523 4325 2543
rect 4314 2503 4321 2506
rect 4330 2503 4333 2536
rect 4338 2533 4341 2543
rect 4318 2436 4321 2503
rect 4338 2493 4341 2526
rect 4314 2433 4321 2436
rect 4290 2403 4293 2413
rect 4290 2303 4293 2376
rect 4194 2173 4213 2176
rect 4250 2193 4261 2196
rect 4266 2253 4273 2256
rect 4194 2096 4197 2173
rect 4210 2133 4213 2146
rect 4194 2093 4205 2096
rect 4186 2043 4193 2046
rect 4150 1963 4157 1966
rect 4162 2033 4177 2036
rect 4138 1943 4141 1956
rect 4138 1923 4141 1936
rect 4122 1913 4133 1916
rect 4082 1843 4093 1846
rect 4082 1733 4085 1843
rect 4106 1813 4109 1826
rect 4090 1793 4093 1806
rect 4090 1733 4093 1746
rect 4074 1723 4085 1726
rect 4098 1723 4101 1806
rect 4002 1613 4013 1616
rect 4018 1613 4021 1626
rect 3986 1603 3993 1606
rect 3990 1536 3993 1603
rect 4002 1543 4005 1606
rect 3990 1533 3997 1536
rect 3994 1476 3997 1533
rect 3994 1473 4001 1476
rect 3958 1433 3965 1436
rect 3958 1296 3961 1433
rect 3970 1343 3973 1416
rect 3970 1313 3973 1326
rect 3978 1323 3981 1436
rect 3986 1413 3989 1466
rect 3998 1406 4001 1473
rect 3994 1403 4001 1406
rect 3994 1366 3997 1403
rect 3990 1363 3997 1366
rect 3990 1306 3993 1363
rect 3990 1303 3997 1306
rect 3958 1293 3965 1296
rect 3962 1236 3965 1293
rect 3994 1286 3997 1303
rect 4010 1296 4013 1613
rect 4018 1566 4021 1606
rect 4034 1593 4037 1606
rect 4018 1563 4029 1566
rect 4026 1466 4029 1563
rect 4074 1536 4077 1716
rect 4082 1656 4085 1723
rect 4082 1653 4101 1656
rect 4082 1613 4085 1626
rect 4098 1566 4101 1653
rect 4070 1533 4077 1536
rect 4094 1563 4101 1566
rect 4018 1463 4029 1466
rect 4018 1433 4021 1463
rect 4058 1413 4061 1526
rect 4026 1393 4029 1406
rect 4018 1313 4021 1326
rect 4010 1293 4017 1296
rect 3994 1283 4005 1286
rect 3938 1233 3965 1236
rect 3938 1073 3941 1233
rect 3954 1213 3957 1226
rect 3962 1213 3973 1216
rect 3994 1213 3997 1226
rect 4002 1206 4005 1283
rect 3994 1203 4005 1206
rect 3946 1123 3949 1136
rect 3962 1123 3965 1146
rect 3970 1133 3973 1156
rect 3978 1133 3981 1146
rect 3926 1053 3941 1056
rect 3906 1003 3913 1006
rect 3866 933 3869 996
rect 3906 966 3909 1003
rect 3938 976 3941 1053
rect 3954 1013 3957 1116
rect 3978 1103 3981 1126
rect 3986 1113 3989 1126
rect 3978 1003 3981 1016
rect 3902 963 3909 966
rect 3930 973 3941 976
rect 3994 973 3997 1203
rect 4014 1166 4017 1293
rect 4034 1266 4037 1356
rect 4058 1333 4061 1396
rect 4070 1366 4073 1533
rect 4082 1463 4085 1526
rect 4070 1363 4077 1366
rect 4074 1296 4077 1363
rect 4094 1356 4097 1563
rect 4066 1293 4077 1296
rect 4086 1353 4097 1356
rect 4034 1263 4045 1266
rect 4042 1203 4045 1263
rect 4066 1236 4069 1293
rect 4086 1286 4089 1353
rect 4106 1333 4109 1756
rect 4114 1733 4117 1886
rect 4114 1713 4117 1726
rect 4114 1603 4117 1616
rect 4122 1613 4125 1816
rect 4130 1723 4133 1913
rect 4150 1846 4153 1963
rect 4150 1843 4157 1846
rect 4146 1813 4149 1826
rect 4138 1733 4141 1746
rect 4146 1706 4149 1766
rect 4138 1703 4149 1706
rect 4138 1636 4141 1703
rect 4138 1633 4149 1636
rect 4146 1613 4149 1633
rect 4154 1613 4157 1843
rect 4162 1773 4165 2033
rect 4170 2003 4173 2026
rect 4178 1933 4181 2006
rect 4190 1966 4193 2043
rect 4186 1963 4193 1966
rect 4186 1933 4189 1963
rect 4202 1946 4205 2093
rect 4194 1943 4205 1946
rect 4170 1733 4173 1926
rect 4194 1813 4197 1943
rect 4218 1933 4221 2016
rect 4226 1996 4229 2026
rect 4234 2013 4237 2126
rect 4250 2086 4253 2193
rect 4266 2166 4269 2253
rect 4298 2233 4301 2406
rect 4290 2193 4293 2226
rect 4266 2163 4285 2166
rect 4250 2083 4257 2086
rect 4226 1993 4233 1996
rect 4230 1926 4233 1993
rect 4226 1923 4233 1926
rect 4226 1863 4229 1923
rect 4194 1783 4197 1806
rect 4114 1513 4117 1536
rect 4122 1413 4125 1606
rect 4138 1546 4141 1606
rect 4146 1603 4157 1606
rect 4138 1543 4149 1546
rect 4130 1513 4133 1526
rect 4138 1496 4141 1536
rect 4134 1493 4141 1496
rect 4134 1406 4137 1493
rect 4134 1403 4141 1406
rect 4138 1383 4141 1403
rect 4146 1393 4149 1543
rect 4154 1366 4157 1526
rect 4162 1506 4165 1726
rect 4170 1623 4173 1726
rect 4178 1696 4181 1736
rect 4186 1713 4189 1726
rect 4202 1723 4205 1746
rect 4178 1693 4185 1696
rect 4182 1626 4185 1693
rect 4178 1623 4185 1626
rect 4170 1523 4173 1616
rect 4178 1603 4181 1623
rect 4162 1503 4169 1506
rect 4166 1436 4169 1503
rect 4194 1493 4197 1656
rect 4202 1613 4205 1626
rect 4210 1513 4213 1776
rect 4218 1753 4221 1806
rect 4218 1476 4221 1736
rect 4226 1576 4229 1746
rect 4234 1713 4237 1736
rect 4226 1573 4233 1576
rect 4210 1473 4221 1476
rect 4162 1433 4169 1436
rect 4162 1403 4165 1433
rect 4150 1363 4157 1366
rect 4170 1366 4173 1416
rect 4178 1413 4181 1466
rect 4178 1383 4181 1406
rect 4210 1396 4213 1473
rect 4230 1436 4233 1573
rect 4230 1433 4237 1436
rect 4226 1403 4229 1426
rect 4210 1393 4229 1396
rect 4170 1363 4177 1366
rect 4082 1283 4089 1286
rect 4066 1233 4077 1236
rect 4014 1163 4021 1166
rect 4018 1116 4021 1163
rect 4018 1113 4037 1116
rect 4010 993 4013 1016
rect 3882 933 3893 936
rect 3858 896 3861 916
rect 3858 893 3865 896
rect 3874 893 3877 926
rect 3890 913 3893 933
rect 3902 906 3905 963
rect 3882 903 3905 906
rect 3862 826 3865 893
rect 3858 823 3865 826
rect 3850 796 3853 816
rect 3858 803 3861 823
rect 3866 796 3869 806
rect 3850 793 3869 796
rect 3838 783 3845 786
rect 3802 703 3813 706
rect 3786 683 3797 686
rect 3778 603 3781 616
rect 3786 596 3789 676
rect 3794 603 3797 683
rect 3810 636 3813 703
rect 3802 633 3813 636
rect 3766 563 3773 566
rect 3778 593 3789 596
rect 3766 486 3769 563
rect 3766 483 3773 486
rect 3754 463 3765 466
rect 3722 403 3725 416
rect 3738 403 3741 416
rect 3706 353 3717 356
rect 3690 343 3709 346
rect 3690 323 3693 343
rect 3698 293 3701 336
rect 3706 333 3709 343
rect 3706 283 3709 326
rect 3586 243 3605 246
rect 3594 213 3597 236
rect 3602 206 3605 243
rect 3594 203 3605 206
rect 3634 243 3653 246
rect 3674 273 3685 276
rect 3634 203 3637 243
rect 3522 123 3525 146
rect 3570 133 3573 156
rect 3618 133 3621 196
rect 3642 123 3645 216
rect 3674 213 3677 273
rect 3714 266 3717 353
rect 3710 263 3717 266
rect 3710 146 3713 263
rect 3710 143 3717 146
rect 3714 123 3717 143
rect 3722 123 3725 326
rect 3730 213 3733 326
rect 3746 316 3749 376
rect 3754 323 3757 336
rect 3762 323 3765 463
rect 3770 333 3773 483
rect 3778 406 3781 593
rect 3786 413 3789 526
rect 3802 503 3805 633
rect 3826 616 3829 776
rect 3842 733 3845 783
rect 3826 613 3837 616
rect 3866 613 3869 726
rect 3818 413 3821 606
rect 3834 546 3837 613
rect 3882 606 3885 903
rect 3906 793 3909 816
rect 3922 813 3925 926
rect 3930 903 3933 973
rect 4010 966 4013 986
rect 4034 983 4037 1113
rect 4042 1103 4045 1126
rect 4066 1123 4069 1216
rect 4074 1203 4077 1233
rect 4082 1136 4085 1283
rect 4090 1203 4093 1226
rect 4130 1213 4133 1326
rect 4150 1316 4153 1363
rect 4146 1313 4153 1316
rect 4146 1216 4149 1313
rect 4174 1306 4177 1363
rect 4202 1333 4205 1356
rect 4170 1303 4177 1306
rect 4170 1286 4173 1303
rect 4162 1283 4173 1286
rect 4138 1213 4149 1216
rect 4154 1213 4157 1226
rect 4106 1193 4109 1206
rect 4138 1186 4141 1206
rect 4146 1203 4157 1206
rect 4130 1183 4141 1186
rect 4074 1133 4085 1136
rect 4058 1013 4061 1026
rect 4006 963 4013 966
rect 3938 836 3941 956
rect 3930 833 3941 836
rect 3922 696 3925 726
rect 3914 693 3925 696
rect 3890 613 3893 626
rect 3858 593 3861 606
rect 3882 603 3893 606
rect 3826 543 3837 546
rect 3858 543 3877 546
rect 3826 506 3829 543
rect 3858 533 3861 543
rect 3850 523 3861 526
rect 3826 503 3837 506
rect 3858 503 3861 523
rect 3866 513 3869 536
rect 3874 523 3877 543
rect 3834 446 3837 503
rect 3826 443 3837 446
rect 3826 413 3829 443
rect 3778 403 3789 406
rect 3850 403 3853 416
rect 3778 323 3781 396
rect 3746 313 3757 316
rect 3754 193 3757 313
rect 3786 283 3789 403
rect 3794 333 3797 346
rect 3826 336 3829 346
rect 3794 313 3797 326
rect 3802 323 3805 336
rect 3810 333 3821 336
rect 3826 333 3837 336
rect 3786 203 3789 216
rect 3802 123 3805 216
rect 3810 213 3813 326
rect 3834 316 3837 333
rect 3826 313 3837 316
rect 3826 296 3829 313
rect 3842 306 3845 326
rect 3834 303 3845 306
rect 3822 293 3829 296
rect 3822 236 3825 293
rect 3834 283 3837 296
rect 3850 283 3853 346
rect 3858 343 3877 346
rect 3890 343 3893 603
rect 3906 593 3909 616
rect 3914 603 3917 693
rect 3930 616 3933 833
rect 3946 803 3949 946
rect 3970 933 3973 946
rect 3978 886 3981 906
rect 3974 883 3981 886
rect 3974 746 3977 883
rect 3974 743 3981 746
rect 3986 743 3989 936
rect 3994 923 3997 936
rect 4006 916 4009 963
rect 4018 933 4021 976
rect 4018 923 4029 926
rect 4006 913 4013 916
rect 4010 856 4013 913
rect 4034 886 4037 936
rect 4026 883 4037 886
rect 4010 853 4017 856
rect 3994 813 3997 826
rect 3946 703 3949 736
rect 3978 726 3981 743
rect 3978 723 3985 726
rect 3926 613 3933 616
rect 3914 533 3917 546
rect 3898 503 3901 526
rect 3926 516 3929 613
rect 3914 513 3929 516
rect 3914 466 3917 513
rect 3938 506 3941 606
rect 3946 603 3949 616
rect 3970 593 3973 716
rect 3982 636 3985 723
rect 3994 713 3997 726
rect 4014 686 4017 853
rect 4026 813 4029 883
rect 4034 813 4037 826
rect 4026 723 4029 746
rect 4034 713 4037 726
rect 4042 703 4045 946
rect 4074 943 4077 1133
rect 4082 1006 4085 1126
rect 4090 1013 4093 1136
rect 4098 1053 4101 1136
rect 4098 1013 4101 1026
rect 4082 1003 4101 1006
rect 4106 986 4109 1126
rect 4098 983 4109 986
rect 4074 933 4085 936
rect 4050 906 4053 926
rect 4050 903 4061 906
rect 4058 836 4061 903
rect 4098 836 4101 983
rect 4114 946 4117 1106
rect 4130 1036 4133 1183
rect 4146 1046 4149 1196
rect 4154 1143 4157 1203
rect 4162 1133 4165 1283
rect 4186 1266 4189 1326
rect 4226 1296 4229 1393
rect 4234 1376 4237 1433
rect 4242 1393 4245 2046
rect 4254 1976 4257 2083
rect 4282 2046 4285 2163
rect 4266 2043 4285 2046
rect 4254 1973 4261 1976
rect 4250 1933 4253 1956
rect 4258 1943 4261 1973
rect 4250 1723 4253 1816
rect 4258 1763 4261 1926
rect 4266 1743 4269 2043
rect 4274 2013 4277 2036
rect 4306 1946 4309 2406
rect 4314 2373 4317 2433
rect 4322 2366 4325 2416
rect 4314 2363 4325 2366
rect 4338 2363 4341 2416
rect 4346 2383 4349 2586
rect 4354 2413 4357 2616
rect 4314 2333 4317 2363
rect 4330 2333 4333 2356
rect 4314 2213 4317 2236
rect 4330 2183 4333 2326
rect 4346 2213 4349 2346
rect 4354 2343 4357 2396
rect 4354 2313 4357 2326
rect 4362 2293 4365 2753
rect 4378 2736 4381 2926
rect 4394 2903 4397 2926
rect 4402 2813 4405 2836
rect 4410 2803 4413 2926
rect 4422 2866 4425 2933
rect 4418 2863 4425 2866
rect 4418 2843 4421 2863
rect 4418 2796 4421 2816
rect 4426 2803 4429 2816
rect 4434 2813 4437 3103
rect 4450 3013 4453 3126
rect 4442 2926 4445 2946
rect 4442 2923 4449 2926
rect 4446 2836 4449 2923
rect 4442 2833 4449 2836
rect 4434 2796 4437 2806
rect 4394 2783 4397 2796
rect 4370 2733 4381 2736
rect 4370 2686 4373 2733
rect 4378 2703 4381 2726
rect 4386 2686 4389 2766
rect 4410 2733 4413 2796
rect 4418 2793 4437 2796
rect 4442 2793 4445 2833
rect 4426 2733 4437 2736
rect 4426 2703 4429 2726
rect 4370 2683 4377 2686
rect 4386 2683 4405 2686
rect 4374 2626 4377 2683
rect 4374 2623 4381 2626
rect 4370 2386 4373 2596
rect 4378 2403 4381 2623
rect 4386 2613 4389 2666
rect 4370 2383 4377 2386
rect 4374 2286 4377 2383
rect 4370 2283 4377 2286
rect 4338 2193 4341 2206
rect 4354 2196 4357 2206
rect 4346 2193 4357 2196
rect 4362 2193 4365 2206
rect 4346 2173 4349 2193
rect 4346 2146 4349 2166
rect 4338 2143 4349 2146
rect 4314 1996 4317 2006
rect 4322 2003 4325 2126
rect 4338 2036 4341 2143
rect 4338 2033 4349 2036
rect 4330 1996 4333 2016
rect 4346 2013 4349 2033
rect 4314 1993 4333 1996
rect 4338 1993 4341 2006
rect 4306 1943 4317 1946
rect 4274 1863 4277 1926
rect 4282 1776 4285 1856
rect 4274 1773 4285 1776
rect 4258 1723 4261 1736
rect 4274 1706 4277 1773
rect 4270 1703 4277 1706
rect 4270 1636 4273 1703
rect 4270 1633 4277 1636
rect 4266 1526 4269 1616
rect 4250 1523 4269 1526
rect 4250 1413 4253 1523
rect 4250 1383 4253 1406
rect 4258 1393 4261 1516
rect 4274 1436 4277 1633
rect 4282 1533 4285 1766
rect 4298 1733 4301 1936
rect 4314 1876 4317 1943
rect 4310 1873 4317 1876
rect 4310 1746 4313 1873
rect 4330 1856 4333 1986
rect 4322 1853 4333 1856
rect 4346 1853 4349 2006
rect 4354 1933 4357 2186
rect 4370 2163 4373 2283
rect 4386 2213 4389 2606
rect 4394 2533 4397 2606
rect 4402 2593 4405 2683
rect 4434 2663 4437 2733
rect 4442 2723 4445 2776
rect 4450 2706 4453 2816
rect 4458 2786 4461 3233
rect 4466 3196 4469 3216
rect 4482 3203 4485 3243
rect 4466 3193 4473 3196
rect 4470 2976 4473 3193
rect 4490 3183 4493 3376
rect 4498 3213 4501 3423
rect 4506 3403 4509 3416
rect 4514 3373 4517 3516
rect 4530 3506 4533 3523
rect 4526 3503 4533 3506
rect 4526 3436 4529 3503
rect 4538 3446 4541 3573
rect 4546 3523 4549 3593
rect 4538 3443 4545 3446
rect 4526 3433 4533 3436
rect 4522 3353 4525 3406
rect 4506 3343 4525 3346
rect 4506 3323 4509 3343
rect 4514 3323 4517 3336
rect 4522 3333 4525 3343
rect 4530 3306 4533 3433
rect 4542 3346 4545 3443
rect 4554 3413 4557 3763
rect 4562 3743 4581 3746
rect 4562 3723 4565 3743
rect 4570 3703 4573 3736
rect 4578 3733 4581 3743
rect 4586 3733 4589 3763
rect 4586 3713 4589 3726
rect 4594 3723 4597 3816
rect 4602 3713 4605 3896
rect 4642 3893 4645 4143
rect 4658 3946 4661 4273
rect 4690 4186 4693 4326
rect 4650 3943 4661 3946
rect 4682 4183 4693 4186
rect 4650 3923 4653 3943
rect 4626 3736 4629 3816
rect 4642 3793 4645 3806
rect 4626 3733 4637 3736
rect 4618 3683 4621 3726
rect 4634 3636 4637 3733
rect 4650 3723 4653 3816
rect 4658 3723 4661 3736
rect 4666 3706 4669 3806
rect 4618 3633 4637 3636
rect 4662 3703 4669 3706
rect 4562 3506 4565 3566
rect 4570 3523 4573 3616
rect 4578 3533 4581 3546
rect 4594 3533 4597 3626
rect 4618 3563 4621 3633
rect 4662 3626 4665 3703
rect 4674 3633 4677 3926
rect 4682 3903 4685 4183
rect 4690 4113 4693 4126
rect 4706 4013 4709 4326
rect 4746 4213 4749 4326
rect 4730 4113 4733 4126
rect 4754 4123 4757 4216
rect 4738 3946 4741 4016
rect 4734 3943 4741 3946
rect 4682 3753 4685 3816
rect 4682 3723 4685 3746
rect 4634 3613 4645 3616
rect 4650 3613 4653 3626
rect 4662 3623 4669 3626
rect 4562 3503 4573 3506
rect 4522 3303 4533 3306
rect 4538 3343 4545 3346
rect 4522 3256 4525 3303
rect 4538 3296 4541 3343
rect 4570 3333 4573 3503
rect 4586 3406 4589 3526
rect 4602 3413 4605 3536
rect 4610 3523 4613 3546
rect 4618 3523 4621 3536
rect 4626 3506 4629 3586
rect 4618 3503 4629 3506
rect 4618 3436 4621 3503
rect 4618 3433 4629 3436
rect 4586 3403 4597 3406
rect 4546 3313 4549 3326
rect 4538 3293 4545 3296
rect 4522 3253 4533 3256
rect 4506 3213 4509 3236
rect 4490 3086 4493 3146
rect 4466 2973 4473 2976
rect 4482 3083 4493 3086
rect 4466 2803 4469 2973
rect 4482 2966 4485 3083
rect 4498 3066 4501 3206
rect 4530 3203 4533 3253
rect 4542 3226 4545 3293
rect 4554 3233 4557 3326
rect 4594 3323 4597 3403
rect 4538 3223 4545 3226
rect 4538 3143 4541 3223
rect 4586 3213 4589 3236
rect 4546 3193 4549 3206
rect 4562 3176 4565 3206
rect 4562 3173 4573 3176
rect 4494 3063 4501 3066
rect 4494 3006 4497 3063
rect 4506 3013 4509 3126
rect 4538 3123 4541 3136
rect 4570 3123 4573 3173
rect 4594 3146 4597 3316
rect 4610 3256 4613 3416
rect 4626 3376 4629 3433
rect 4634 3383 4637 3606
rect 4642 3403 4645 3546
rect 4650 3496 4653 3606
rect 4658 3553 4661 3606
rect 4666 3583 4669 3623
rect 4674 3603 4677 3626
rect 4658 3516 4661 3536
rect 4674 3533 4677 3546
rect 4666 3523 4677 3526
rect 4658 3513 4669 3516
rect 4650 3493 4657 3496
rect 4654 3426 4657 3493
rect 4654 3423 4661 3426
rect 4626 3373 4637 3376
rect 4634 3356 4637 3373
rect 4634 3353 4641 3356
rect 4638 3286 4641 3353
rect 4650 3323 4653 3416
rect 4658 3323 4661 3423
rect 4606 3253 4613 3256
rect 4634 3283 4641 3286
rect 4606 3176 4609 3253
rect 4606 3173 4613 3176
rect 4594 3143 4601 3146
rect 4598 3096 4601 3143
rect 4594 3093 4601 3096
rect 4494 3003 4501 3006
rect 4482 2963 4489 2966
rect 4486 2886 4489 2963
rect 4482 2883 4489 2886
rect 4458 2783 4465 2786
rect 4446 2703 4453 2706
rect 4446 2656 4449 2703
rect 4462 2696 4465 2783
rect 4418 2626 4421 2656
rect 4442 2653 4449 2656
rect 4458 2693 4465 2696
rect 4418 2623 4429 2626
rect 4410 2563 4413 2616
rect 4426 2576 4429 2623
rect 4442 2603 4445 2653
rect 4458 2616 4461 2693
rect 4458 2613 4465 2616
rect 4418 2573 4429 2576
rect 4418 2546 4421 2573
rect 4414 2543 4421 2546
rect 4394 2513 4397 2526
rect 4394 2403 4397 2416
rect 4402 2413 4405 2526
rect 4414 2466 4417 2543
rect 4434 2513 4437 2526
rect 4414 2463 4421 2466
rect 4410 2413 4413 2446
rect 4418 2423 4421 2463
rect 4402 2386 4405 2406
rect 4418 2393 4421 2406
rect 4426 2403 4429 2486
rect 4398 2383 4405 2386
rect 4398 2156 4401 2383
rect 4410 2203 4413 2386
rect 4418 2306 4421 2326
rect 4426 2323 4429 2336
rect 4418 2303 4425 2306
rect 4410 2183 4413 2196
rect 4398 2153 4405 2156
rect 4378 2133 4381 2146
rect 4402 2076 4405 2153
rect 4394 2073 4405 2076
rect 4362 2013 4365 2026
rect 4394 2006 4397 2073
rect 4394 2003 4405 2006
rect 4402 1983 4405 2003
rect 4410 1966 4413 2176
rect 4422 2146 4425 2303
rect 4434 2163 4437 2426
rect 4442 2423 4445 2596
rect 4442 2333 4445 2416
rect 4450 2363 4453 2606
rect 4462 2556 4465 2613
rect 4474 2583 4477 2816
rect 4482 2593 4485 2883
rect 4498 2846 4501 3003
rect 4530 2933 4533 2946
rect 4494 2843 4501 2846
rect 4494 2756 4497 2843
rect 4506 2813 4509 2926
rect 4530 2813 4533 2916
rect 4490 2753 4497 2756
rect 4490 2593 4493 2753
rect 4506 2743 4509 2806
rect 4546 2803 4549 3006
rect 4554 2913 4557 3016
rect 4562 2993 4565 3006
rect 4578 3003 4581 3056
rect 4570 2813 4573 2906
rect 4586 2903 4589 3016
rect 4594 2896 4597 3093
rect 4610 3026 4613 3173
rect 4618 3123 4621 3136
rect 4634 3086 4637 3283
rect 4642 3213 4645 3226
rect 4650 3136 4653 3206
rect 4626 3083 4637 3086
rect 4642 3133 4653 3136
rect 4658 3133 4661 3216
rect 4610 3023 4621 3026
rect 4602 2923 4605 3006
rect 4586 2893 4597 2896
rect 4586 2876 4589 2893
rect 4602 2886 4605 2916
rect 4582 2873 4589 2876
rect 4594 2883 4605 2886
rect 4562 2783 4565 2806
rect 4582 2776 4585 2873
rect 4582 2773 4589 2776
rect 4498 2696 4501 2736
rect 4498 2693 4509 2696
rect 4506 2626 4509 2693
rect 4498 2623 4509 2626
rect 4458 2553 4465 2556
rect 4458 2476 4461 2553
rect 4482 2533 4485 2556
rect 4498 2523 4501 2623
rect 4522 2606 4525 2746
rect 4554 2613 4557 2726
rect 4586 2693 4589 2773
rect 4514 2603 4525 2606
rect 4514 2533 4517 2603
rect 4458 2473 4469 2476
rect 4466 2386 4469 2473
rect 4498 2413 4501 2436
rect 4514 2413 4517 2526
rect 4562 2513 4565 2526
rect 4578 2493 4581 2636
rect 4586 2603 4589 2626
rect 4594 2586 4597 2883
rect 4610 2866 4613 3006
rect 4606 2863 4613 2866
rect 4606 2756 4609 2863
rect 4606 2753 4613 2756
rect 4610 2733 4613 2753
rect 4618 2733 4621 3023
rect 4626 2933 4629 3083
rect 4642 3013 4645 3133
rect 4650 2993 4653 3126
rect 4666 3116 4669 3513
rect 4682 3413 4685 3686
rect 4690 3593 4693 3806
rect 4698 3803 4701 3926
rect 4722 3913 4725 3926
rect 4722 3856 4725 3906
rect 4734 3876 4737 3943
rect 4762 3933 4765 3946
rect 4778 3943 4781 4383
rect 4786 4123 4789 4146
rect 4734 3873 4741 3876
rect 4718 3853 4725 3856
rect 4738 3856 4741 3873
rect 4738 3853 4749 3856
rect 4706 3793 4709 3816
rect 4718 3776 4721 3853
rect 4746 3776 4749 3853
rect 4718 3773 4725 3776
rect 4698 3733 4701 3746
rect 4722 3726 4725 3773
rect 4738 3773 4749 3776
rect 4698 3713 4701 3726
rect 4690 3523 4693 3536
rect 4698 3533 4701 3616
rect 4706 3613 4709 3726
rect 4722 3723 4729 3726
rect 4698 3423 4701 3526
rect 4706 3523 4709 3556
rect 4714 3516 4717 3716
rect 4726 3666 4729 3723
rect 4710 3513 4717 3516
rect 4722 3663 4729 3666
rect 4674 3393 4677 3406
rect 4682 3333 4685 3406
rect 4690 3376 4693 3416
rect 4698 3393 4701 3416
rect 4710 3406 4713 3513
rect 4706 3403 4713 3406
rect 4706 3383 4709 3403
rect 4690 3373 4717 3376
rect 4690 3343 4709 3346
rect 4674 3313 4677 3326
rect 4674 3193 4677 3216
rect 4682 3186 4685 3326
rect 4690 3323 4693 3343
rect 4698 3223 4701 3336
rect 4706 3333 4709 3343
rect 4706 3296 4709 3326
rect 4714 3323 4717 3373
rect 4722 3313 4725 3663
rect 4738 3456 4741 3773
rect 4746 3733 4749 3756
rect 4746 3706 4749 3726
rect 4762 3723 4765 3816
rect 4746 3703 4757 3706
rect 4754 3636 4757 3703
rect 4746 3633 4757 3636
rect 4746 3613 4749 3633
rect 4746 3523 4749 3536
rect 4738 3453 4745 3456
rect 4742 3376 4745 3453
rect 4754 3413 4757 3426
rect 4738 3373 4745 3376
rect 4706 3293 4717 3296
rect 4714 3216 4717 3293
rect 4662 3113 4669 3116
rect 4678 3183 4685 3186
rect 4698 3213 4717 3216
rect 4662 3046 4665 3113
rect 4678 3106 4681 3183
rect 4698 3136 4701 3213
rect 4698 3133 4705 3136
rect 4674 3103 4681 3106
rect 4662 3043 4669 3046
rect 4658 3013 4661 3026
rect 4658 2983 4661 3006
rect 4642 2943 4661 2946
rect 4626 2813 4629 2846
rect 4626 2793 4629 2806
rect 4634 2803 4637 2936
rect 4642 2923 4645 2943
rect 4650 2923 4653 2936
rect 4658 2933 4661 2943
rect 4642 2743 4645 2816
rect 4658 2813 4661 2926
rect 4650 2793 4653 2806
rect 4590 2583 4597 2586
rect 4590 2466 4593 2583
rect 4602 2556 4605 2726
rect 4610 2693 4613 2726
rect 4634 2716 4637 2736
rect 4626 2713 4637 2716
rect 4626 2626 4629 2713
rect 4610 2613 4613 2626
rect 4626 2623 4637 2626
rect 4602 2553 4621 2556
rect 4590 2463 4597 2466
rect 4458 2383 4469 2386
rect 4418 2143 4425 2146
rect 4418 2096 4421 2143
rect 4426 2113 4429 2126
rect 4418 2093 4425 2096
rect 4402 1963 4413 1966
rect 4378 1943 4381 1956
rect 4322 1786 4325 1853
rect 4338 1793 4341 1806
rect 4322 1783 4333 1786
rect 4306 1743 4313 1746
rect 4290 1713 4293 1726
rect 4290 1533 4293 1596
rect 4274 1433 4285 1436
rect 4274 1413 4277 1426
rect 4282 1406 4285 1433
rect 4290 1413 4293 1436
rect 4274 1403 4285 1406
rect 4298 1403 4301 1536
rect 4234 1373 4241 1376
rect 4178 1263 4189 1266
rect 4218 1293 4229 1296
rect 4170 1133 4173 1236
rect 4178 1133 4181 1263
rect 4186 1193 4189 1216
rect 4194 1186 4197 1216
rect 4190 1183 4197 1186
rect 4146 1043 4157 1046
rect 4130 1033 4141 1036
rect 4110 943 4117 946
rect 4110 856 4113 943
rect 4110 853 4117 856
rect 4050 833 4061 836
rect 4050 776 4053 833
rect 4058 793 4061 816
rect 4050 773 4057 776
rect 4054 696 4057 773
rect 4066 726 4069 806
rect 4074 796 4077 806
rect 4082 803 4085 836
rect 4098 833 4109 836
rect 4090 796 4093 816
rect 4074 793 4093 796
rect 4098 773 4101 806
rect 4074 743 4093 746
rect 4074 733 4077 743
rect 4066 723 4077 726
rect 4082 723 4085 736
rect 4090 723 4093 743
rect 4098 733 4101 756
rect 4074 713 4077 723
rect 3978 633 3985 636
rect 4010 683 4017 686
rect 4050 693 4057 696
rect 3978 603 3981 633
rect 3954 533 3957 546
rect 3930 503 3941 506
rect 3946 506 3949 526
rect 3978 506 3981 576
rect 3946 503 3957 506
rect 3914 463 3925 466
rect 3898 413 3901 426
rect 3922 376 3925 463
rect 3930 413 3933 503
rect 3954 426 3957 503
rect 3938 413 3941 426
rect 3946 423 3957 426
rect 3970 503 3981 506
rect 3970 426 3973 503
rect 3970 423 3981 426
rect 3946 403 3949 423
rect 3910 373 3925 376
rect 3858 323 3861 343
rect 3866 293 3869 336
rect 3874 333 3877 343
rect 3890 333 3901 336
rect 3874 283 3877 326
rect 3834 256 3837 276
rect 3834 253 3841 256
rect 3822 233 3829 236
rect 3826 213 3829 233
rect 3838 206 3841 253
rect 3882 213 3885 326
rect 3898 313 3901 326
rect 3910 306 3913 373
rect 3970 336 3973 406
rect 3922 333 3941 336
rect 3906 303 3913 306
rect 3834 203 3841 206
rect 3906 203 3909 303
rect 3930 273 3933 333
rect 3946 326 3949 336
rect 3962 333 3973 336
rect 3978 333 3981 423
rect 3986 413 3989 616
rect 3994 603 3997 616
rect 4010 586 4013 683
rect 4042 613 4045 646
rect 4002 583 4013 586
rect 4002 426 4005 583
rect 4002 423 4013 426
rect 4010 403 4013 423
rect 4018 413 4021 596
rect 4026 513 4029 586
rect 4034 566 4037 606
rect 4050 583 4053 693
rect 4034 563 4045 566
rect 4042 506 4045 563
rect 4058 533 4061 616
rect 4066 573 4069 706
rect 4106 683 4109 833
rect 4074 613 4077 626
rect 4114 623 4117 853
rect 4122 723 4125 936
rect 4130 913 4133 1016
rect 4138 933 4141 1033
rect 4154 956 4157 1043
rect 4170 1013 4173 1126
rect 4178 1013 4181 1126
rect 4190 1076 4193 1183
rect 4202 1096 4205 1206
rect 4218 1203 4221 1293
rect 4238 1286 4241 1373
rect 4250 1313 4253 1326
rect 4234 1283 4241 1286
rect 4218 1123 4221 1136
rect 4226 1113 4229 1216
rect 4234 1213 4237 1283
rect 4258 1213 4261 1226
rect 4234 1133 4237 1206
rect 4242 1203 4253 1206
rect 4250 1186 4253 1203
rect 4266 1193 4269 1216
rect 4250 1183 4261 1186
rect 4242 1103 4245 1126
rect 4258 1123 4261 1183
rect 4266 1133 4269 1146
rect 4274 1106 4277 1403
rect 4282 1303 4285 1326
rect 4290 1313 4293 1326
rect 4298 1213 4301 1226
rect 4266 1103 4277 1106
rect 4202 1093 4213 1096
rect 4186 1073 4193 1076
rect 4186 1006 4189 1073
rect 4194 1013 4197 1056
rect 4210 1036 4213 1093
rect 4202 1033 4213 1036
rect 4202 1013 4205 1033
rect 4146 953 4157 956
rect 4146 923 4149 953
rect 4130 693 4133 816
rect 4146 733 4149 746
rect 4090 603 4093 616
rect 4138 613 4141 636
rect 4154 606 4157 726
rect 4162 676 4165 936
rect 4170 813 4173 1006
rect 4182 1003 4189 1006
rect 4266 1006 4269 1103
rect 4282 1013 4285 1126
rect 4290 1123 4293 1136
rect 4306 1083 4309 1743
rect 4314 1703 4317 1726
rect 4314 1516 4317 1646
rect 4322 1533 4325 1616
rect 4314 1513 4321 1516
rect 4330 1513 4333 1783
rect 4362 1723 4365 1816
rect 4378 1716 4381 1936
rect 4402 1866 4405 1963
rect 4422 1946 4425 2093
rect 4422 1943 4429 1946
rect 4402 1863 4409 1866
rect 4406 1766 4409 1863
rect 4406 1763 4413 1766
rect 4386 1743 4405 1746
rect 4386 1733 4389 1743
rect 4394 1723 4397 1736
rect 4402 1723 4405 1743
rect 4370 1713 4381 1716
rect 4346 1583 4349 1606
rect 4318 1456 4321 1513
rect 4314 1453 4321 1456
rect 4314 1403 4317 1453
rect 4338 1436 4341 1556
rect 4370 1553 4373 1713
rect 4378 1626 4381 1706
rect 4378 1623 4385 1626
rect 4382 1556 4385 1623
rect 4394 1613 4397 1626
rect 4378 1553 4385 1556
rect 4346 1543 4373 1546
rect 4346 1533 4349 1543
rect 4354 1523 4357 1536
rect 4378 1506 4381 1553
rect 4370 1503 4381 1506
rect 4370 1446 4373 1503
rect 4386 1456 4389 1536
rect 4410 1533 4413 1763
rect 4418 1733 4421 1936
rect 4418 1703 4421 1726
rect 4426 1646 4429 1943
rect 4434 1933 4437 2016
rect 4434 1876 4437 1926
rect 4442 1896 4445 2216
rect 4458 2213 4461 2383
rect 4490 2373 4493 2406
rect 4546 2403 4549 2416
rect 4466 2313 4469 2326
rect 4482 2296 4485 2366
rect 4482 2293 4493 2296
rect 4466 2213 4477 2216
rect 4490 2213 4493 2293
rect 4506 2223 4509 2336
rect 4538 2296 4541 2376
rect 4546 2333 4549 2386
rect 4530 2293 4541 2296
rect 4530 2226 4533 2293
rect 4554 2243 4557 2446
rect 4562 2403 4565 2426
rect 4530 2223 4541 2226
rect 4466 2143 4469 2206
rect 4482 2186 4485 2206
rect 4530 2193 4533 2206
rect 4482 2183 4489 2186
rect 4450 2133 4469 2136
rect 4450 2086 4453 2133
rect 4458 2093 4461 2126
rect 4466 2113 4469 2126
rect 4450 2083 4469 2086
rect 4450 2013 4453 2066
rect 4466 2013 4469 2083
rect 4474 2063 4477 2166
rect 4486 2116 4489 2183
rect 4506 2146 4509 2156
rect 4498 2126 4501 2146
rect 4506 2143 4517 2146
rect 4522 2143 4525 2156
rect 4498 2123 4505 2126
rect 4482 2113 4489 2116
rect 4482 2056 4485 2113
rect 4474 2053 4485 2056
rect 4450 1996 4453 2006
rect 4458 2003 4469 2006
rect 4450 1993 4469 1996
rect 4458 1933 4461 1956
rect 4450 1913 4453 1926
rect 4466 1923 4469 1993
rect 4442 1893 4453 1896
rect 4434 1873 4441 1876
rect 4438 1796 4441 1873
rect 4434 1793 4441 1796
rect 4434 1706 4437 1793
rect 4450 1776 4453 1893
rect 4474 1836 4477 2053
rect 4482 2013 4485 2036
rect 4490 1966 4493 2096
rect 4482 1963 4493 1966
rect 4482 1933 4485 1963
rect 4502 1956 4505 2123
rect 4498 1953 4505 1956
rect 4498 1933 4501 1953
rect 4514 1936 4517 2143
rect 4538 2133 4541 2223
rect 4546 2186 4549 2206
rect 4562 2203 4565 2336
rect 4570 2286 4573 2416
rect 4586 2413 4589 2446
rect 4578 2403 4589 2406
rect 4586 2323 4589 2336
rect 4570 2283 4581 2286
rect 4570 2203 4573 2216
rect 4546 2183 4553 2186
rect 4538 2106 4541 2126
rect 4530 2103 4541 2106
rect 4530 1976 4533 2103
rect 4550 2096 4553 2183
rect 4578 2166 4581 2283
rect 4586 2193 4589 2206
rect 4594 2176 4597 2463
rect 4602 2413 4605 2526
rect 4610 2523 4613 2546
rect 4618 2516 4621 2553
rect 4634 2533 4637 2623
rect 4626 2523 4637 2526
rect 4610 2513 4621 2516
rect 4602 2393 4605 2406
rect 4610 2376 4613 2513
rect 4642 2503 4645 2736
rect 4658 2706 4661 2726
rect 4654 2703 4661 2706
rect 4654 2636 4657 2703
rect 4654 2633 4661 2636
rect 4606 2373 4613 2376
rect 4606 2266 4609 2373
rect 4606 2263 4613 2266
rect 4570 2163 4581 2166
rect 4590 2173 4597 2176
rect 4546 2093 4553 2096
rect 4530 1973 4541 1976
rect 4510 1933 4517 1936
rect 4510 1856 4513 1933
rect 4510 1853 4517 1856
rect 4466 1833 4477 1836
rect 4466 1786 4469 1833
rect 4490 1793 4493 1806
rect 4514 1796 4517 1853
rect 4522 1806 4525 1946
rect 4530 1943 4533 1956
rect 4538 1926 4541 1973
rect 4534 1923 4541 1926
rect 4534 1846 4537 1923
rect 4546 1853 4549 2093
rect 4554 1886 4557 1926
rect 4562 1906 4565 2136
rect 4570 2106 4573 2163
rect 4578 2133 4581 2156
rect 4570 2103 4581 2106
rect 4570 1913 4573 1936
rect 4562 1903 4573 1906
rect 4578 1903 4581 2103
rect 4590 1976 4593 2173
rect 4590 1973 4597 1976
rect 4586 1933 4589 1956
rect 4554 1883 4561 1886
rect 4534 1843 4541 1846
rect 4530 1813 4533 1826
rect 4522 1803 4533 1806
rect 4514 1793 4525 1796
rect 4466 1783 4477 1786
rect 4442 1773 4453 1776
rect 4442 1743 4445 1773
rect 4442 1723 4445 1736
rect 4466 1733 4469 1756
rect 4474 1716 4477 1783
rect 4522 1766 4525 1793
rect 4514 1763 4525 1766
rect 4466 1713 4477 1716
rect 4434 1703 4445 1706
rect 4418 1643 4429 1646
rect 4386 1453 4393 1456
rect 4370 1443 4381 1446
rect 4322 1433 4341 1436
rect 4322 1046 4325 1433
rect 4338 1323 4341 1426
rect 4378 1423 4381 1443
rect 4346 1343 4365 1346
rect 4346 1333 4349 1343
rect 4354 1303 4357 1336
rect 4362 1323 4365 1343
rect 4378 1323 4381 1396
rect 4390 1366 4393 1453
rect 4386 1363 4393 1366
rect 4386 1303 4389 1363
rect 4394 1333 4397 1346
rect 4346 1156 4349 1206
rect 4370 1186 4373 1206
rect 4338 1153 4349 1156
rect 4354 1183 4373 1186
rect 4338 1073 4341 1153
rect 4322 1043 4329 1046
rect 4266 1003 4277 1006
rect 4182 836 4185 1003
rect 4274 983 4277 1003
rect 4202 886 4205 956
rect 4202 883 4213 886
rect 4250 883 4253 926
rect 4290 906 4293 926
rect 4282 903 4293 906
rect 4178 833 4185 836
rect 4170 713 4173 736
rect 4178 703 4181 833
rect 4186 723 4189 816
rect 4210 803 4213 883
rect 4226 813 4229 856
rect 4282 846 4285 903
rect 4306 896 4309 1016
rect 4326 956 4329 1043
rect 4326 953 4333 956
rect 4302 893 4309 896
rect 4282 843 4293 846
rect 4218 706 4221 786
rect 4226 743 4245 746
rect 4226 733 4229 743
rect 4234 723 4237 736
rect 4242 723 4245 743
rect 4202 703 4221 706
rect 4162 673 4173 676
rect 4170 613 4173 673
rect 4178 613 4181 636
rect 4154 603 4181 606
rect 4034 503 4045 506
rect 4034 413 4037 503
rect 4090 413 4093 526
rect 4138 436 4141 536
rect 4146 523 4149 546
rect 4154 533 4157 596
rect 4202 566 4205 703
rect 4226 636 4229 706
rect 4250 653 4253 806
rect 4258 733 4261 746
rect 4258 693 4261 726
rect 4266 723 4269 816
rect 4274 796 4277 816
rect 4282 813 4285 826
rect 4274 793 4281 796
rect 4278 736 4281 793
rect 4290 743 4293 843
rect 4302 836 4305 893
rect 4302 833 4309 836
rect 4298 783 4301 816
rect 4306 763 4309 833
rect 4314 813 4317 886
rect 4330 853 4333 953
rect 4338 886 4341 1066
rect 4346 906 4349 1086
rect 4354 1013 4357 1183
rect 4386 1013 4389 1126
rect 4394 1063 4397 1326
rect 4370 976 4373 996
rect 4370 973 4377 976
rect 4354 913 4357 926
rect 4346 903 4357 906
rect 4338 883 4345 886
rect 4330 803 4333 826
rect 4342 776 4345 883
rect 4338 773 4345 776
rect 4338 753 4341 773
rect 4274 733 4281 736
rect 4274 716 4277 733
rect 4306 723 4317 726
rect 4322 723 4325 736
rect 4266 713 4277 716
rect 4218 633 4229 636
rect 4218 586 4221 633
rect 4218 583 4229 586
rect 4202 563 4221 566
rect 4162 523 4165 536
rect 4138 433 4149 436
rect 4026 356 4029 406
rect 4114 403 4117 416
rect 4026 353 4037 356
rect 3938 323 3949 326
rect 3954 306 3957 326
rect 3946 303 3957 306
rect 3946 226 3949 303
rect 3946 223 3957 226
rect 3834 133 3837 203
rect 3898 133 3901 146
rect 3930 123 3933 216
rect 3954 203 3957 223
rect 3962 126 3965 333
rect 3970 263 3973 326
rect 3994 313 3997 336
rect 4002 333 4013 336
rect 4002 213 4005 326
rect 4018 323 4021 336
rect 4034 333 4037 353
rect 4026 313 4029 326
rect 4042 303 4045 326
rect 4050 313 4053 386
rect 4106 346 4109 376
rect 4106 343 4117 346
rect 4058 213 4061 336
rect 4082 296 4085 336
rect 4114 296 4117 343
rect 4130 323 4133 416
rect 4146 346 4149 433
rect 4146 343 4153 346
rect 4074 293 4085 296
rect 4106 293 4117 296
rect 3978 193 3981 206
rect 4018 133 4021 156
rect 3962 123 3981 126
rect 4066 123 4069 216
rect 4074 193 4077 293
rect 4082 213 4085 256
rect 4082 196 4085 206
rect 4090 203 4093 276
rect 4098 196 4101 216
rect 4082 193 4101 196
rect 4106 123 4109 293
rect 4150 286 4153 343
rect 4170 336 4173 536
rect 4178 513 4181 526
rect 4194 413 4197 546
rect 4202 513 4205 526
rect 4218 496 4221 563
rect 4210 493 4221 496
rect 4210 426 4213 493
rect 4210 423 4221 426
rect 4162 333 4173 336
rect 4162 323 4165 333
rect 4170 303 4173 326
rect 4186 323 4189 406
rect 4194 373 4197 406
rect 4218 403 4221 423
rect 4226 403 4229 583
rect 4234 516 4237 576
rect 4242 566 4245 616
rect 4266 586 4269 713
rect 4314 706 4317 723
rect 4330 716 4333 736
rect 4310 703 4317 706
rect 4322 713 4333 716
rect 4262 583 4269 586
rect 4242 563 4253 566
rect 4234 513 4241 516
rect 4238 456 4241 513
rect 4234 453 4241 456
rect 4234 383 4237 453
rect 4250 436 4253 563
rect 4262 516 4265 583
rect 4274 526 4277 656
rect 4310 626 4313 703
rect 4290 613 4293 626
rect 4310 623 4317 626
rect 4314 606 4317 623
rect 4322 613 4325 713
rect 4330 613 4333 626
rect 4314 603 4333 606
rect 4282 533 4285 556
rect 4274 523 4285 526
rect 4262 513 4269 516
rect 4242 433 4253 436
rect 4194 323 4197 336
rect 4146 283 4153 286
rect 4114 213 4117 266
rect 4130 123 4133 206
rect 4146 203 4149 283
rect 4202 236 4205 366
rect 4218 303 4221 326
rect 4234 306 4237 326
rect 4230 303 4237 306
rect 4178 233 4205 236
rect 4230 236 4233 303
rect 4230 233 4237 236
rect 4154 196 4157 216
rect 4162 203 4165 216
rect 4178 213 4181 233
rect 4170 196 4173 206
rect 4154 193 4173 196
rect 4186 123 4189 216
rect 4202 193 4205 216
rect 4234 213 4237 233
rect 4242 206 4245 433
rect 4250 253 4253 416
rect 4266 413 4269 513
rect 4274 393 4277 406
rect 4258 343 4277 346
rect 4282 343 4285 523
rect 4290 506 4293 526
rect 4290 503 4301 506
rect 4298 436 4301 503
rect 4290 433 4301 436
rect 4290 413 4293 433
rect 4322 426 4325 546
rect 4322 423 4329 426
rect 4258 333 4261 343
rect 4258 313 4261 326
rect 4266 323 4269 336
rect 4274 323 4277 343
rect 4282 213 4285 336
rect 4290 303 4293 406
rect 4298 393 4301 406
rect 4314 403 4317 416
rect 4306 323 4309 386
rect 4314 333 4317 396
rect 4326 356 4329 423
rect 4338 373 4341 726
rect 4346 613 4349 636
rect 4354 393 4357 903
rect 4374 886 4377 973
rect 4386 923 4389 946
rect 4402 936 4405 1526
rect 4410 1513 4413 1526
rect 4418 1376 4421 1643
rect 4442 1636 4445 1703
rect 4466 1656 4469 1713
rect 4466 1653 4477 1656
rect 4426 1533 4429 1636
rect 4442 1633 4461 1636
rect 4434 1613 4437 1626
rect 4442 1566 4445 1616
rect 4438 1563 4445 1566
rect 4438 1496 4441 1563
rect 4458 1556 4461 1633
rect 4474 1573 4477 1653
rect 4450 1553 4461 1556
rect 4438 1493 4445 1496
rect 4442 1433 4445 1493
rect 4410 1373 4421 1376
rect 4410 1206 4413 1373
rect 4426 1333 4429 1356
rect 4450 1246 4453 1553
rect 4458 1533 4477 1536
rect 4482 1533 4485 1746
rect 4490 1613 4493 1706
rect 4514 1656 4517 1763
rect 4530 1746 4533 1803
rect 4526 1743 4533 1746
rect 4526 1676 4529 1743
rect 4526 1673 4533 1676
rect 4514 1653 4525 1656
rect 4490 1596 4493 1606
rect 4498 1603 4501 1636
rect 4506 1596 4509 1616
rect 4490 1593 4509 1596
rect 4514 1593 4517 1606
rect 4458 1393 4461 1533
rect 4466 1506 4469 1526
rect 4466 1503 4473 1506
rect 4470 1436 4473 1503
rect 4482 1493 4485 1526
rect 4466 1433 4473 1436
rect 4466 1336 4469 1433
rect 4458 1333 4469 1336
rect 4458 1306 4461 1333
rect 4466 1313 4469 1326
rect 4458 1303 4465 1306
rect 4418 1213 4421 1226
rect 4410 1203 4421 1206
rect 4418 1166 4421 1203
rect 4418 1163 4425 1166
rect 4422 1106 4425 1163
rect 4418 1103 4425 1106
rect 4402 933 4409 936
rect 4394 913 4397 926
rect 4370 883 4377 886
rect 4370 763 4373 883
rect 4322 353 4329 356
rect 4322 323 4325 353
rect 4370 346 4373 756
rect 4378 723 4381 776
rect 4386 733 4389 796
rect 4394 706 4397 896
rect 4406 886 4409 933
rect 4402 883 4409 886
rect 4402 766 4405 883
rect 4418 866 4421 1103
rect 4434 1086 4437 1246
rect 4442 1243 4453 1246
rect 4462 1246 4465 1303
rect 4462 1243 4469 1246
rect 4474 1243 4477 1416
rect 4482 1396 4485 1486
rect 4490 1403 4493 1536
rect 4498 1483 4501 1536
rect 4482 1393 4493 1396
rect 4490 1303 4493 1393
rect 4442 1193 4445 1243
rect 4450 1213 4453 1236
rect 4458 1213 4461 1226
rect 4466 1186 4469 1243
rect 4410 863 4421 866
rect 4430 1083 4437 1086
rect 4446 1183 4469 1186
rect 4430 866 4433 1083
rect 4446 1076 4449 1183
rect 4442 1073 4449 1076
rect 4430 863 4437 866
rect 4410 793 4413 863
rect 4418 813 4421 826
rect 4402 763 4413 766
rect 4402 733 4405 746
rect 4410 726 4413 763
rect 4386 703 4397 706
rect 4402 723 4413 726
rect 4386 636 4389 703
rect 4386 633 4397 636
rect 4378 543 4381 616
rect 4386 533 4389 606
rect 4394 603 4397 633
rect 4386 516 4389 526
rect 4394 523 4397 536
rect 4402 533 4405 723
rect 4410 613 4413 656
rect 4410 516 4413 606
rect 4426 583 4429 766
rect 4434 723 4437 863
rect 4442 786 4445 1073
rect 4458 946 4461 1136
rect 4474 1023 4477 1216
rect 4482 1196 4485 1206
rect 4490 1203 4493 1236
rect 4498 1223 4501 1416
rect 4506 1413 4509 1426
rect 4506 1323 4509 1406
rect 4514 1333 4517 1546
rect 4522 1533 4525 1653
rect 4530 1603 4533 1673
rect 4530 1543 4533 1556
rect 4538 1483 4541 1843
rect 4558 1796 4561 1883
rect 4554 1793 4561 1796
rect 4554 1736 4557 1793
rect 4570 1776 4573 1903
rect 4578 1813 4581 1826
rect 4546 1733 4557 1736
rect 4562 1773 4573 1776
rect 4562 1733 4565 1773
rect 4578 1756 4581 1806
rect 4570 1753 4581 1756
rect 4546 1716 4549 1733
rect 4554 1723 4565 1726
rect 4570 1723 4573 1753
rect 4546 1713 4557 1716
rect 4546 1476 4549 1686
rect 4538 1473 4549 1476
rect 4538 1416 4541 1473
rect 4522 1333 4525 1416
rect 4530 1413 4541 1416
rect 4546 1413 4549 1426
rect 4530 1333 4533 1396
rect 4538 1343 4541 1406
rect 4554 1396 4557 1713
rect 4578 1706 4581 1746
rect 4574 1703 4581 1706
rect 4574 1656 4577 1703
rect 4586 1666 4589 1856
rect 4594 1683 4597 1973
rect 4602 1923 4605 2246
rect 4610 2203 4613 2263
rect 4618 2146 4621 2496
rect 4626 2403 4629 2416
rect 4634 2403 4645 2406
rect 4626 2213 4629 2396
rect 4634 2286 4637 2403
rect 4650 2393 4653 2616
rect 4658 2493 4661 2633
rect 4658 2403 4661 2416
rect 4642 2343 4661 2346
rect 4642 2323 4645 2343
rect 4650 2323 4653 2336
rect 4658 2333 4661 2343
rect 4658 2306 4661 2326
rect 4654 2303 4661 2306
rect 4634 2283 4645 2286
rect 4642 2236 4645 2283
rect 4634 2233 4645 2236
rect 4654 2236 4657 2303
rect 4654 2233 4661 2236
rect 4634 2203 4637 2233
rect 4642 2196 4645 2216
rect 4650 2203 4653 2216
rect 4658 2213 4661 2233
rect 4658 2196 4661 2206
rect 4642 2193 4661 2196
rect 4618 2143 4629 2146
rect 4618 2123 4621 2136
rect 4618 1906 4621 2116
rect 4626 2056 4629 2143
rect 4642 2143 4661 2146
rect 4634 2066 4637 2136
rect 4642 2123 4645 2143
rect 4650 2123 4653 2136
rect 4658 2133 4661 2143
rect 4634 2063 4653 2066
rect 4626 2053 4637 2056
rect 4610 1903 4621 1906
rect 4610 1836 4613 1903
rect 4610 1833 4621 1836
rect 4602 1743 4605 1806
rect 4610 1726 4613 1816
rect 4606 1723 4613 1726
rect 4586 1663 4597 1666
rect 4574 1653 4581 1656
rect 4562 1533 4565 1626
rect 4570 1583 4573 1596
rect 4550 1393 4557 1396
rect 4514 1313 4517 1326
rect 4498 1196 4501 1216
rect 4482 1193 4501 1196
rect 4506 1173 4509 1306
rect 4514 1133 4517 1206
rect 4522 1203 4525 1236
rect 4530 1186 4533 1216
rect 4526 1183 4533 1186
rect 4490 1106 4493 1126
rect 4526 1116 4529 1183
rect 4522 1113 4529 1116
rect 4490 1103 4501 1106
rect 4498 1046 4501 1103
rect 4490 1043 4501 1046
rect 4466 993 4469 1006
rect 4474 1003 4477 1016
rect 4482 993 4485 1016
rect 4490 1003 4493 1043
rect 4458 943 4469 946
rect 4458 913 4461 936
rect 4450 793 4453 816
rect 4458 813 4461 826
rect 4466 813 4469 943
rect 4474 853 4477 936
rect 4490 933 4493 946
rect 4482 913 4485 926
rect 4498 923 4501 1026
rect 4522 946 4525 1113
rect 4538 1096 4541 1336
rect 4550 1236 4553 1393
rect 4550 1233 4557 1236
rect 4534 1093 4541 1096
rect 4534 966 4537 1093
rect 4534 963 4541 966
rect 4522 943 4533 946
rect 4522 906 4525 926
rect 4514 903 4525 906
rect 4514 836 4517 903
rect 4514 833 4525 836
rect 4442 783 4453 786
rect 4450 736 4453 783
rect 4446 733 4453 736
rect 4446 656 4449 733
rect 4446 653 4453 656
rect 4450 606 4453 653
rect 4458 613 4461 726
rect 4474 633 4477 816
rect 4490 796 4493 806
rect 4498 803 4501 816
rect 4506 796 4509 816
rect 4490 793 4509 796
rect 4514 793 4517 806
rect 4482 743 4501 746
rect 4482 733 4485 743
rect 4490 656 4493 736
rect 4498 723 4501 743
rect 4490 653 4497 656
rect 4450 603 4461 606
rect 4458 566 4461 603
rect 4494 576 4497 653
rect 4506 613 4509 736
rect 4522 726 4525 833
rect 4530 813 4533 943
rect 4514 723 4525 726
rect 4514 653 4517 723
rect 4538 646 4541 963
rect 4546 906 4549 1216
rect 4554 1203 4557 1233
rect 4562 1223 4565 1526
rect 4570 1416 4573 1536
rect 4578 1426 4581 1653
rect 4594 1586 4597 1663
rect 4606 1646 4609 1723
rect 4606 1643 4613 1646
rect 4610 1623 4613 1643
rect 4586 1583 4597 1586
rect 4586 1543 4589 1583
rect 4586 1493 4589 1536
rect 4594 1533 4597 1556
rect 4602 1513 4605 1566
rect 4610 1426 4613 1616
rect 4618 1613 4621 1833
rect 4626 1703 4629 1906
rect 4634 1813 4637 2053
rect 4642 1933 4645 1946
rect 4650 1906 4653 2063
rect 4658 2033 4661 2126
rect 4666 2086 4669 3043
rect 4674 2826 4677 3103
rect 4682 2996 4685 3016
rect 4690 3013 4693 3126
rect 4702 3036 4705 3133
rect 4698 3033 4705 3036
rect 4698 3013 4701 3033
rect 4730 3023 4733 3126
rect 4714 2996 4717 3016
rect 4722 3003 4725 3016
rect 4730 2996 4733 3006
rect 4682 2993 4689 2996
rect 4714 2993 4733 2996
rect 4686 2866 4689 2993
rect 4698 2913 4701 2926
rect 4706 2923 4717 2926
rect 4682 2863 4689 2866
rect 4682 2843 4685 2863
rect 4714 2826 4717 2846
rect 4674 2823 4685 2826
rect 4682 2766 4685 2823
rect 4706 2823 4717 2826
rect 4706 2776 4709 2823
rect 4706 2773 4717 2776
rect 4674 2763 4685 2766
rect 4674 2706 4677 2763
rect 4714 2756 4717 2773
rect 4738 2766 4741 3373
rect 4754 3213 4757 3326
rect 4734 2763 4741 2766
rect 4714 2753 4725 2756
rect 4682 2743 4701 2746
rect 4682 2723 4685 2743
rect 4674 2703 4681 2706
rect 4678 2636 4681 2703
rect 4690 2686 4693 2736
rect 4698 2733 4701 2743
rect 4690 2683 4701 2686
rect 4674 2633 4681 2636
rect 4674 2613 4677 2633
rect 4674 2513 4677 2526
rect 4682 2523 4685 2536
rect 4674 2413 4677 2456
rect 4690 2423 4693 2526
rect 4674 2393 4677 2406
rect 4674 2276 4677 2376
rect 4682 2296 4685 2406
rect 4690 2323 4693 2416
rect 4698 2383 4701 2683
rect 4706 2633 4709 2726
rect 4722 2666 4725 2753
rect 4714 2663 4725 2666
rect 4714 2576 4717 2663
rect 4734 2576 4737 2763
rect 4746 2586 4749 3206
rect 4786 3203 4789 3806
rect 4754 3013 4757 3026
rect 4762 3023 4765 3036
rect 4770 3006 4773 3136
rect 4802 3096 4805 3186
rect 4762 3003 4773 3006
rect 4794 3093 4805 3096
rect 4754 2913 4757 2926
rect 4762 2906 4765 3003
rect 4794 2976 4797 3093
rect 4810 3076 4813 3096
rect 4806 3073 4813 3076
rect 4806 2996 4809 3073
rect 4806 2993 4813 2996
rect 4794 2973 4805 2976
rect 4758 2903 4765 2906
rect 4758 2836 4761 2903
rect 4754 2833 4761 2836
rect 4754 2773 4757 2833
rect 4754 2733 4757 2746
rect 4754 2613 4757 2726
rect 4762 2723 4765 2816
rect 4786 2776 4789 2946
rect 4802 2813 4805 2973
rect 4810 2796 4813 2993
rect 4806 2793 4813 2796
rect 4746 2583 4753 2586
rect 4778 2583 4781 2776
rect 4786 2773 4797 2776
rect 4794 2586 4797 2773
rect 4786 2583 4797 2586
rect 4714 2573 4721 2576
rect 4734 2573 4741 2576
rect 4706 2413 4709 2506
rect 4718 2486 4721 2573
rect 4718 2483 4725 2486
rect 4706 2393 4709 2406
rect 4714 2373 4717 2416
rect 4722 2383 4725 2483
rect 4730 2413 4733 2426
rect 4738 2413 4741 2573
rect 4750 2476 4753 2583
rect 4746 2473 4753 2476
rect 4730 2403 4741 2406
rect 4698 2313 4701 2326
rect 4706 2323 4717 2326
rect 4682 2293 4693 2296
rect 4674 2273 4681 2276
rect 4678 2166 4681 2273
rect 4674 2163 4681 2166
rect 4674 2103 4677 2163
rect 4690 2146 4693 2293
rect 4738 2276 4741 2396
rect 4730 2273 4741 2276
rect 4686 2143 4693 2146
rect 4686 2096 4689 2143
rect 4698 2113 4701 2126
rect 4706 2123 4709 2216
rect 4730 2176 4733 2273
rect 4730 2173 4741 2176
rect 4682 2093 4689 2096
rect 4666 2083 4673 2086
rect 4658 1923 4661 2006
rect 4670 1966 4673 2083
rect 4666 1963 4673 1966
rect 4646 1903 4653 1906
rect 4646 1846 4649 1903
rect 4642 1843 4649 1846
rect 4634 1633 4637 1776
rect 4642 1706 4645 1843
rect 4650 1813 4653 1826
rect 4658 1803 4661 1916
rect 4666 1803 4669 1963
rect 4674 1933 4677 1946
rect 4674 1903 4677 1926
rect 4674 1803 4677 1826
rect 4682 1786 4685 2093
rect 4690 1923 4693 2036
rect 4698 2003 4701 2016
rect 4678 1783 4685 1786
rect 4650 1713 4653 1726
rect 4642 1703 4649 1706
rect 4646 1636 4649 1703
rect 4646 1633 4653 1636
rect 4618 1453 4621 1606
rect 4626 1533 4629 1616
rect 4634 1583 4637 1606
rect 4578 1423 4589 1426
rect 4610 1423 4617 1426
rect 4570 1413 4581 1416
rect 4570 1373 4573 1406
rect 4554 933 4557 1196
rect 4546 903 4553 906
rect 4550 846 4553 903
rect 4562 893 4565 1216
rect 4578 1213 4581 1413
rect 4586 1383 4589 1423
rect 4594 1393 4597 1416
rect 4602 1333 4605 1406
rect 4614 1346 4617 1423
rect 4614 1343 4621 1346
rect 4570 1193 4573 1206
rect 4578 1186 4581 1206
rect 4578 1183 4585 1186
rect 4546 843 4553 846
rect 4546 773 4549 843
rect 4570 826 4573 1176
rect 4582 1036 4585 1183
rect 4578 1033 4585 1036
rect 4578 1003 4581 1033
rect 4586 1003 4589 1016
rect 4594 996 4597 1226
rect 4610 1213 4613 1326
rect 4610 1133 4613 1146
rect 4618 1036 4621 1343
rect 4626 1223 4629 1486
rect 4634 1396 4637 1576
rect 4642 1563 4645 1616
rect 4642 1533 4645 1556
rect 4650 1533 4653 1633
rect 4658 1603 4661 1736
rect 4666 1703 4669 1726
rect 4678 1716 4681 1783
rect 4690 1723 4693 1816
rect 4698 1813 4701 1826
rect 4714 1813 4717 2006
rect 4698 1776 4701 1806
rect 4714 1793 4717 1806
rect 4738 1783 4741 2173
rect 4746 1873 4749 2473
rect 4754 2433 4757 2456
rect 4754 2403 4757 2426
rect 4762 2413 4765 2526
rect 4754 2313 4757 2326
rect 4754 2123 4757 2206
rect 4754 2013 4757 2116
rect 4754 1923 4757 2006
rect 4762 1856 4765 2386
rect 4786 2133 4789 2583
rect 4806 2496 4809 2793
rect 4802 2493 4809 2496
rect 4802 2366 4805 2493
rect 4802 2363 4813 2366
rect 4810 2296 4813 2363
rect 4802 2293 4813 2296
rect 4802 2166 4805 2293
rect 4802 2163 4809 2166
rect 4786 2106 4789 2126
rect 4786 2103 4797 2106
rect 4794 2013 4797 2103
rect 4794 1923 4797 1946
rect 4758 1853 4765 1856
rect 4746 1813 4749 1826
rect 4758 1796 4761 1853
rect 4806 1836 4809 2163
rect 4758 1793 4765 1796
rect 4698 1773 4705 1776
rect 4762 1773 4765 1793
rect 4702 1716 4705 1773
rect 4678 1713 4685 1716
rect 4682 1646 4685 1713
rect 4674 1643 4685 1646
rect 4698 1713 4705 1716
rect 4714 1713 4717 1736
rect 4674 1576 4677 1643
rect 4674 1573 4685 1576
rect 4634 1393 4641 1396
rect 4638 1256 4641 1393
rect 4634 1253 4641 1256
rect 4650 1253 4653 1526
rect 4658 1523 4661 1546
rect 4666 1533 4669 1556
rect 4674 1533 4677 1546
rect 4674 1473 4677 1526
rect 4682 1496 4685 1573
rect 4690 1533 4693 1636
rect 4698 1593 4701 1713
rect 4738 1613 4741 1726
rect 4778 1656 4781 1816
rect 4794 1813 4797 1836
rect 4806 1833 4813 1836
rect 4810 1813 4813 1833
rect 4778 1653 4785 1656
rect 4714 1566 4717 1606
rect 4706 1563 4717 1566
rect 4706 1533 4709 1563
rect 4690 1513 4693 1526
rect 4730 1513 4733 1526
rect 4682 1493 4693 1496
rect 4626 1113 4629 1216
rect 4578 993 4597 996
rect 4578 906 4581 993
rect 4586 923 4589 936
rect 4578 903 4585 906
rect 4594 903 4597 926
rect 4582 836 4585 903
rect 4602 896 4605 1036
rect 4618 1033 4625 1036
rect 4634 1033 4637 1253
rect 4658 1203 4661 1356
rect 4674 1333 4677 1456
rect 4690 1396 4693 1493
rect 4746 1426 4749 1616
rect 4782 1586 4785 1653
rect 4794 1613 4797 1626
rect 4778 1583 4785 1586
rect 4778 1566 4781 1583
rect 4774 1563 4781 1566
rect 4774 1516 4777 1563
rect 4786 1523 4789 1556
rect 4774 1513 4781 1516
rect 4778 1456 4781 1513
rect 4778 1453 4785 1456
rect 4746 1423 4757 1426
rect 4682 1393 4693 1396
rect 4666 1313 4669 1326
rect 4674 1203 4677 1216
rect 4650 1143 4669 1146
rect 4610 1013 4613 1026
rect 4554 823 4573 826
rect 4578 833 4585 836
rect 4594 893 4605 896
rect 4554 756 4557 823
rect 4550 753 4557 756
rect 4550 656 4553 753
rect 4550 653 4557 656
rect 4514 643 4541 646
rect 4450 563 4461 566
rect 4490 573 4497 576
rect 4418 523 4421 536
rect 4426 533 4429 546
rect 4386 513 4397 516
rect 4410 513 4421 516
rect 4394 413 4397 513
rect 4418 446 4421 513
rect 4450 466 4453 563
rect 4450 463 4461 466
rect 4414 443 4421 446
rect 4370 343 4381 346
rect 4298 296 4301 316
rect 4298 293 4309 296
rect 4306 236 4309 293
rect 4298 233 4309 236
rect 4234 203 4245 206
rect 4290 203 4293 226
rect 4298 213 4301 233
rect 4210 133 4213 156
rect 4234 133 4237 203
rect 4282 113 4285 126
rect 4314 123 4317 196
rect 4322 133 4325 216
rect 4330 193 4333 336
rect 4338 213 4341 266
rect 4362 203 4365 336
rect 4378 276 4381 343
rect 4402 313 4405 436
rect 4414 366 4417 443
rect 4414 363 4421 366
rect 4410 323 4413 336
rect 4418 323 4421 363
rect 4426 333 4429 396
rect 4434 323 4437 376
rect 4442 333 4445 406
rect 4458 393 4461 463
rect 4466 413 4469 556
rect 4490 456 4493 573
rect 4482 453 4493 456
rect 4482 386 4485 453
rect 4506 413 4509 526
rect 4514 496 4517 643
rect 4554 633 4557 653
rect 4546 603 4549 626
rect 4514 493 4521 496
rect 4518 386 4521 493
rect 4530 413 4533 586
rect 4554 523 4557 616
rect 4562 533 4565 816
rect 4570 733 4573 816
rect 4578 803 4581 833
rect 4586 776 4589 816
rect 4594 803 4597 893
rect 4602 803 4605 816
rect 4610 793 4613 986
rect 4622 976 4625 1033
rect 4634 993 4637 1006
rect 4642 983 4645 1136
rect 4650 1123 4653 1143
rect 4658 1123 4661 1136
rect 4666 1133 4669 1143
rect 4650 1013 4653 1116
rect 4658 993 4661 1006
rect 4622 973 4645 976
rect 4618 943 4637 946
rect 4618 923 4621 943
rect 4626 923 4629 936
rect 4634 933 4637 943
rect 4578 773 4589 776
rect 4570 613 4573 646
rect 4570 506 4573 606
rect 4578 573 4581 773
rect 4594 733 4597 746
rect 4594 713 4597 726
rect 4602 666 4605 736
rect 4618 733 4621 916
rect 4634 906 4637 926
rect 4642 913 4645 973
rect 4666 926 4669 1126
rect 4674 1123 4677 1196
rect 4682 1026 4685 1393
rect 4690 1323 4693 1376
rect 4714 1353 4717 1406
rect 4714 1313 4717 1336
rect 4738 1323 4741 1416
rect 4754 1316 4757 1423
rect 4782 1376 4785 1453
rect 4794 1413 4797 1426
rect 4746 1313 4757 1316
rect 4778 1373 4785 1376
rect 4714 1236 4717 1256
rect 4710 1233 4717 1236
rect 4746 1236 4749 1313
rect 4746 1233 4753 1236
rect 4690 1213 4693 1226
rect 4690 1123 4693 1206
rect 4698 1193 4701 1216
rect 4682 1023 4689 1026
rect 4650 923 4669 926
rect 4626 903 4637 906
rect 4626 813 4629 903
rect 4626 793 4629 806
rect 4634 803 4637 816
rect 4642 786 4645 806
rect 4650 796 4653 816
rect 4658 803 4661 816
rect 4666 813 4669 836
rect 4666 796 4669 806
rect 4674 803 4677 1016
rect 4686 946 4689 1023
rect 4698 1003 4701 1126
rect 4710 1096 4713 1233
rect 4730 1203 4733 1216
rect 4738 1123 4741 1226
rect 4750 1116 4753 1233
rect 4746 1113 4753 1116
rect 4710 1093 4717 1096
rect 4714 1076 4717 1093
rect 4714 1073 4725 1076
rect 4722 996 4725 1073
rect 4746 1013 4749 1113
rect 4682 943 4689 946
rect 4714 993 4725 996
rect 4650 793 4669 796
rect 4642 783 4653 786
rect 4626 703 4629 726
rect 4602 663 4613 666
rect 4586 566 4589 636
rect 4602 613 4605 626
rect 4594 603 4605 606
rect 4562 503 4573 506
rect 4578 563 4589 566
rect 4562 456 4565 503
rect 4562 453 4573 456
rect 4570 433 4573 453
rect 4554 403 4557 416
rect 4482 383 4493 386
rect 4490 363 4493 383
rect 4482 343 4501 346
rect 4434 296 4437 316
rect 4370 273 4381 276
rect 4430 293 4437 296
rect 4370 253 4373 273
rect 4430 236 4433 293
rect 4430 233 4437 236
rect 4410 213 4413 226
rect 4434 216 4437 233
rect 4442 223 4445 326
rect 4450 266 4453 336
rect 4482 333 4485 343
rect 4466 303 4469 326
rect 4490 323 4493 336
rect 4498 323 4501 343
rect 4506 333 4509 386
rect 4514 383 4521 386
rect 4514 363 4517 383
rect 4450 263 4461 266
rect 4434 213 4445 216
rect 4450 213 4453 236
rect 4458 166 4461 263
rect 4450 163 4461 166
rect 4370 133 4373 156
rect 4322 113 4325 126
rect 4418 113 4421 126
rect 4450 123 4453 163
rect 4466 133 4469 216
rect 4474 203 4477 216
rect 4482 213 4485 246
rect 4514 243 4517 326
rect 4522 306 4525 336
rect 4530 323 4533 376
rect 4570 373 4573 416
rect 4522 303 4529 306
rect 4526 246 4529 303
rect 4538 296 4541 356
rect 4546 333 4549 366
rect 4554 323 4557 356
rect 4570 323 4573 336
rect 4578 313 4581 563
rect 4610 523 4613 663
rect 4618 613 4621 656
rect 4626 603 4629 616
rect 4538 293 4549 296
rect 4522 243 4529 246
rect 4498 213 4501 236
rect 4522 226 4525 243
rect 4546 236 4549 293
rect 4514 223 4525 226
rect 4538 233 4549 236
rect 4458 113 4461 126
rect 4498 123 4501 206
rect 4514 203 4517 223
rect 4522 196 4525 216
rect 4530 203 4533 216
rect 4538 213 4541 233
rect 4538 196 4541 206
rect 4522 193 4541 196
rect 4554 123 4557 216
rect 4578 213 4581 236
rect 4586 153 4589 406
rect 4610 403 4613 516
rect 4618 503 4621 526
rect 4634 513 4637 756
rect 4650 736 4653 783
rect 4682 753 4685 943
rect 4690 913 4693 926
rect 4698 923 4709 926
rect 4714 886 4717 993
rect 4730 913 4733 926
rect 4778 896 4781 1373
rect 4778 893 4789 896
rect 4714 883 4725 886
rect 4690 746 4693 836
rect 4698 813 4701 826
rect 4706 813 4717 816
rect 4642 703 4645 736
rect 4650 733 4661 736
rect 4674 733 4677 746
rect 4682 743 4693 746
rect 4650 693 4653 726
rect 4642 613 4645 686
rect 4658 626 4661 733
rect 4666 713 4669 726
rect 4650 623 4661 626
rect 4650 533 4653 623
rect 4658 596 4661 616
rect 4666 603 4669 706
rect 4674 596 4677 606
rect 4658 593 4677 596
rect 4658 543 4677 546
rect 4658 523 4661 543
rect 4594 333 4597 386
rect 4618 353 4621 416
rect 4666 413 4669 536
rect 4674 533 4677 543
rect 4682 523 4685 743
rect 4690 713 4693 736
rect 4698 723 4701 736
rect 4706 723 4709 746
rect 4714 706 4717 806
rect 4710 703 4717 706
rect 4690 613 4693 626
rect 4698 613 4701 636
rect 4710 576 4713 703
rect 4722 683 4725 883
rect 4738 813 4741 826
rect 4738 723 4741 736
rect 4786 636 4789 893
rect 4778 633 4789 636
rect 4730 613 4733 626
rect 4710 573 4717 576
rect 4674 496 4677 516
rect 4714 513 4717 573
rect 4674 493 4693 496
rect 4690 406 4693 493
rect 4746 413 4749 526
rect 4618 343 4637 346
rect 4610 293 4613 336
rect 4618 323 4621 343
rect 4626 323 4629 336
rect 4634 333 4637 343
rect 4610 176 4613 216
rect 4618 203 4621 216
rect 4626 203 4629 216
rect 4634 213 4637 326
rect 4642 203 4645 406
rect 4674 403 4693 406
rect 4778 403 4781 633
rect 4650 196 4653 216
rect 4658 203 4661 296
rect 4666 196 4669 206
rect 4674 203 4677 403
rect 4690 313 4693 326
rect 4706 246 4709 346
rect 4730 313 4733 326
rect 4778 323 4789 326
rect 4706 243 4717 246
rect 4698 213 4701 226
rect 4714 203 4717 243
rect 4738 213 4741 226
rect 4794 213 4797 236
rect 4650 193 4669 196
rect 4594 173 4613 176
rect 4578 133 4581 146
rect 4594 133 4597 173
rect 4618 133 4621 146
rect 4602 113 4605 126
rect 4642 113 4645 126
rect 4698 123 4701 156
rect 4817 37 4837 4703
rect 4841 13 4861 4727
rect 4866 2823 4877 2826
rect 4866 1663 4869 2816
rect 4874 606 4877 2823
rect 4866 603 4877 606
rect 4866 593 4869 603
<< metal3 >>
rect 2001 4682 2318 4687
rect 937 4652 1086 4657
rect 497 4642 686 4647
rect 497 4637 502 4642
rect 473 4632 502 4637
rect 681 4637 686 4642
rect 937 4637 942 4652
rect 1081 4637 1086 4652
rect 2233 4652 2310 4657
rect 2233 4647 2238 4652
rect 1129 4642 1206 4647
rect 1937 4642 2238 4647
rect 2305 4647 2310 4652
rect 2369 4652 2446 4657
rect 2369 4647 2374 4652
rect 2305 4642 2374 4647
rect 2441 4647 2446 4652
rect 2441 4642 2494 4647
rect 1129 4637 1134 4642
rect 681 4632 942 4637
rect 977 4632 1062 4637
rect 1081 4632 1134 4637
rect 1201 4637 1206 4642
rect 1201 4632 1310 4637
rect 3649 4632 3686 4637
rect 4193 4632 4310 4637
rect 977 4627 982 4632
rect 545 4622 590 4627
rect 953 4622 982 4627
rect 1057 4627 1062 4632
rect 1057 4622 1190 4627
rect 1777 4622 1822 4627
rect 1945 4622 1990 4627
rect 2249 4622 2294 4627
rect 2385 4622 2430 4627
rect 2657 4622 2702 4627
rect 2801 4622 2846 4627
rect 3761 4622 3790 4627
rect 3929 4622 3958 4627
rect 4193 4622 4238 4627
rect 4561 4622 4646 4627
rect 4753 4617 4758 4627
rect 505 4612 670 4617
rect 689 4612 902 4617
rect 937 4612 1118 4617
rect 3233 4612 3390 4617
rect 4753 4612 4877 4617
rect 689 4607 694 4612
rect 249 4602 294 4607
rect 401 4602 438 4607
rect 489 4602 534 4607
rect 649 4602 694 4607
rect 897 4607 902 4612
rect 1137 4607 1246 4612
rect 897 4602 1142 4607
rect 1241 4602 1270 4607
rect 1313 4602 1390 4607
rect 1745 4602 1798 4607
rect 2121 4602 2406 4607
rect 2545 4602 2590 4607
rect 2121 4597 2126 4602
rect 161 4592 246 4597
rect 313 4592 358 4597
rect 593 4592 782 4597
rect 825 4592 918 4597
rect 1001 4592 1102 4597
rect 1113 4592 1222 4597
rect 1433 4592 1566 4597
rect 1649 4592 1734 4597
rect 241 4587 246 4592
rect 417 4587 486 4592
rect 1729 4587 1734 4592
rect 1809 4592 1910 4597
rect 1953 4592 1990 4597
rect 2097 4592 2126 4597
rect 2401 4597 2406 4602
rect 3233 4597 3238 4612
rect 2401 4592 2430 4597
rect 2449 4592 2662 4597
rect 2825 4592 3046 4597
rect 3177 4592 3238 4597
rect 3385 4597 3390 4612
rect 3577 4602 3694 4607
rect 3713 4602 3806 4607
rect 4209 4602 4366 4607
rect 3713 4597 3718 4602
rect 3385 4592 3582 4597
rect 1809 4587 1814 4592
rect 241 4582 422 4587
rect 481 4582 510 4587
rect 657 4582 694 4587
rect 873 4582 1142 4587
rect 1473 4582 1510 4587
rect 1729 4582 1814 4587
rect 1905 4587 1910 4592
rect 2449 4587 2454 4592
rect 3577 4587 3582 4592
rect 3649 4592 3718 4597
rect 3801 4597 3806 4602
rect 3801 4592 3934 4597
rect 3649 4587 3654 4592
rect 1905 4582 2454 4587
rect 3249 4582 3374 4587
rect 3577 4582 3654 4587
rect 3673 4582 3830 4587
rect 529 4577 638 4582
rect 3825 4577 3830 4582
rect 4049 4582 4190 4587
rect 4049 4577 4054 4582
rect 0 4572 70 4577
rect 433 4572 534 4577
rect 633 4572 678 4577
rect 777 4572 958 4577
rect 1073 4572 1150 4577
rect 1257 4572 1414 4577
rect 1969 4572 2102 4577
rect 2681 4572 2878 4577
rect 3097 4572 3222 4577
rect 3825 4572 4054 4577
rect 4185 4577 4190 4582
rect 4385 4582 4486 4587
rect 4385 4577 4390 4582
rect 4185 4572 4390 4577
rect 4481 4577 4486 4582
rect 4481 4572 4782 4577
rect 329 4567 438 4572
rect 1257 4567 1262 4572
rect 185 4562 334 4567
rect 457 4562 686 4567
rect 897 4562 1094 4567
rect 1121 4562 1262 4567
rect 1409 4567 1414 4572
rect 2681 4567 2686 4572
rect 1409 4562 1622 4567
rect 1841 4562 2006 4567
rect 721 4557 814 4562
rect 1841 4557 1846 4562
rect 2001 4557 2006 4562
rect 2081 4562 2278 4567
rect 2609 4562 2686 4567
rect 2873 4567 2878 4572
rect 2873 4562 3086 4567
rect 3233 4562 3406 4567
rect 3521 4562 3662 4567
rect 2081 4557 2086 4562
rect 3081 4557 3238 4562
rect 3657 4557 3662 4562
rect 3809 4562 3926 4567
rect 3961 4562 4110 4567
rect 3809 4557 3814 4562
rect 4129 4557 4262 4562
rect 297 4552 566 4557
rect 601 4552 726 4557
rect 809 4552 838 4557
rect 905 4552 942 4557
rect 1057 4552 1134 4557
rect 1289 4552 1334 4557
rect 1345 4552 1438 4557
rect 1753 4552 1846 4557
rect 1945 4552 1982 4557
rect 2001 4552 2086 4557
rect 2233 4552 2414 4557
rect 2729 4552 2862 4557
rect 2945 4552 2974 4557
rect 3377 4552 3574 4557
rect 3657 4552 3814 4557
rect 3833 4552 3894 4557
rect 3929 4552 4134 4557
rect 4257 4552 4470 4557
rect 3377 4547 3382 4552
rect 129 4542 190 4547
rect 273 4542 518 4547
rect 529 4542 622 4547
rect 513 4537 518 4542
rect 641 4537 646 4547
rect 737 4542 782 4547
rect 913 4542 1070 4547
rect 1089 4542 1182 4547
rect 1273 4542 1374 4547
rect 1393 4542 1438 4547
rect 1513 4542 1590 4547
rect 1793 4542 1838 4547
rect 1921 4542 1974 4547
rect 2241 4542 2262 4547
rect 2449 4542 2590 4547
rect 2633 4542 2766 4547
rect 2857 4542 3382 4547
rect 3401 4542 3582 4547
rect 4017 4542 4046 4547
rect 2449 4537 2454 4542
rect 345 4532 486 4537
rect 513 4532 646 4537
rect 849 4532 886 4537
rect 897 4532 926 4537
rect 1017 4532 1046 4537
rect 1193 4532 1390 4537
rect 2425 4532 2454 4537
rect 2585 4537 2590 4542
rect 4041 4537 4046 4542
rect 4137 4542 4166 4547
rect 4193 4542 4270 4547
rect 4137 4537 4142 4542
rect 2585 4532 2830 4537
rect 3529 4532 3574 4537
rect 4041 4532 4142 4537
rect 4401 4532 4510 4537
rect 1041 4527 1198 4532
rect 321 4522 454 4527
rect 817 4522 990 4527
rect 1257 4522 1502 4527
rect 1817 4522 1966 4527
rect 2129 4522 2222 4527
rect 2545 4522 2590 4527
rect 2617 4522 2718 4527
rect 2849 4522 2958 4527
rect 3121 4522 3286 4527
rect 3313 4522 3502 4527
rect 4297 4522 4390 4527
rect 4401 4517 4406 4532
rect 4505 4527 4510 4532
rect 4505 4522 4614 4527
rect 4753 4522 4877 4527
rect 305 4512 406 4517
rect 465 4512 574 4517
rect 593 4512 702 4517
rect 721 4512 766 4517
rect 881 4512 926 4517
rect 977 4512 1102 4517
rect 1193 4512 1230 4517
rect 1345 4512 1374 4517
rect 1393 4512 1422 4517
rect 1433 4512 1510 4517
rect 1521 4512 1654 4517
rect 1665 4512 1814 4517
rect 1825 4512 1982 4517
rect 2009 4512 2038 4517
rect 2145 4512 2174 4517
rect 2441 4512 2678 4517
rect 2825 4512 2878 4517
rect 3057 4512 3102 4517
rect 3265 4512 3326 4517
rect 3337 4512 3446 4517
rect 3545 4512 3598 4517
rect 4097 4512 4142 4517
rect 4161 4512 4206 4517
rect 4265 4512 4406 4517
rect 4441 4512 4494 4517
rect 4753 4512 4758 4522
rect 401 4507 470 4512
rect 593 4507 598 4512
rect 153 4502 382 4507
rect 545 4502 598 4507
rect 697 4507 702 4512
rect 697 4502 910 4507
rect 1049 4502 1326 4507
rect 1489 4502 1534 4507
rect 1745 4502 1774 4507
rect 281 4492 310 4497
rect 305 4487 310 4492
rect 401 4492 478 4497
rect 553 4492 750 4497
rect 1209 4492 1238 4497
rect 401 4487 406 4492
rect 1233 4487 1238 4492
rect 1441 4492 1470 4497
rect 1441 4487 1446 4492
rect 305 4482 406 4487
rect 537 4482 734 4487
rect 1233 4482 1446 4487
rect 1769 4487 1774 4502
rect 1913 4502 1942 4507
rect 1969 4502 2086 4507
rect 2537 4502 2662 4507
rect 3001 4502 3158 4507
rect 3201 4502 3270 4507
rect 4097 4502 4150 4507
rect 4169 4502 4398 4507
rect 1913 4487 1918 4502
rect 2033 4492 2070 4497
rect 2521 4492 2630 4497
rect 2961 4492 3606 4497
rect 3625 4492 3766 4497
rect 4193 4492 4222 4497
rect 1769 4482 1918 4487
rect 2681 4482 2942 4487
rect 3081 4482 3254 4487
rect 3625 4482 3630 4492
rect 2681 4477 2686 4482
rect 2937 4477 3062 4482
rect 3489 4477 3630 4482
rect 3761 4477 3766 4492
rect 4217 4487 4222 4492
rect 4409 4492 4702 4497
rect 4409 4487 4414 4492
rect 4217 4482 4414 4487
rect 425 4472 654 4477
rect 801 4472 934 4477
rect 953 4472 1142 4477
rect 2657 4472 2686 4477
rect 3057 4472 3494 4477
rect 3649 4472 3734 4477
rect 3761 4472 3790 4477
rect 3809 4472 4038 4477
rect 801 4467 806 4472
rect 481 4462 510 4467
rect 665 4462 806 4467
rect 929 4467 934 4472
rect 3649 4467 3654 4472
rect 929 4462 998 4467
rect 505 4457 670 4462
rect 993 4457 998 4462
rect 1153 4462 1214 4467
rect 1937 4462 2030 4467
rect 1153 4457 1158 4462
rect 1937 4457 1942 4462
rect 849 4452 894 4457
rect 993 4452 1158 4457
rect 1857 4452 1942 4457
rect 2025 4457 2030 4462
rect 2209 4462 2278 4467
rect 2209 4457 2214 4462
rect 2025 4452 2214 4457
rect 2273 4457 2278 4462
rect 2385 4462 2606 4467
rect 2625 4462 3654 4467
rect 3729 4467 3734 4472
rect 3729 4462 3758 4467
rect 2385 4457 2390 4462
rect 2273 4452 2390 4457
rect 2601 4457 2606 4462
rect 3809 4457 3814 4472
rect 2601 4452 2734 4457
rect 2873 4452 3814 4457
rect 4033 4457 4038 4472
rect 4161 4462 4246 4467
rect 4161 4457 4166 4462
rect 4033 4452 4062 4457
rect 4137 4452 4166 4457
rect 4241 4457 4246 4462
rect 4289 4462 4438 4467
rect 4241 4452 4270 4457
rect 2729 4447 2878 4452
rect 4289 4447 4294 4462
rect 553 4442 750 4447
rect 817 4442 974 4447
rect 1721 4442 1782 4447
rect 2425 4442 2518 4447
rect 2561 4442 2614 4447
rect 2681 4442 2710 4447
rect 2425 4437 2430 4442
rect 545 4432 590 4437
rect 625 4432 926 4437
rect 985 4432 1150 4437
rect 1689 4432 1782 4437
rect 1793 4432 1910 4437
rect 1945 4432 2014 4437
rect 2225 4432 2262 4437
rect 2401 4432 2430 4437
rect 2513 4437 2518 4442
rect 2705 4437 2710 4442
rect 2897 4442 2966 4447
rect 3073 4442 3126 4447
rect 3441 4442 3678 4447
rect 3809 4442 4030 4447
rect 4257 4442 4294 4447
rect 4433 4447 4438 4462
rect 4561 4452 4606 4457
rect 4433 4442 4550 4447
rect 2897 4437 2902 4442
rect 3217 4437 3318 4442
rect 3673 4437 3814 4442
rect 2513 4432 2542 4437
rect 2705 4432 2902 4437
rect 2921 4432 2966 4437
rect 3113 4432 3222 4437
rect 3313 4432 3366 4437
rect 3545 4432 3654 4437
rect 4129 4432 4198 4437
rect 4233 4432 4598 4437
rect 4609 4432 4646 4437
rect 1793 4427 1798 4432
rect 4609 4427 4614 4432
rect 241 4422 342 4427
rect 465 4412 526 4417
rect 561 4402 566 4427
rect 585 4422 726 4427
rect 769 4422 998 4427
rect 1057 4422 1094 4427
rect 1241 4422 1326 4427
rect 1425 4422 1590 4427
rect 1657 4422 1702 4427
rect 1761 4422 1798 4427
rect 1825 4422 1966 4427
rect 2193 4422 2238 4427
rect 2385 4422 2454 4427
rect 2473 4422 2518 4427
rect 2953 4422 2998 4427
rect 3233 4422 3334 4427
rect 3385 4422 3430 4427
rect 3585 4422 3630 4427
rect 3729 4422 3774 4427
rect 3793 4422 3862 4427
rect 4033 4422 4182 4427
rect 4401 4422 4502 4427
rect 3041 4417 3190 4422
rect 3793 4417 3798 4422
rect 689 4412 718 4417
rect 881 4412 910 4417
rect 1225 4412 1486 4417
rect 1889 4412 2022 4417
rect 2041 4412 2134 4417
rect 713 4407 886 4412
rect 1025 4407 1110 4412
rect 2041 4407 2046 4412
rect 937 4402 1030 4407
rect 1105 4402 1134 4407
rect 1809 4402 1886 4407
rect 1881 4397 1886 4402
rect 1985 4402 2046 4407
rect 2129 4407 2134 4412
rect 2665 4412 2846 4417
rect 2665 4407 2670 4412
rect 2129 4402 2198 4407
rect 1985 4397 1990 4402
rect 2193 4397 2198 4402
rect 2257 4402 2350 4407
rect 2369 4402 2406 4407
rect 2641 4402 2670 4407
rect 2841 4407 2846 4412
rect 3017 4412 3046 4417
rect 3185 4412 3214 4417
rect 3265 4412 3310 4417
rect 3369 4412 3478 4417
rect 3497 4412 3798 4417
rect 3857 4417 3862 4422
rect 4497 4417 4502 4422
rect 4561 4422 4614 4427
rect 4633 4422 4678 4427
rect 4561 4417 4566 4422
rect 3857 4412 4166 4417
rect 3017 4407 3022 4412
rect 2841 4402 3022 4407
rect 3209 4407 3214 4412
rect 4161 4407 4166 4412
rect 4225 4412 4254 4417
rect 4337 4412 4422 4417
rect 4433 4412 4478 4417
rect 4497 4412 4566 4417
rect 4657 4412 4877 4417
rect 4225 4407 4230 4412
rect 4433 4407 4438 4412
rect 3209 4402 3302 4407
rect 3329 4402 3726 4407
rect 3769 4402 4142 4407
rect 4161 4402 4230 4407
rect 4329 4402 4438 4407
rect 2257 4397 2262 4402
rect 193 4392 318 4397
rect 361 4392 470 4397
rect 497 4392 718 4397
rect 737 4392 766 4397
rect 833 4392 862 4397
rect 857 4387 862 4392
rect 1041 4392 1070 4397
rect 1089 4392 1166 4397
rect 1217 4392 1270 4397
rect 1433 4392 1510 4397
rect 1609 4392 1654 4397
rect 1793 4392 1846 4397
rect 1881 4392 1990 4397
rect 2009 4392 2110 4397
rect 2193 4392 2262 4397
rect 2345 4397 2350 4402
rect 2689 4397 2822 4402
rect 2345 4392 2694 4397
rect 2817 4392 3286 4397
rect 1041 4387 1046 4392
rect 3281 4387 3286 4392
rect 3449 4392 3566 4397
rect 3769 4392 3862 4397
rect 4017 4392 4046 4397
rect 4441 4392 4566 4397
rect 3449 4387 3454 4392
rect 3561 4387 3774 4392
rect 3857 4387 4022 4392
rect 393 4382 486 4387
rect 553 4382 798 4387
rect 857 4382 1046 4387
rect 2145 4382 2182 4387
rect 2177 4377 2182 4382
rect 2257 4382 2286 4387
rect 2297 4382 2430 4387
rect 2593 4382 2774 4387
rect 2785 4382 3006 4387
rect 3161 4382 3262 4387
rect 3281 4382 3454 4387
rect 3513 4382 3542 4387
rect 3793 4382 3838 4387
rect 2257 4377 2262 4382
rect 3001 4377 3166 4382
rect 0 4372 174 4377
rect 185 4372 382 4377
rect 377 4367 382 4372
rect 449 4372 542 4377
rect 625 4372 750 4377
rect 2089 4372 2158 4377
rect 2177 4372 2262 4377
rect 2449 4372 2574 4377
rect 2753 4372 2854 4377
rect 3473 4372 3782 4377
rect 3849 4372 4126 4377
rect 4673 4372 4726 4377
rect 449 4367 454 4372
rect 537 4367 630 4372
rect 2449 4367 2454 4372
rect 377 4362 454 4367
rect 961 4362 1006 4367
rect 1177 4362 1422 4367
rect 1937 4362 2142 4367
rect 2329 4362 2398 4367
rect 2409 4362 2454 4367
rect 2569 4367 2574 4372
rect 2633 4367 2702 4372
rect 2873 4367 2982 4372
rect 3185 4367 3334 4372
rect 3777 4367 3854 4372
rect 2569 4362 2638 4367
rect 2697 4362 2790 4367
rect 2801 4362 2878 4367
rect 2977 4362 3190 4367
rect 3329 4362 3574 4367
rect 3873 4362 3902 4367
rect 3977 4362 4118 4367
rect 649 4357 726 4362
rect 3569 4357 3574 4362
rect 169 4352 230 4357
rect 473 4352 526 4357
rect 625 4352 654 4357
rect 721 4352 798 4357
rect 969 4352 1006 4357
rect 1281 4352 1398 4357
rect 2105 4352 2558 4357
rect 2649 4352 2686 4357
rect 2761 4352 2966 4357
rect 3201 4352 3318 4357
rect 3497 4352 3526 4357
rect 3569 4352 3638 4357
rect 3665 4352 3894 4357
rect 4081 4352 4238 4357
rect 4297 4352 4374 4357
rect 4393 4352 4454 4357
rect 1137 4347 1286 4352
rect 3201 4347 3206 4352
rect 3337 4347 3454 4352
rect 4297 4347 4302 4352
rect 129 4342 190 4347
rect 281 4342 374 4347
rect 473 4342 542 4347
rect 681 4342 710 4347
rect 841 4342 886 4347
rect 897 4342 974 4347
rect 1009 4342 1142 4347
rect 1297 4342 1502 4347
rect 1673 4342 1806 4347
rect 2433 4342 2598 4347
rect 2673 4342 2718 4347
rect 2817 4342 2950 4347
rect 3041 4342 3206 4347
rect 3305 4342 3342 4347
rect 3449 4342 3726 4347
rect 897 4337 902 4342
rect 3041 4337 3046 4342
rect 3721 4337 3726 4342
rect 3809 4342 4206 4347
rect 4273 4342 4302 4347
rect 4369 4347 4374 4352
rect 4369 4342 4462 4347
rect 3809 4337 3814 4342
rect 113 4332 142 4337
rect 201 4332 270 4337
rect 137 4327 206 4332
rect 265 4327 270 4332
rect 329 4332 694 4337
rect 833 4332 902 4337
rect 1153 4332 1638 4337
rect 2481 4332 2534 4337
rect 2609 4332 2662 4337
rect 2753 4332 3046 4337
rect 3065 4332 3094 4337
rect 3209 4332 3246 4337
rect 3257 4332 3670 4337
rect 3721 4332 3814 4337
rect 4041 4332 4142 4337
rect 4409 4332 4446 4337
rect 329 4327 334 4332
rect 937 4327 1014 4332
rect 4289 4327 4358 4332
rect 265 4322 334 4327
rect 369 4322 654 4327
rect 777 4322 942 4327
rect 1009 4322 1038 4327
rect 1281 4322 1454 4327
rect 2705 4322 2774 4327
rect 2913 4322 3006 4327
rect 3129 4322 3358 4327
rect 3457 4322 3494 4327
rect 3881 4322 3926 4327
rect 2913 4317 2918 4322
rect 3001 4317 3134 4322
rect 3921 4317 3926 4322
rect 4033 4322 4294 4327
rect 4353 4322 4710 4327
rect 4033 4317 4038 4322
rect 129 4312 182 4317
rect 353 4312 494 4317
rect 609 4312 638 4317
rect 809 4312 854 4317
rect 953 4312 1270 4317
rect 1497 4312 1526 4317
rect 1697 4312 1742 4317
rect 1913 4312 1958 4317
rect 1969 4312 2358 4317
rect 2545 4312 2654 4317
rect 2673 4312 2718 4317
rect 2737 4312 2918 4317
rect 2937 4312 2982 4317
rect 3321 4312 3366 4317
rect 3545 4312 3590 4317
rect 3601 4312 3702 4317
rect 3857 4312 3902 4317
rect 3921 4312 4038 4317
rect 4057 4312 4182 4317
rect 4305 4312 4342 4317
rect 4441 4312 4486 4317
rect 4577 4312 4630 4317
rect 1265 4307 1382 4312
rect 1497 4307 1502 4312
rect 2545 4307 2550 4312
rect 193 4302 766 4307
rect 889 4302 942 4307
rect 761 4297 766 4302
rect 937 4297 942 4302
rect 1065 4302 1094 4307
rect 1377 4302 1502 4307
rect 1841 4302 1902 4307
rect 1065 4297 1070 4302
rect 1897 4297 1902 4302
rect 1969 4302 1998 4307
rect 2393 4302 2502 4307
rect 2521 4302 2550 4307
rect 2649 4307 2654 4312
rect 2649 4302 2710 4307
rect 2913 4302 3126 4307
rect 1969 4297 1974 4302
rect 2393 4297 2398 4302
rect 393 4292 422 4297
rect 417 4277 422 4292
rect 561 4292 590 4297
rect 761 4292 870 4297
rect 937 4292 1070 4297
rect 1225 4292 1294 4297
rect 1897 4292 1974 4297
rect 2361 4292 2398 4297
rect 2497 4297 2502 4302
rect 3121 4297 3126 4302
rect 3273 4302 3478 4307
rect 3521 4302 3614 4307
rect 4097 4302 4214 4307
rect 4321 4302 4374 4307
rect 3273 4297 3278 4302
rect 2497 4292 2870 4297
rect 3121 4292 3278 4297
rect 3313 4292 3414 4297
rect 561 4277 566 4292
rect 585 4282 622 4287
rect 417 4272 566 4277
rect 865 4277 870 4292
rect 1225 4287 1230 4292
rect 3409 4287 3414 4292
rect 3529 4292 3622 4297
rect 3529 4287 3534 4292
rect 1105 4282 1230 4287
rect 1249 4282 1358 4287
rect 2409 4282 2566 4287
rect 2601 4282 2734 4287
rect 3409 4282 3534 4287
rect 3929 4282 4078 4287
rect 1105 4277 1110 4282
rect 865 4272 1110 4277
rect 1889 4272 2094 4277
rect 1889 4267 1894 4272
rect 1865 4262 1894 4267
rect 2089 4267 2094 4272
rect 2185 4272 2342 4277
rect 2561 4272 2846 4277
rect 2985 4272 3102 4277
rect 3297 4272 3390 4277
rect 3553 4272 3694 4277
rect 2185 4267 2190 4272
rect 2089 4262 2190 4267
rect 2337 4267 2342 4272
rect 2337 4262 2678 4267
rect 2689 4262 2918 4267
rect 3177 4262 3294 4267
rect 3409 4262 3510 4267
rect 3409 4257 3414 4262
rect 209 4252 350 4257
rect 761 4252 790 4257
rect 1937 4252 2078 4257
rect 2185 4252 2262 4257
rect 2609 4252 2750 4257
rect 2841 4252 2894 4257
rect 3129 4252 3174 4257
rect 3241 4252 3414 4257
rect 3505 4257 3510 4262
rect 3553 4257 3558 4272
rect 3505 4252 3558 4257
rect 3689 4257 3694 4272
rect 3929 4267 3934 4282
rect 4073 4277 4078 4282
rect 4073 4272 4270 4277
rect 3905 4262 3934 4267
rect 4265 4267 4270 4272
rect 4265 4262 4326 4267
rect 3689 4252 4254 4257
rect 4321 4252 4454 4257
rect 209 4247 214 4252
rect 185 4242 214 4247
rect 345 4247 350 4252
rect 4249 4247 4326 4252
rect 345 4242 374 4247
rect 601 4242 742 4247
rect 961 4242 1078 4247
rect 1745 4242 1798 4247
rect 1833 4242 1934 4247
rect 2193 4242 3278 4247
rect 2057 4237 2158 4242
rect 3273 4237 3278 4242
rect 3425 4242 3590 4247
rect 3697 4242 3846 4247
rect 3425 4237 3430 4242
rect 3585 4237 3702 4242
rect 329 4232 382 4237
rect 401 4232 478 4237
rect 625 4232 678 4237
rect 785 4232 806 4237
rect 1785 4232 2022 4237
rect 2033 4232 2062 4237
rect 2153 4232 2182 4237
rect 2649 4232 2758 4237
rect 2825 4232 2910 4237
rect 3073 4232 3254 4237
rect 3273 4232 3430 4237
rect 3521 4232 3566 4237
rect 3721 4232 3766 4237
rect 3881 4232 4094 4237
rect 4273 4232 4318 4237
rect 4329 4232 4366 4237
rect 193 4227 310 4232
rect 401 4227 406 4232
rect 169 4222 198 4227
rect 305 4222 406 4227
rect 473 4227 478 4232
rect 473 4222 678 4227
rect 729 4222 862 4227
rect 889 4222 982 4227
rect 993 4222 1094 4227
rect 1361 4222 1470 4227
rect 1649 4222 1694 4227
rect 1705 4222 1814 4227
rect 1921 4222 1982 4227
rect 1977 4217 1982 4222
rect 2057 4222 2150 4227
rect 2169 4222 2206 4227
rect 2345 4222 2406 4227
rect 2521 4222 2702 4227
rect 2809 4222 2854 4227
rect 2953 4222 3030 4227
rect 3049 4222 3094 4227
rect 3153 4222 3198 4227
rect 3633 4222 3678 4227
rect 3889 4222 3918 4227
rect 2057 4217 2062 4222
rect 0 4212 70 4217
rect 233 4212 462 4217
rect 593 4212 806 4217
rect 865 4212 926 4217
rect 1025 4212 1118 4217
rect 1225 4212 1302 4217
rect 1713 4212 1750 4217
rect 1769 4212 1894 4217
rect 1937 4212 1958 4217
rect 1977 4212 2062 4217
rect 2145 4217 2150 4222
rect 2145 4212 2470 4217
rect 2497 4212 2526 4217
rect 2625 4212 3214 4217
rect 3353 4212 3630 4217
rect 3745 4212 3878 4217
rect 1745 4207 1750 4212
rect 361 4202 422 4207
rect 633 4202 694 4207
rect 817 4202 846 4207
rect 969 4202 1358 4207
rect 1745 4202 1766 4207
rect 1793 4202 1870 4207
rect 417 4197 422 4202
rect 841 4197 950 4202
rect 161 4192 190 4197
rect 201 4192 238 4197
rect 281 4192 374 4197
rect 417 4192 622 4197
rect 657 4192 758 4197
rect 945 4192 1086 4197
rect 1177 4192 1254 4197
rect 1289 4192 1406 4197
rect 1601 4192 1702 4197
rect 1713 4192 1886 4197
rect 1937 4192 1942 4212
rect 2521 4207 2630 4212
rect 3913 4207 3918 4222
rect 4081 4222 4198 4227
rect 4417 4222 4694 4227
rect 4081 4207 4086 4222
rect 4297 4212 4358 4217
rect 4489 4212 4542 4217
rect 4745 4212 4877 4217
rect 2145 4202 2182 4207
rect 2649 4202 3062 4207
rect 3913 4202 4086 4207
rect 2321 4197 2454 4202
rect 3081 4197 3254 4202
rect 3321 4197 3750 4202
rect 2209 4192 2326 4197
rect 2449 4192 2678 4197
rect 2761 4192 3086 4197
rect 3249 4192 3278 4197
rect 3297 4192 3326 4197
rect 3745 4192 3774 4197
rect 4201 4192 4374 4197
rect 4545 4192 4582 4197
rect 377 4182 462 4187
rect 777 4182 886 4187
rect 881 4177 886 4182
rect 969 4182 1046 4187
rect 1057 4182 1390 4187
rect 1681 4182 1782 4187
rect 1929 4182 2014 4187
rect 2337 4182 2438 4187
rect 2945 4182 3894 4187
rect 4209 4182 4246 4187
rect 4561 4182 4630 4187
rect 969 4177 974 4182
rect 2465 4177 2806 4182
rect 2849 4177 2950 4182
rect 705 4172 862 4177
rect 881 4172 974 4177
rect 1729 4172 1790 4177
rect 2017 4172 2086 4177
rect 2449 4172 2470 4177
rect 2801 4172 2854 4177
rect 2961 4172 2990 4177
rect 3209 4172 3710 4177
rect 1225 4167 1350 4172
rect 2337 4167 2454 4172
rect 2985 4167 3214 4172
rect 561 4162 606 4167
rect 785 4162 822 4167
rect 1113 4162 1182 4167
rect 1201 4162 1230 4167
rect 1345 4162 1446 4167
rect 2241 4162 2342 4167
rect 2473 4162 2790 4167
rect 2865 4162 2942 4167
rect 3329 4162 3534 4167
rect 3729 4162 3886 4167
rect 4025 4162 4310 4167
rect 1113 4157 1118 4162
rect 553 4152 862 4157
rect 993 4152 1118 4157
rect 1177 4157 1182 4162
rect 1785 4157 1870 4162
rect 3233 4157 3310 4162
rect 3553 4157 3734 4162
rect 3881 4157 3886 4162
rect 1177 4152 1302 4157
rect 1321 4152 1350 4157
rect 1585 4152 1790 4157
rect 1865 4152 2062 4157
rect 2297 4152 2462 4157
rect 2529 4152 2910 4157
rect 2457 4147 2534 4152
rect 2905 4147 2910 4152
rect 3017 4152 3238 4157
rect 3305 4152 3558 4157
rect 3881 4152 3910 4157
rect 4169 4152 4206 4157
rect 4417 4152 4638 4157
rect 3017 4147 3022 4152
rect 129 4142 222 4147
rect 313 4142 414 4147
rect 537 4142 654 4147
rect 833 4142 854 4147
rect 905 4142 926 4147
rect 969 4142 1014 4147
rect 1129 4142 1190 4147
rect 1329 4142 1398 4147
rect 1473 4142 1518 4147
rect 1801 4142 1854 4147
rect 2169 4142 2254 4147
rect 2385 4142 2406 4147
rect 2553 4142 2638 4147
rect 2737 4142 2886 4147
rect 2905 4142 3022 4147
rect 3041 4142 3078 4147
rect 3249 4142 3478 4147
rect 3529 4142 3598 4147
rect 3657 4142 3870 4147
rect 3905 4142 4046 4147
rect 4169 4142 4198 4147
rect 4321 4142 4350 4147
rect 4409 4142 4446 4147
rect 4601 4142 4790 4147
rect 2401 4137 2406 4142
rect 0 4132 182 4137
rect 209 4132 302 4137
rect 297 4127 302 4132
rect 377 4132 718 4137
rect 769 4132 806 4137
rect 985 4132 1110 4137
rect 1209 4132 1310 4137
rect 1337 4132 1502 4137
rect 2153 4132 2198 4137
rect 2257 4132 2302 4137
rect 2401 4132 2566 4137
rect 377 4127 382 4132
rect 1209 4127 1214 4132
rect 297 4122 382 4127
rect 569 4122 646 4127
rect 705 4122 742 4127
rect 777 4122 982 4127
rect 1145 4122 1214 4127
rect 1305 4127 1310 4132
rect 2561 4127 2566 4132
rect 2649 4132 2726 4137
rect 2649 4127 2654 4132
rect 1305 4122 1350 4127
rect 1585 4122 1862 4127
rect 2017 4122 2038 4127
rect 2561 4122 2654 4127
rect 2721 4127 2726 4132
rect 2817 4132 2846 4137
rect 3137 4132 3270 4137
rect 3337 4132 3366 4137
rect 3513 4132 3542 4137
rect 4057 4132 4390 4137
rect 2817 4127 2822 4132
rect 2721 4122 2822 4127
rect 3049 4122 3094 4127
rect 3209 4122 3286 4127
rect 2129 4117 2246 4122
rect 3281 4117 3286 4122
rect 401 4112 582 4117
rect 697 4112 734 4117
rect 1113 4112 1286 4117
rect 1321 4112 1366 4117
rect 1361 4107 1366 4112
rect 1513 4112 1566 4117
rect 1841 4112 1910 4117
rect 2057 4112 2134 4117
rect 2241 4112 2542 4117
rect 2977 4112 3014 4117
rect 3225 4112 3270 4117
rect 3281 4112 3342 4117
rect 1513 4107 1518 4112
rect 3361 4107 3366 4132
rect 3537 4127 4062 4132
rect 4473 4122 4606 4127
rect 4753 4122 4877 4127
rect 3401 4112 3446 4117
rect 3481 4112 3526 4117
rect 3569 4112 3606 4117
rect 3713 4112 4022 4117
rect 4177 4112 4222 4117
rect 4353 4112 4390 4117
rect 4689 4112 4734 4117
rect 3713 4107 3718 4112
rect 225 4102 390 4107
rect 385 4097 390 4102
rect 449 4102 534 4107
rect 545 4102 654 4107
rect 889 4102 1046 4107
rect 1137 4102 1190 4107
rect 1361 4102 1518 4107
rect 1817 4102 1894 4107
rect 2145 4102 2206 4107
rect 2561 4102 2894 4107
rect 2913 4102 3038 4107
rect 3145 4102 3318 4107
rect 3345 4102 3366 4107
rect 3433 4102 3494 4107
rect 3641 4102 3718 4107
rect 4017 4107 4022 4112
rect 4017 4102 4166 4107
rect 4233 4102 4422 4107
rect 449 4097 454 4102
rect 385 4092 454 4097
rect 529 4097 534 4102
rect 2233 4097 2302 4102
rect 2561 4097 2566 4102
rect 529 4092 558 4097
rect 665 4092 878 4097
rect 1057 4092 1342 4097
rect 1905 4092 2134 4097
rect 2217 4092 2238 4097
rect 2297 4092 2566 4097
rect 2889 4097 2894 4102
rect 4161 4097 4238 4102
rect 2889 4092 4006 4097
rect 553 4087 670 4092
rect 873 4087 974 4092
rect 1057 4087 1062 4092
rect 2129 4087 2222 4092
rect 2585 4087 2870 4092
rect 4001 4087 4006 4092
rect 4329 4092 4358 4097
rect 4377 4092 4630 4097
rect 4329 4087 4334 4092
rect 969 4082 1062 4087
rect 1097 4082 1126 4087
rect 625 4072 654 4077
rect 649 4067 654 4072
rect 721 4072 950 4077
rect 721 4067 726 4072
rect 649 4062 726 4067
rect 1121 4067 1126 4082
rect 1281 4082 1310 4087
rect 2249 4082 2286 4087
rect 2545 4082 2590 4087
rect 2865 4082 3238 4087
rect 3297 4082 3518 4087
rect 3633 4082 3678 4087
rect 4001 4082 4334 4087
rect 1281 4067 1286 4082
rect 2449 4077 2526 4082
rect 1657 4072 2454 4077
rect 2521 4072 3118 4077
rect 3241 4072 3982 4077
rect 1121 4062 1286 4067
rect 2273 4062 2302 4067
rect 2465 4062 3374 4067
rect 4001 4062 4118 4067
rect 4137 4062 4182 4067
rect 4201 4062 4350 4067
rect 2113 4057 2254 4062
rect 2321 4057 2446 4062
rect 3473 4057 4006 4062
rect 4113 4057 4118 4062
rect 4201 4057 4206 4062
rect 249 4052 398 4057
rect 249 4037 254 4052
rect 225 4032 254 4037
rect 393 4037 398 4052
rect 969 4052 1078 4057
rect 1889 4052 2118 4057
rect 2249 4052 2326 4057
rect 2441 4052 3478 4057
rect 4113 4052 4206 4057
rect 4345 4057 4350 4062
rect 4393 4062 4478 4067
rect 4393 4057 4398 4062
rect 4345 4052 4398 4057
rect 4473 4057 4478 4062
rect 4473 4052 4534 4057
rect 969 4047 974 4052
rect 745 4042 974 4047
rect 1073 4047 1078 4052
rect 1073 4042 1102 4047
rect 1993 4042 2022 4047
rect 2017 4037 2022 4042
rect 2129 4042 2342 4047
rect 2129 4037 2134 4042
rect 393 4032 422 4037
rect 1017 4032 1062 4037
rect 1297 4032 1398 4037
rect 2017 4032 2134 4037
rect 2337 4037 2342 4042
rect 2417 4042 2790 4047
rect 2417 4037 2422 4042
rect 2337 4032 2422 4037
rect 2593 4032 2670 4037
rect 1297 4027 1302 4032
rect 209 4022 574 4027
rect 617 4022 662 4027
rect 801 4022 966 4027
rect 1025 4022 1302 4027
rect 1393 4027 1398 4032
rect 2177 4027 2270 4032
rect 2665 4027 2670 4032
rect 2737 4032 2766 4037
rect 2737 4027 2742 4032
rect 1393 4022 1558 4027
rect 1617 4022 1662 4027
rect 2153 4022 2182 4027
rect 2265 4022 2294 4027
rect 2441 4022 2518 4027
rect 2529 4022 2646 4027
rect 2665 4022 2742 4027
rect 2785 4027 2790 4042
rect 2961 4042 3110 4047
rect 3169 4042 3342 4047
rect 3489 4042 3958 4047
rect 4145 4042 4222 4047
rect 4353 4042 4462 4047
rect 2961 4027 2966 4042
rect 3105 4037 3110 4042
rect 3337 4037 3494 4042
rect 3977 4037 4054 4042
rect 3105 4032 3182 4037
rect 3193 4032 3254 4037
rect 3273 4032 3318 4037
rect 3513 4032 3982 4037
rect 4049 4032 4342 4037
rect 4417 4032 4446 4037
rect 4337 4027 4422 4032
rect 2785 4022 2966 4027
rect 2985 4022 3046 4027
rect 3097 4022 4038 4027
rect 4121 4022 4166 4027
rect 4449 4022 4510 4027
rect 4561 4022 4606 4027
rect 4033 4017 4126 4022
rect 553 4012 790 4017
rect 785 4007 790 4012
rect 905 4012 934 4017
rect 961 4012 1102 4017
rect 1609 4012 1742 4017
rect 2169 4012 2342 4017
rect 2569 4012 2646 4017
rect 3017 4012 3134 4017
rect 3201 4012 3342 4017
rect 3505 4012 3558 4017
rect 4145 4012 4326 4017
rect 4585 4012 4742 4017
rect 905 4007 910 4012
rect 2377 4007 2478 4012
rect 3553 4007 4014 4012
rect 345 4002 374 4007
rect 441 4002 470 4007
rect 641 4002 710 4007
rect 785 4002 910 4007
rect 985 4002 1126 4007
rect 1313 4002 1422 4007
rect 1617 4002 1646 4007
rect 1641 3997 1646 4002
rect 1753 4002 1798 4007
rect 2353 4002 2382 4007
rect 2473 4002 2542 4007
rect 2817 4002 2846 4007
rect 3137 4002 3190 4007
rect 3321 4002 3366 4007
rect 3449 4002 3534 4007
rect 4009 4002 4174 4007
rect 4281 4002 4430 4007
rect 4497 4002 4526 4007
rect 1753 3997 1758 4002
rect 2241 3997 2334 4002
rect 2969 3997 3118 4002
rect 3209 3997 3302 4002
rect 4169 3997 4286 4002
rect 129 3992 222 3997
rect 297 3992 414 3997
rect 537 3992 582 3997
rect 609 3992 654 3997
rect 937 3992 1030 3997
rect 1217 3992 1270 3997
rect 1409 3992 1494 3997
rect 1641 3992 1758 3997
rect 2217 3992 2246 3997
rect 2329 3992 2590 3997
rect 2633 3992 2734 3997
rect 2865 3992 2894 3997
rect 2945 3992 2974 3997
rect 3113 3992 3214 3997
rect 3297 3992 3486 3997
rect 3649 3992 3718 3997
rect 3777 3992 3854 3997
rect 3865 3992 3998 3997
rect 4121 3992 4150 3997
rect 4305 3992 4334 3997
rect 4393 3992 4478 3997
rect 609 3987 614 3992
rect 3993 3987 4126 3992
rect 249 3982 318 3987
rect 425 3982 614 3987
rect 633 3982 806 3987
rect 897 3982 934 3987
rect 1425 3982 1454 3987
rect 1873 3982 2582 3987
rect 313 3977 430 3982
rect 2577 3977 2582 3982
rect 2689 3982 3302 3987
rect 3593 3982 3654 3987
rect 3705 3982 3830 3987
rect 3841 3982 3886 3987
rect 2689 3977 2694 3982
rect 3321 3977 3454 3982
rect 3841 3977 3846 3982
rect 457 3972 510 3977
rect 817 3972 886 3977
rect 209 3967 286 3972
rect 505 3967 510 3972
rect 713 3967 822 3972
rect 881 3967 886 3972
rect 945 3972 1358 3977
rect 2273 3972 2398 3977
rect 2521 3972 2558 3977
rect 2577 3972 2694 3977
rect 2713 3972 2774 3977
rect 2881 3972 2910 3977
rect 945 3967 950 3972
rect 2905 3967 2910 3972
rect 3001 3972 3030 3977
rect 3105 3972 3326 3977
rect 3449 3972 3478 3977
rect 3521 3972 3582 3977
rect 3001 3967 3006 3972
rect 3521 3967 3526 3972
rect 0 3962 174 3967
rect 185 3962 214 3967
rect 281 3962 406 3967
rect 505 3962 718 3967
rect 881 3962 950 3967
rect 1137 3962 1230 3967
rect 1729 3962 1806 3967
rect 2185 3962 2310 3967
rect 2433 3962 2518 3967
rect 2905 3962 3006 3967
rect 3249 3962 3310 3967
rect 3353 3962 3526 3967
rect 3577 3967 3582 3972
rect 3801 3972 3846 3977
rect 3881 3977 3886 3982
rect 4273 3982 4382 3987
rect 4273 3977 4278 3982
rect 3881 3972 4278 3977
rect 4297 3972 4350 3977
rect 3801 3967 3806 3972
rect 3577 3962 3806 3967
rect 3825 3962 3862 3967
rect 1001 3957 1118 3962
rect 1729 3957 1734 3962
rect 169 3952 198 3957
rect 225 3952 270 3957
rect 353 3952 486 3957
rect 737 3952 806 3957
rect 977 3952 1006 3957
rect 1113 3952 1222 3957
rect 1705 3952 1734 3957
rect 1801 3957 1806 3962
rect 3145 3957 3230 3962
rect 1801 3952 1830 3957
rect 2097 3952 2382 3957
rect 2465 3952 2686 3957
rect 2769 3952 2854 3957
rect 3057 3952 3150 3957
rect 3225 3952 3254 3957
rect 225 3947 230 3952
rect 737 3947 742 3952
rect 81 3942 230 3947
rect 241 3942 302 3947
rect 385 3942 422 3947
rect 553 3942 742 3947
rect 801 3947 806 3952
rect 2769 3947 2774 3952
rect 801 3942 942 3947
rect 969 3942 1070 3947
rect 1081 3942 1350 3947
rect 1361 3942 1478 3947
rect 1697 3942 1750 3947
rect 1961 3942 2254 3947
rect 2265 3942 2350 3947
rect 2529 3942 2566 3947
rect 2681 3942 2718 3947
rect 2745 3942 2774 3947
rect 2849 3947 2854 3952
rect 3249 3947 3254 3952
rect 3385 3952 3430 3957
rect 3849 3952 3950 3957
rect 4641 3952 4742 3957
rect 3385 3947 3390 3952
rect 4641 3947 4646 3952
rect 2849 3942 2878 3947
rect 3161 3942 3198 3947
rect 3249 3942 3390 3947
rect 3409 3942 3542 3947
rect 3681 3942 3726 3947
rect 3817 3942 3846 3947
rect 4001 3942 4046 3947
rect 4153 3942 4198 3947
rect 4313 3942 4358 3947
rect 4617 3942 4646 3947
rect 4737 3947 4742 3952
rect 4737 3942 4782 3947
rect 1345 3937 1350 3942
rect 361 3932 390 3937
rect 753 3932 790 3937
rect 1033 3932 1134 3937
rect 1345 3932 1422 3937
rect 1489 3932 1582 3937
rect 1713 3932 2206 3937
rect 2393 3932 2422 3937
rect 2657 3932 2686 3937
rect 2785 3932 2838 3937
rect 2897 3932 2926 3937
rect 3129 3932 3214 3937
rect 3433 3932 3454 3937
rect 385 3927 390 3932
rect 1153 3927 1270 3932
rect 1417 3927 1494 3932
rect 2681 3927 2790 3932
rect 2833 3927 2902 3932
rect 369 3922 390 3927
rect 625 3922 790 3927
rect 913 3922 942 3927
rect 1049 3922 1158 3927
rect 1265 3922 1390 3927
rect 1753 3922 1966 3927
rect 2041 3922 2062 3927
rect 2305 3922 2358 3927
rect 2401 3922 2446 3927
rect 2513 3922 2550 3927
rect 2977 3922 3014 3927
rect 3049 3922 3230 3927
rect 3585 3922 3638 3927
rect 3681 3917 3686 3942
rect 3729 3932 3918 3937
rect 4209 3932 4270 3937
rect 4337 3932 4366 3937
rect 4481 3932 4542 3937
rect 3921 3922 4326 3927
rect 4337 3922 4342 3932
rect 4369 3922 4494 3927
rect 4529 3922 4702 3927
rect 4721 3922 4877 3927
rect 4321 3917 4326 3922
rect 4369 3917 4374 3922
rect 129 3912 222 3917
rect 361 3912 582 3917
rect 833 3912 902 3917
rect 969 3912 998 3917
rect 1041 3912 1462 3917
rect 897 3907 974 3912
rect 1457 3907 1462 3912
rect 1537 3912 1566 3917
rect 1673 3912 1734 3917
rect 1817 3912 1878 3917
rect 2033 3912 2062 3917
rect 2201 3912 2414 3917
rect 2521 3912 2550 3917
rect 2729 3912 2782 3917
rect 2849 3912 2886 3917
rect 2993 3912 3030 3917
rect 3169 3912 3214 3917
rect 3281 3912 3390 3917
rect 3449 3912 3494 3917
rect 3633 3912 3686 3917
rect 3705 3912 3734 3917
rect 3825 3912 3902 3917
rect 3985 3912 4014 3917
rect 4153 3912 4198 3917
rect 4321 3912 4374 3917
rect 4385 3912 4526 3917
rect 4721 3912 4726 3922
rect 1537 3907 1542 3912
rect 3825 3907 3830 3912
rect 177 3902 646 3907
rect 1001 3902 1150 3907
rect 1209 3902 1310 3907
rect 1345 3902 1438 3907
rect 1457 3902 1542 3907
rect 1633 3902 1694 3907
rect 2401 3902 2486 3907
rect 2297 3897 2406 3902
rect 2609 3897 2614 3907
rect 2785 3902 2814 3907
rect 2897 3902 3062 3907
rect 3113 3902 3294 3907
rect 3377 3902 3462 3907
rect 3513 3902 3614 3907
rect 3713 3902 3830 3907
rect 3897 3907 3902 3912
rect 4009 3907 4158 3912
rect 3897 3902 3950 3907
rect 4177 3902 4310 3907
rect 4473 3902 4502 3907
rect 4681 3902 4726 3907
rect 2809 3897 2902 3902
rect 3513 3897 3518 3902
rect 3609 3897 3694 3902
rect 4305 3897 4478 3902
rect 377 3892 590 3897
rect 657 3892 822 3897
rect 585 3887 662 3892
rect 817 3887 822 3892
rect 1145 3892 1326 3897
rect 1145 3887 1150 3892
rect 1321 3887 1326 3892
rect 1401 3892 1430 3897
rect 2209 3892 2302 3897
rect 2425 3892 2614 3897
rect 2649 3892 2758 3897
rect 3009 3892 3086 3897
rect 3177 3892 3222 3897
rect 3313 3892 3342 3897
rect 3489 3892 3518 3897
rect 3689 3892 3894 3897
rect 1401 3887 1406 3892
rect 2649 3887 2654 3892
rect 449 3882 566 3887
rect 817 3882 1150 3887
rect 1169 3882 1238 3887
rect 1321 3882 1406 3887
rect 1761 3882 2198 3887
rect 2193 3877 2198 3882
rect 2313 3882 2398 3887
rect 2625 3882 2654 3887
rect 2753 3887 2758 3892
rect 3337 3887 3494 3892
rect 3889 3887 3894 3892
rect 3961 3892 4246 3897
rect 4601 3892 4646 3897
rect 3961 3887 3966 3892
rect 2753 3882 2998 3887
rect 2313 3877 2318 3882
rect 2393 3877 2502 3882
rect 2625 3877 2630 3882
rect 2993 3877 2998 3882
rect 3097 3882 3318 3887
rect 3521 3882 3606 3887
rect 3617 3882 3870 3887
rect 3889 3882 3966 3887
rect 4161 3882 4190 3887
rect 4257 3882 4494 3887
rect 3097 3877 3102 3882
rect 3617 3877 3622 3882
rect 4185 3877 4262 3882
rect 321 3872 366 3877
rect 361 3867 366 3872
rect 433 3872 462 3877
rect 545 3872 678 3877
rect 2193 3872 2318 3877
rect 2337 3872 2374 3877
rect 2497 3872 2630 3877
rect 2665 3872 2742 3877
rect 2993 3872 3102 3877
rect 3153 3872 3190 3877
rect 3233 3872 3374 3877
rect 3481 3872 3622 3877
rect 3705 3872 3742 3877
rect 433 3867 438 3872
rect 3761 3867 3918 3872
rect 361 3862 438 3867
rect 2337 3862 2478 3867
rect 3329 3862 3766 3867
rect 3913 3862 4150 3867
rect 4145 3857 4150 3862
rect 4217 3862 4510 3867
rect 4217 3857 4222 3862
rect 521 3852 678 3857
rect 521 3847 526 3852
rect 489 3842 526 3847
rect 673 3847 678 3852
rect 969 3852 1118 3857
rect 2121 3852 2174 3857
rect 2297 3852 2366 3857
rect 2497 3852 2566 3857
rect 2577 3852 3318 3857
rect 3529 3852 3630 3857
rect 3729 3852 3814 3857
rect 3849 3852 3902 3857
rect 4145 3852 4222 3857
rect 969 3847 974 3852
rect 673 3842 782 3847
rect 841 3842 974 3847
rect 841 3837 846 3842
rect 169 3832 190 3837
rect 537 3832 662 3837
rect 817 3832 846 3837
rect 1113 3837 1118 3852
rect 2577 3847 2582 3852
rect 1913 3842 2358 3847
rect 2377 3842 2406 3847
rect 2401 3837 2406 3842
rect 2513 3842 2582 3847
rect 3313 3847 3318 3852
rect 3313 3842 3510 3847
rect 3617 3842 3654 3847
rect 4265 3842 4350 3847
rect 4377 3842 4406 3847
rect 2513 3837 2518 3842
rect 3505 3837 3598 3842
rect 4265 3837 4270 3842
rect 1113 3832 1142 3837
rect 1169 3832 1310 3837
rect 2161 3832 2230 3837
rect 2401 3832 2518 3837
rect 2569 3832 2630 3837
rect 3137 3832 3294 3837
rect 3593 3832 3686 3837
rect 3697 3832 3726 3837
rect 3801 3832 3846 3837
rect 4241 3832 4270 3837
rect 4345 3837 4350 3842
rect 4345 3832 4406 3837
rect 1169 3827 1174 3832
rect 225 3807 230 3827
rect 249 3822 382 3827
rect 457 3822 550 3827
rect 713 3822 774 3827
rect 985 3822 1070 3827
rect 1105 3822 1174 3827
rect 1305 3827 1310 3832
rect 1305 3822 1334 3827
rect 1417 3822 1566 3827
rect 2129 3822 2174 3827
rect 2537 3822 2582 3827
rect 2673 3822 2870 3827
rect 3241 3822 3598 3827
rect 3737 3822 4158 3827
rect 4185 3822 4214 3827
rect 4297 3822 4334 3827
rect 4481 3822 4518 3827
rect 817 3817 950 3822
rect 3593 3817 3742 3822
rect 4209 3817 4302 3822
rect 689 3812 734 3817
rect 761 3812 822 3817
rect 945 3812 974 3817
rect 1041 3812 1430 3817
rect 1769 3812 1982 3817
rect 2009 3812 2118 3817
rect 2185 3812 2246 3817
rect 2113 3807 2190 3812
rect 2705 3807 2710 3817
rect 3161 3812 3206 3817
rect 3457 3812 3510 3817
rect 3537 3812 3574 3817
rect 4321 3812 4470 3817
rect 4529 3812 4630 3817
rect 3249 3807 3358 3812
rect 3825 3807 3934 3812
rect 4465 3807 4534 3812
rect 137 3802 214 3807
rect 225 3802 326 3807
rect 321 3797 326 3802
rect 393 3802 558 3807
rect 833 3802 1118 3807
rect 1361 3802 1470 3807
rect 1561 3802 1670 3807
rect 2705 3802 2806 3807
rect 3017 3802 3254 3807
rect 3353 3802 3446 3807
rect 3585 3802 3830 3807
rect 3929 3802 3958 3807
rect 3977 3802 4054 3807
rect 4145 3802 4206 3807
rect 4665 3802 4702 3807
rect 393 3797 398 3802
rect 3441 3797 3590 3802
rect 3977 3797 3982 3802
rect 161 3792 190 3797
rect 185 3787 190 3792
rect 273 3792 302 3797
rect 321 3792 398 3797
rect 521 3792 574 3797
rect 705 3792 798 3797
rect 953 3792 1062 3797
rect 1177 3792 1246 3797
rect 1449 3792 1574 3797
rect 1729 3792 1774 3797
rect 1873 3792 1910 3797
rect 1961 3792 2118 3797
rect 273 3787 278 3792
rect 2113 3787 2118 3792
rect 2201 3792 2294 3797
rect 2497 3792 2534 3797
rect 2705 3792 2926 3797
rect 3121 3792 3166 3797
rect 3265 3792 3342 3797
rect 3721 3792 3750 3797
rect 3841 3792 3870 3797
rect 3889 3792 3982 3797
rect 4049 3797 4054 3802
rect 4049 3792 4110 3797
rect 4409 3792 4430 3797
rect 4505 3792 4534 3797
rect 2201 3787 2206 3792
rect 4529 3787 4534 3792
rect 4617 3792 4710 3797
rect 4617 3787 4622 3792
rect 185 3782 278 3787
rect 633 3782 926 3787
rect 1217 3782 1302 3787
rect 2113 3782 2206 3787
rect 2225 3782 2334 3787
rect 2401 3782 2422 3787
rect 3089 3782 3278 3787
rect 3417 3782 4118 3787
rect 4113 3777 4118 3782
rect 4217 3782 4294 3787
rect 4529 3782 4622 3787
rect 4217 3777 4222 3782
rect 649 3772 718 3777
rect 865 3772 1222 3777
rect 745 3767 870 3772
rect 1217 3767 1222 3772
rect 1313 3772 1406 3777
rect 1745 3772 1782 3777
rect 1881 3772 1918 3777
rect 2057 3772 2094 3777
rect 3073 3772 3150 3777
rect 3233 3772 3406 3777
rect 3889 3772 4006 3777
rect 4065 3772 4094 3777
rect 4113 3772 4222 3777
rect 1313 3767 1318 3772
rect 3145 3767 3238 3772
rect 3401 3767 3894 3772
rect 553 3762 750 3767
rect 889 3762 910 3767
rect 1217 3762 1318 3767
rect 1665 3762 1734 3767
rect 1729 3757 1734 3762
rect 1793 3762 1870 3767
rect 1793 3757 1798 3762
rect 193 3752 286 3757
rect 697 3752 910 3757
rect 1049 3752 1198 3757
rect 1193 3747 1198 3752
rect 1361 3752 1390 3757
rect 1729 3752 1798 3757
rect 1865 3757 1870 3762
rect 1929 3762 1958 3767
rect 3097 3762 3126 3767
rect 3257 3762 3302 3767
rect 3913 3762 3942 3767
rect 3953 3762 3982 3767
rect 4025 3762 4086 3767
rect 1929 3757 1934 3762
rect 1865 3752 1934 3757
rect 2625 3752 2718 3757
rect 2801 3752 2902 3757
rect 3249 3752 3662 3757
rect 3721 3752 3902 3757
rect 3929 3752 4078 3757
rect 4337 3752 4422 3757
rect 4681 3752 4750 3757
rect 1361 3747 1366 3752
rect 4337 3747 4342 3752
rect 233 3742 350 3747
rect 465 3742 550 3747
rect 609 3742 710 3747
rect 777 3742 806 3747
rect 953 3742 1070 3747
rect 1193 3742 1366 3747
rect 1577 3742 1606 3747
rect 2425 3742 2518 3747
rect 2769 3742 2822 3747
rect 3065 3742 3158 3747
rect 3201 3742 3326 3747
rect 3441 3742 3470 3747
rect 3569 3742 3598 3747
rect 3713 3742 3742 3747
rect 3737 3737 3742 3742
rect 3921 3742 3990 3747
rect 3921 3737 3926 3742
rect 201 3732 278 3737
rect 361 3732 654 3737
rect 673 3732 790 3737
rect 833 3732 942 3737
rect 273 3727 366 3732
rect 225 3722 254 3727
rect 393 3722 422 3727
rect 545 3722 798 3727
rect 881 3722 910 3727
rect 937 3717 942 3732
rect 1081 3732 1134 3737
rect 1489 3732 1630 3737
rect 2321 3732 2398 3737
rect 2945 3732 3038 3737
rect 3073 3732 3102 3737
rect 3385 3732 3414 3737
rect 3737 3732 3926 3737
rect 3985 3737 3990 3742
rect 4073 3742 4174 3747
rect 4249 3742 4342 3747
rect 4417 3747 4422 3752
rect 4417 3742 4446 3747
rect 4489 3742 4534 3747
rect 4681 3742 4702 3747
rect 4073 3737 4078 3742
rect 3985 3732 4078 3737
rect 4097 3732 4174 3737
rect 4353 3732 4390 3737
rect 4585 3732 4726 3737
rect 1081 3717 1086 3732
rect 3433 3727 3574 3732
rect 4721 3727 4726 3732
rect 1153 3722 1174 3727
rect 1617 3722 1646 3727
rect 1681 3722 1838 3727
rect 1849 3722 1910 3727
rect 2625 3722 2926 3727
rect 2625 3717 2630 3722
rect 321 3712 718 3717
rect 937 3712 1086 3717
rect 1121 3712 1166 3717
rect 1401 3712 1470 3717
rect 1633 3712 1662 3717
rect 1729 3712 1774 3717
rect 1825 3712 1886 3717
rect 2105 3712 2142 3717
rect 2313 3712 2334 3717
rect 2417 3712 2438 3717
rect 2497 3712 2582 3717
rect 2601 3712 2630 3717
rect 2921 3717 2926 3722
rect 3121 3722 3286 3727
rect 3305 3722 3438 3727
rect 3569 3722 3662 3727
rect 3945 3722 3966 3727
rect 4161 3722 4190 3727
rect 4217 3722 4254 3727
rect 4393 3722 4414 3727
rect 4521 3722 4710 3727
rect 4721 3722 4877 3727
rect 3121 3717 3126 3722
rect 2921 3712 2982 3717
rect 3001 3712 3030 3717
rect 3057 3712 3126 3717
rect 3281 3717 3286 3722
rect 3281 3712 3662 3717
rect 3841 3712 3902 3717
rect 4057 3712 4158 3717
rect 4249 3712 4278 3717
rect 4465 3712 4534 3717
rect 4585 3712 4718 3717
rect 2497 3707 2502 3712
rect 241 3702 694 3707
rect 1169 3702 1254 3707
rect 1273 3702 1414 3707
rect 1409 3697 1414 3702
rect 1481 3702 1622 3707
rect 1481 3697 1486 3702
rect 337 3692 366 3697
rect 361 3687 366 3692
rect 465 3692 582 3697
rect 465 3687 470 3692
rect 577 3687 582 3692
rect 729 3692 766 3697
rect 1409 3692 1486 3697
rect 729 3687 734 3692
rect 273 3682 326 3687
rect 361 3682 470 3687
rect 489 3682 550 3687
rect 577 3682 734 3687
rect 1617 3687 1622 3702
rect 1897 3702 2094 3707
rect 1897 3687 1902 3702
rect 2089 3697 2094 3702
rect 2153 3702 2406 3707
rect 2473 3702 2502 3707
rect 2577 3707 2582 3712
rect 2977 3707 2982 3712
rect 3145 3707 3262 3712
rect 2577 3702 2966 3707
rect 2977 3702 3150 3707
rect 3257 3702 3310 3707
rect 3425 3702 3454 3707
rect 2153 3697 2158 3702
rect 2401 3697 2478 3702
rect 3449 3697 3454 3702
rect 3529 3702 3558 3707
rect 3745 3702 4054 3707
rect 4545 3702 4574 3707
rect 3529 3697 3534 3702
rect 2089 3692 2158 3697
rect 3081 3692 3286 3697
rect 3449 3692 3534 3697
rect 3681 3692 3734 3697
rect 2537 3687 2702 3692
rect 3729 3687 3734 3692
rect 3817 3692 3870 3697
rect 3817 3687 3822 3692
rect 1617 3682 1902 3687
rect 2417 3682 2494 3687
rect 2513 3682 2542 3687
rect 2697 3682 2726 3687
rect 2817 3682 3182 3687
rect 3297 3682 3422 3687
rect 321 3667 326 3682
rect 489 3667 494 3682
rect 2417 3677 2422 3682
rect 1153 3672 1390 3677
rect 2137 3672 2422 3677
rect 2489 3677 2494 3682
rect 2817 3677 2822 3682
rect 3177 3677 3302 3682
rect 3417 3677 3422 3682
rect 3569 3682 3646 3687
rect 3729 3682 3822 3687
rect 3569 3677 3574 3682
rect 2489 3672 2822 3677
rect 3089 3672 3158 3677
rect 321 3662 494 3667
rect 785 3662 990 3667
rect 545 3652 694 3657
rect 257 3642 278 3647
rect 545 3637 550 3652
rect 201 3632 246 3637
rect 425 3632 494 3637
rect 521 3632 550 3637
rect 689 3637 694 3652
rect 785 3647 790 3662
rect 985 3657 990 3662
rect 1153 3657 1158 3672
rect 985 3652 1078 3657
rect 1129 3652 1158 3657
rect 1385 3657 1390 3672
rect 2889 3667 2990 3672
rect 3153 3667 3158 3672
rect 3353 3672 3398 3677
rect 3417 3672 3574 3677
rect 3865 3677 3870 3692
rect 4169 3692 4382 3697
rect 4169 3687 4174 3692
rect 4065 3682 4174 3687
rect 4329 3682 4686 3687
rect 4065 3677 4070 3682
rect 3865 3672 4070 3677
rect 3353 3667 3358 3672
rect 2433 3662 2614 3667
rect 2769 3662 2894 3667
rect 2985 3662 3134 3667
rect 3153 3662 3358 3667
rect 2609 3657 2774 3662
rect 1385 3652 1414 3657
rect 2097 3652 2190 3657
rect 713 3642 750 3647
rect 761 3642 790 3647
rect 1073 3647 1078 3652
rect 2185 3647 2190 3652
rect 2329 3652 2590 3657
rect 2329 3647 2334 3652
rect 2585 3647 2590 3652
rect 2793 3652 2822 3657
rect 2905 3652 2974 3657
rect 2793 3647 2798 3652
rect 1073 3642 1414 3647
rect 1801 3642 1902 3647
rect 2185 3642 2334 3647
rect 2377 3642 2430 3647
rect 1801 3637 1806 3642
rect 689 3632 742 3637
rect 785 3632 974 3637
rect 1737 3632 1806 3637
rect 1897 3637 1902 3642
rect 2425 3637 2430 3642
rect 2537 3642 2566 3647
rect 2585 3642 2798 3647
rect 2937 3642 3014 3647
rect 3129 3642 3238 3647
rect 3257 3642 3318 3647
rect 3961 3642 3982 3647
rect 4393 3642 4494 3647
rect 2537 3637 2542 3642
rect 3129 3637 3134 3642
rect 1897 3632 1998 3637
rect 2425 3632 2542 3637
rect 2969 3632 3134 3637
rect 3233 3637 3238 3642
rect 4393 3637 4398 3642
rect 3233 3632 3350 3637
rect 3881 3632 3926 3637
rect 4369 3632 4398 3637
rect 4489 3637 4494 3642
rect 4489 3632 4518 3637
rect 4673 3632 4694 3637
rect 425 3627 430 3632
rect 129 3622 270 3627
rect 377 3622 430 3627
rect 489 3627 494 3632
rect 489 3622 638 3627
rect 681 3622 774 3627
rect 857 3622 902 3627
rect 1025 3622 1062 3627
rect 1081 3622 1166 3627
rect 1257 3622 1326 3627
rect 1433 3622 1542 3627
rect 1817 3622 1886 3627
rect 2129 3622 2166 3627
rect 2353 3622 2406 3627
rect 2585 3622 2614 3627
rect 2697 3622 2726 3627
rect 2865 3622 2990 3627
rect 3145 3622 3286 3627
rect 3841 3622 3894 3627
rect 3905 3622 3950 3627
rect 4201 3622 4374 3627
rect 4433 3622 4598 3627
rect 4649 3622 4678 3627
rect 1081 3617 1086 3622
rect 617 3612 926 3617
rect 1001 3612 1086 3617
rect 1161 3617 1166 3622
rect 1433 3617 1438 3622
rect 1161 3612 1190 3617
rect 1225 3612 1270 3617
rect 1369 3612 1438 3617
rect 1537 3617 1542 3622
rect 1537 3612 1590 3617
rect 1609 3612 1638 3617
rect 1961 3612 1998 3617
rect 2161 3612 2222 3617
rect 2305 3612 2374 3617
rect 2457 3612 2494 3617
rect 2961 3612 3102 3617
rect 3233 3612 3398 3617
rect 4465 3612 4646 3617
rect 4689 3607 4694 3632
rect 313 3602 414 3607
rect 441 3602 486 3607
rect 545 3602 710 3607
rect 1073 3602 1150 3607
rect 1281 3602 1430 3607
rect 2289 3602 2358 3607
rect 2489 3602 2662 3607
rect 2761 3602 2942 3607
rect 2993 3602 3054 3607
rect 3129 3602 3206 3607
rect 3265 3602 3430 3607
rect 3617 3602 3678 3607
rect 3737 3602 3822 3607
rect 4649 3602 4694 3607
rect 313 3597 318 3602
rect 289 3592 318 3597
rect 409 3597 414 3602
rect 1281 3597 1286 3602
rect 409 3592 430 3597
rect 425 3587 430 3592
rect 513 3592 542 3597
rect 673 3592 822 3597
rect 833 3592 862 3597
rect 953 3592 1022 3597
rect 1033 3592 1286 3597
rect 1329 3592 1526 3597
rect 1633 3592 1654 3597
rect 1929 3592 2046 3597
rect 2337 3592 2422 3597
rect 2537 3592 2558 3597
rect 513 3587 518 3592
rect 2761 3587 2766 3602
rect 241 3582 398 3587
rect 425 3582 518 3587
rect 633 3582 686 3587
rect 961 3582 982 3587
rect 993 3582 1110 3587
rect 1241 3582 1358 3587
rect 1385 3582 1414 3587
rect 1841 3582 1878 3587
rect 2257 3582 2510 3587
rect 2505 3577 2510 3582
rect 2585 3582 2766 3587
rect 2937 3587 2942 3602
rect 3737 3597 3742 3602
rect 3113 3592 3190 3597
rect 3337 3592 3518 3597
rect 3713 3592 3742 3597
rect 3817 3597 3822 3602
rect 4417 3597 4502 3602
rect 3817 3592 3918 3597
rect 3969 3592 4046 3597
rect 4161 3592 4198 3597
rect 4393 3592 4422 3597
rect 4497 3592 4694 3597
rect 2937 3582 3094 3587
rect 3225 3582 3278 3587
rect 3329 3582 3366 3587
rect 3377 3582 3414 3587
rect 3537 3582 3638 3587
rect 3657 3582 3742 3587
rect 4057 3582 4486 3587
rect 4625 3582 4670 3587
rect 2585 3577 2590 3582
rect 3441 3577 3542 3582
rect 3633 3577 3638 3582
rect 345 3572 406 3577
rect 881 3572 1094 3577
rect 1153 3572 1238 3577
rect 1313 3572 1422 3577
rect 2249 3572 2374 3577
rect 2457 3572 2486 3577
rect 2505 3572 2590 3577
rect 2777 3572 2806 3577
rect 2369 3567 2462 3572
rect 2801 3567 2806 3572
rect 3017 3572 3046 3577
rect 3417 3572 3446 3577
rect 3633 3572 3822 3577
rect 3841 3572 4046 3577
rect 4153 3572 4182 3577
rect 4417 3572 4438 3577
rect 3017 3567 3022 3572
rect 4041 3567 4158 3572
rect 729 3562 862 3567
rect 1049 3562 1102 3567
rect 1761 3562 2022 3567
rect 2305 3562 2350 3567
rect 2801 3562 3022 3567
rect 3265 3562 3294 3567
rect 3385 3562 3654 3567
rect 3761 3562 3878 3567
rect 3945 3562 3966 3567
rect 4561 3562 4622 3567
rect 729 3557 734 3562
rect 857 3557 1030 3562
rect 3649 3557 3766 3562
rect 105 3552 214 3557
rect 705 3552 734 3557
rect 1025 3552 1262 3557
rect 1673 3552 1742 3557
rect 2017 3552 2054 3557
rect 2073 3552 2230 3557
rect 2377 3552 2414 3557
rect 3785 3552 3870 3557
rect 4113 3552 4238 3557
rect 4417 3552 4510 3557
rect 4521 3552 4710 3557
rect 105 3547 110 3552
rect 81 3542 110 3547
rect 209 3547 214 3552
rect 1673 3547 1678 3552
rect 209 3542 238 3547
rect 281 3542 390 3547
rect 465 3542 558 3547
rect 601 3542 814 3547
rect 865 3542 894 3547
rect 889 3537 894 3542
rect 953 3542 998 3547
rect 1009 3542 1110 3547
rect 1393 3542 1486 3547
rect 1529 3542 1574 3547
rect 1649 3542 1678 3547
rect 1737 3547 1742 3552
rect 2073 3547 2078 3552
rect 1737 3542 2078 3547
rect 2225 3547 2230 3552
rect 3473 3547 3630 3552
rect 2225 3542 2366 3547
rect 2425 3542 2790 3547
rect 2897 3542 2982 3547
rect 3185 3542 3382 3547
rect 3417 3542 3478 3547
rect 3625 3542 3654 3547
rect 3777 3542 3966 3547
rect 3985 3542 4094 3547
rect 4161 3542 4398 3547
rect 4473 3542 4534 3547
rect 4577 3542 4614 3547
rect 4641 3542 4678 3547
rect 953 3537 958 3542
rect 1105 3537 1110 3542
rect 1225 3537 1326 3542
rect 2361 3537 2430 3542
rect 3985 3537 3990 3542
rect 1 3532 70 3537
rect 137 3532 166 3537
rect 393 3532 478 3537
rect 593 3532 678 3537
rect 889 3532 958 3537
rect 1001 3532 1030 3537
rect 1105 3532 1230 3537
rect 1321 3532 1406 3537
rect 2113 3532 2142 3537
rect 3489 3532 3622 3537
rect 3969 3532 3990 3537
rect 4089 3537 4094 3542
rect 4089 3532 4150 3537
rect 4233 3532 4262 3537
rect 4497 3532 4662 3537
rect 4697 3532 4750 3537
rect 65 3527 142 3532
rect 1769 3527 1878 3532
rect 3785 3527 3974 3532
rect 4145 3527 4238 3532
rect 193 3522 334 3527
rect 601 3522 718 3527
rect 977 3522 1086 3527
rect 1225 3522 1310 3527
rect 1569 3522 1606 3527
rect 1657 3522 1774 3527
rect 1873 3522 2350 3527
rect 3081 3522 3150 3527
rect 3177 3522 3278 3527
rect 3273 3517 3278 3522
rect 3409 3522 3534 3527
rect 3409 3517 3414 3522
rect 3529 3517 3534 3522
rect 3633 3522 3670 3527
rect 3705 3522 3790 3527
rect 3985 3522 4118 3527
rect 4393 3522 4414 3527
rect 4425 3522 4622 3527
rect 4673 3522 4694 3527
rect 3633 3517 3638 3522
rect 3985 3517 3990 3522
rect 129 3512 182 3517
rect 377 3512 646 3517
rect 833 3512 966 3517
rect 961 3497 966 3512
rect 1097 3512 1190 3517
rect 1097 3497 1102 3512
rect 1185 3507 1190 3512
rect 1249 3512 1278 3517
rect 1617 3512 1678 3517
rect 1729 3512 2334 3517
rect 2497 3512 2630 3517
rect 2841 3512 2934 3517
rect 3201 3512 3254 3517
rect 3273 3512 3414 3517
rect 3433 3512 3510 3517
rect 3529 3512 3638 3517
rect 3801 3512 3870 3517
rect 3929 3512 3990 3517
rect 4185 3512 4302 3517
rect 4313 3512 4518 3517
rect 1249 3507 1254 3512
rect 1185 3502 1254 3507
rect 2817 3502 2838 3507
rect 2913 3502 3094 3507
rect 3761 3502 3830 3507
rect 4153 3502 4198 3507
rect 4377 3502 4398 3507
rect 217 3492 254 3497
rect 961 3492 1102 3497
rect 3097 3492 3142 3497
rect 3569 3492 3726 3497
rect 3745 3492 3774 3497
rect 3937 3492 4190 3497
rect 3569 3487 3574 3492
rect 473 3482 686 3487
rect 2433 3482 2462 3487
rect 2481 3482 2710 3487
rect 2729 3482 2782 3487
rect 3545 3482 3574 3487
rect 3721 3487 3726 3492
rect 3793 3487 3862 3492
rect 3721 3482 3798 3487
rect 3857 3482 3974 3487
rect 2105 3472 2174 3477
rect 2257 3472 2366 3477
rect 2385 3472 2422 3477
rect 2257 3467 2262 3472
rect 233 3462 366 3467
rect 1329 3462 1366 3467
rect 2009 3462 2086 3467
rect 2233 3462 2262 3467
rect 2361 3467 2366 3472
rect 2481 3467 2486 3482
rect 2705 3467 2710 3482
rect 3657 3472 3702 3477
rect 3793 3472 3846 3477
rect 3985 3472 4118 3477
rect 3697 3467 3798 3472
rect 3841 3467 3990 3472
rect 2361 3462 2486 3467
rect 2505 3462 2654 3467
rect 2705 3462 2774 3467
rect 3225 3462 3478 3467
rect 3561 3462 3678 3467
rect 233 3447 238 3462
rect 185 3442 238 3447
rect 361 3447 366 3462
rect 2009 3457 2014 3462
rect 1481 3452 1534 3457
rect 1865 3452 2014 3457
rect 2081 3457 2086 3462
rect 2505 3457 2510 3462
rect 2081 3452 2382 3457
rect 2473 3452 2510 3457
rect 2649 3457 2654 3462
rect 3673 3457 3678 3462
rect 4129 3462 4414 3467
rect 4129 3457 4134 3462
rect 2649 3452 2758 3457
rect 3145 3452 3318 3457
rect 3569 3452 3654 3457
rect 3673 3452 4134 3457
rect 2377 3447 2478 3452
rect 361 3442 390 3447
rect 409 3442 518 3447
rect 409 3437 414 3442
rect 249 3432 414 3437
rect 513 3437 518 3442
rect 889 3442 958 3447
rect 1393 3442 1414 3447
rect 1585 3442 1662 3447
rect 2041 3442 2078 3447
rect 2281 3442 2358 3447
rect 889 3437 894 3442
rect 513 3432 654 3437
rect 681 3432 894 3437
rect 953 3437 958 3442
rect 2073 3437 2286 3442
rect 2353 3437 2358 3442
rect 2497 3442 2638 3447
rect 2801 3442 2934 3447
rect 3513 3442 3566 3447
rect 4505 3442 4766 3447
rect 2497 3437 2502 3442
rect 2801 3437 2806 3442
rect 953 3432 1390 3437
rect 1777 3432 1846 3437
rect 2025 3432 2054 3437
rect 2305 3432 2334 3437
rect 2353 3432 2502 3437
rect 2521 3432 2622 3437
rect 2657 3432 2806 3437
rect 2929 3437 2934 3442
rect 3161 3437 3262 3442
rect 4505 3437 4510 3442
rect 2929 3432 2958 3437
rect 3073 3432 3118 3437
rect 3137 3432 3166 3437
rect 3257 3432 3350 3437
rect 3561 3432 3694 3437
rect 3705 3432 3798 3437
rect 4329 3432 4366 3437
rect 4481 3432 4510 3437
rect 4761 3437 4766 3442
rect 4761 3432 4790 3437
rect 2657 3427 2662 3432
rect 225 3422 454 3427
rect 617 3422 670 3427
rect 1169 3422 1222 3427
rect 1401 3422 1454 3427
rect 1777 3422 1854 3427
rect 1913 3422 2030 3427
rect 2081 3422 2150 3427
rect 2193 3422 2270 3427
rect 2289 3422 2318 3427
rect 2609 3422 2662 3427
rect 2817 3422 2974 3427
rect 2993 3422 3038 3427
rect 3201 3422 3246 3427
rect 3585 3422 3638 3427
rect 3953 3422 4038 3427
rect 4233 3422 4302 3427
rect 4321 3422 4390 3427
rect 4697 3422 4758 3427
rect 2193 3417 2198 3422
rect 129 3412 166 3417
rect 361 3412 502 3417
rect 905 3412 942 3417
rect 1817 3412 1846 3417
rect 1993 3412 2062 3417
rect 257 3407 342 3412
rect 1841 3407 1998 3412
rect 2057 3407 2062 3412
rect 2161 3412 2198 3417
rect 2265 3417 2270 3422
rect 2513 3417 2590 3422
rect 2265 3412 2518 3417
rect 2585 3412 3118 3417
rect 2161 3407 2166 3412
rect 3113 3407 3118 3412
rect 3361 3412 3430 3417
rect 3537 3412 3582 3417
rect 3785 3412 3998 3417
rect 4217 3412 4486 3417
rect 4505 3412 4654 3417
rect 3361 3407 3366 3412
rect 169 3402 262 3407
rect 337 3402 654 3407
rect 689 3402 878 3407
rect 897 3402 942 3407
rect 2017 3402 2038 3407
rect 2057 3402 2166 3407
rect 2209 3402 2326 3407
rect 2529 3402 2678 3407
rect 2873 3402 3014 3407
rect 3113 3402 3366 3407
rect 3969 3402 4046 3407
rect 4249 3402 4342 3407
rect 4401 3402 4454 3407
rect 689 3397 694 3402
rect 161 3392 198 3397
rect 273 3392 382 3397
rect 433 3392 478 3397
rect 625 3392 694 3397
rect 873 3397 878 3402
rect 2321 3397 2326 3402
rect 2673 3397 2878 3402
rect 873 3392 934 3397
rect 1193 3392 1262 3397
rect 1305 3392 1350 3397
rect 1569 3392 1670 3397
rect 1857 3392 1958 3397
rect 2193 3392 2310 3397
rect 2321 3392 2382 3397
rect 2617 3392 2654 3397
rect 2897 3392 2950 3397
rect 2945 3387 2950 3392
rect 3025 3392 3094 3397
rect 3537 3392 3686 3397
rect 3953 3392 3982 3397
rect 4185 3392 4262 3397
rect 4305 3392 4358 3397
rect 4673 3392 4702 3397
rect 3025 3387 3030 3392
rect 217 3382 254 3387
rect 417 3382 446 3387
rect 961 3382 1142 3387
rect 1425 3382 1486 3387
rect 1665 3382 1694 3387
rect 1705 3382 1846 3387
rect 633 3377 750 3382
rect 961 3377 966 3382
rect 209 3372 406 3377
rect 449 3372 638 3377
rect 745 3372 966 3377
rect 1137 3377 1142 3382
rect 1841 3377 1846 3382
rect 1969 3382 2102 3387
rect 2193 3382 2238 3387
rect 2249 3382 2398 3387
rect 2481 3382 2614 3387
rect 2641 3382 2910 3387
rect 2945 3382 3030 3387
rect 3969 3382 4014 3387
rect 4145 3382 4246 3387
rect 4337 3382 4422 3387
rect 4633 3382 4686 3387
rect 1969 3377 1974 3382
rect 1137 3372 1166 3377
rect 1313 3372 1550 3377
rect 1569 3372 1702 3377
rect 1841 3372 1974 3377
rect 2049 3372 2094 3377
rect 2377 3372 2406 3377
rect 2505 3372 2534 3377
rect 3561 3372 3694 3377
rect 3873 3372 4110 3377
rect 4489 3372 4518 3377
rect 1569 3367 1574 3372
rect 2225 3367 2294 3372
rect 2561 3367 2638 3372
rect 2769 3367 2862 3372
rect 3561 3367 3566 3372
rect 649 3362 734 3367
rect 1273 3362 1406 3367
rect 1401 3357 1406 3362
rect 1489 3362 1574 3367
rect 1601 3362 1630 3367
rect 2113 3362 2230 3367
rect 2289 3362 2566 3367
rect 2633 3362 2774 3367
rect 2857 3362 2886 3367
rect 2929 3362 3030 3367
rect 3449 3362 3566 3367
rect 3689 3367 3694 3372
rect 3689 3362 3814 3367
rect 4009 3362 4038 3367
rect 4121 3362 4222 3367
rect 4313 3362 4438 3367
rect 1489 3357 1494 3362
rect 1625 3357 1734 3362
rect 2113 3357 2118 3362
rect 2929 3357 2934 3362
rect 361 3352 454 3357
rect 633 3352 998 3357
rect 1057 3352 1086 3357
rect 1113 3352 1326 3357
rect 1401 3352 1494 3357
rect 1729 3352 2118 3357
rect 2241 3352 2302 3357
rect 2353 3352 2390 3357
rect 2577 3352 2622 3357
rect 2785 3352 2934 3357
rect 3025 3357 3030 3362
rect 3833 3357 3910 3362
rect 4033 3357 4126 3362
rect 3025 3352 3054 3357
rect 3257 3352 3294 3357
rect 3393 3352 3438 3357
rect 137 3342 262 3347
rect 353 3342 382 3347
rect 377 3337 382 3342
rect 465 3342 662 3347
rect 713 3342 742 3347
rect 841 3342 862 3347
rect 1033 3342 1142 3347
rect 1177 3342 1230 3347
rect 1289 3342 1382 3347
rect 1513 3342 1630 3347
rect 1641 3342 1710 3347
rect 2201 3342 2486 3347
rect 2497 3342 2590 3347
rect 2729 3342 2822 3347
rect 2889 3342 2918 3347
rect 465 3337 470 3342
rect 945 3337 1014 3342
rect 2913 3337 2918 3342
rect 2985 3342 3014 3347
rect 3257 3342 3390 3347
rect 2985 3337 2990 3342
rect 377 3332 470 3337
rect 569 3332 646 3337
rect 785 3332 950 3337
rect 1009 3332 1054 3337
rect 1209 3332 1246 3337
rect 665 3327 734 3332
rect 193 3322 310 3327
rect 561 3322 670 3327
rect 729 3322 774 3327
rect 961 3322 998 3327
rect 1041 3322 1222 3327
rect 769 3317 838 3322
rect 961 3317 966 3322
rect 1241 3317 1246 3332
rect 1377 3332 1478 3337
rect 1377 3317 1382 3332
rect 1489 3327 1494 3337
rect 2273 3332 2566 3337
rect 2625 3332 2814 3337
rect 2913 3332 2990 3337
rect 3433 3337 3438 3352
rect 3577 3352 3678 3357
rect 3809 3352 3838 3357
rect 3905 3352 3966 3357
rect 4217 3352 4526 3357
rect 3577 3337 3582 3352
rect 3633 3342 3670 3347
rect 3785 3342 3894 3347
rect 4081 3342 4318 3347
rect 4345 3342 4398 3347
rect 3433 3332 3582 3337
rect 3641 3332 3670 3337
rect 3881 3332 3966 3337
rect 4209 3332 4238 3337
rect 4337 3332 4366 3337
rect 3665 3327 3670 3332
rect 4233 3327 4342 3332
rect 1425 3322 1494 3327
rect 2145 3322 2214 3327
rect 2353 3322 2382 3327
rect 2377 3317 2382 3322
rect 2457 3322 2534 3327
rect 2633 3322 2662 3327
rect 2793 3322 2822 3327
rect 3049 3322 3118 3327
rect 3649 3322 3670 3327
rect 4417 3322 4518 3327
rect 4657 3322 4686 3327
rect 4705 3322 4710 3387
rect 2457 3317 2462 3322
rect 2529 3317 2638 3322
rect 249 3312 646 3317
rect 689 3312 718 3317
rect 833 3312 966 3317
rect 985 3312 1054 3317
rect 1241 3312 1382 3317
rect 1457 3312 1558 3317
rect 1609 3312 1638 3317
rect 1985 3312 2006 3317
rect 2073 3312 2310 3317
rect 2377 3312 2462 3317
rect 2481 3312 2510 3317
rect 2505 3307 2510 3312
rect 2673 3312 2774 3317
rect 2809 3312 2846 3317
rect 3265 3312 3326 3317
rect 3601 3312 3814 3317
rect 4129 3312 4198 3317
rect 2673 3307 2678 3312
rect 4193 3307 4198 3312
rect 4265 3312 4310 3317
rect 4369 3312 4430 3317
rect 4545 3312 4726 3317
rect 4265 3307 4270 3312
rect 265 3302 294 3307
rect 289 3297 294 3302
rect 401 3302 430 3307
rect 577 3302 814 3307
rect 1617 3302 1710 3307
rect 2505 3302 2678 3307
rect 2865 3302 3030 3307
rect 3297 3302 3430 3307
rect 4193 3302 4270 3307
rect 401 3297 406 3302
rect 2865 3297 2870 3302
rect 289 3292 406 3297
rect 593 3292 870 3297
rect 2353 3292 2462 3297
rect 2353 3287 2358 3292
rect 145 3282 206 3287
rect 673 3282 1134 3287
rect 1649 3282 2358 3287
rect 2457 3287 2462 3292
rect 2761 3292 2870 3297
rect 2761 3287 2766 3292
rect 2457 3282 2518 3287
rect 2537 3282 2718 3287
rect 2737 3282 2766 3287
rect 3025 3287 3030 3302
rect 4305 3297 4310 3312
rect 4417 3302 4446 3307
rect 4417 3297 4422 3302
rect 3217 3292 3286 3297
rect 3345 3292 3430 3297
rect 4305 3292 4422 3297
rect 3281 3287 3350 3292
rect 3025 3282 3070 3287
rect 3449 3282 3542 3287
rect 3641 3282 3662 3287
rect 4001 3282 4030 3287
rect 2537 3277 2542 3282
rect 2409 3272 2542 3277
rect 2713 3277 2718 3282
rect 3449 3277 3454 3282
rect 2713 3272 3014 3277
rect 3081 3272 3454 3277
rect 3537 3277 3542 3282
rect 3537 3272 3566 3277
rect 641 3267 846 3272
rect 2249 3267 2358 3272
rect 3009 3267 3086 3272
rect 89 3262 438 3267
rect 457 3262 598 3267
rect 617 3262 646 3267
rect 841 3262 870 3267
rect 1177 3262 1318 3267
rect 2081 3262 2254 3267
rect 2353 3262 2542 3267
rect 2609 3262 2694 3267
rect 457 3257 462 3262
rect 425 3252 462 3257
rect 593 3257 598 3262
rect 1177 3257 1182 3262
rect 593 3252 1182 3257
rect 1313 3257 1318 3262
rect 2609 3257 2614 3262
rect 1313 3252 1374 3257
rect 2017 3252 2062 3257
rect 2265 3252 2342 3257
rect 2585 3252 2614 3257
rect 2689 3257 2694 3262
rect 3185 3257 3606 3262
rect 2689 3252 3030 3257
rect 3161 3252 3190 3257
rect 3601 3252 3750 3257
rect 2361 3247 2446 3252
rect 153 3242 182 3247
rect 609 3242 862 3247
rect 1961 3242 1990 3247
rect 2073 3242 2142 3247
rect 1049 3237 1166 3242
rect 1985 3237 2078 3242
rect 2137 3237 2142 3242
rect 2257 3242 2366 3247
rect 2441 3242 2710 3247
rect 2257 3237 2262 3242
rect 2705 3237 2710 3242
rect 2825 3242 2854 3247
rect 3113 3242 3134 3247
rect 3185 3242 3590 3247
rect 2825 3237 2830 3242
rect 385 3232 1054 3237
rect 1161 3232 1302 3237
rect 1665 3232 1726 3237
rect 2137 3232 2262 3237
rect 2281 3232 2430 3237
rect 2705 3232 2830 3237
rect 2969 3232 3158 3237
rect 3209 3232 3350 3237
rect 3521 3232 3550 3237
rect 4505 3232 4534 3237
rect 4553 3232 4590 3237
rect 1665 3227 1670 3232
rect 3345 3227 3526 3232
rect 617 3222 726 3227
rect 849 3222 886 3227
rect 1065 3222 1150 3227
rect 1217 3222 1286 3227
rect 1385 3222 1542 3227
rect 1609 3222 1670 3227
rect 1689 3222 1782 3227
rect 1945 3222 2054 3227
rect 2393 3222 2414 3227
rect 2425 3222 2686 3227
rect 3009 3222 3078 3227
rect 3177 3222 3214 3227
rect 3281 3222 3326 3227
rect 3609 3222 3958 3227
rect 4025 3222 4054 3227
rect 4481 3222 4646 3227
rect 361 3217 454 3222
rect 3609 3217 3614 3222
rect 313 3212 366 3217
rect 449 3212 494 3217
rect 945 3212 1014 3217
rect 1785 3212 1830 3217
rect 2025 3212 2118 3217
rect 2385 3212 2502 3217
rect 3033 3212 3510 3217
rect 3529 3212 3614 3217
rect 609 3207 686 3212
rect 3529 3207 3534 3212
rect 3953 3207 3958 3222
rect 4465 3212 4502 3217
rect 4553 3207 4694 3212
rect 177 3202 214 3207
rect 361 3202 390 3207
rect 385 3197 390 3202
rect 449 3202 614 3207
rect 681 3202 710 3207
rect 729 3202 806 3207
rect 841 3202 1070 3207
rect 1705 3202 1758 3207
rect 2481 3202 2502 3207
rect 2521 3202 2670 3207
rect 2689 3202 2726 3207
rect 2745 3202 2838 3207
rect 3177 3202 3534 3207
rect 3721 3202 3862 3207
rect 3953 3202 3982 3207
rect 4529 3202 4558 3207
rect 4689 3202 4750 3207
rect 449 3197 454 3202
rect 729 3197 734 3202
rect 273 3192 326 3197
rect 385 3192 454 3197
rect 473 3192 526 3197
rect 625 3192 734 3197
rect 801 3197 806 3202
rect 2521 3197 2526 3202
rect 801 3192 830 3197
rect 905 3192 950 3197
rect 1041 3192 1174 3197
rect 1193 3192 1270 3197
rect 1377 3192 1470 3197
rect 1609 3192 1662 3197
rect 1681 3192 1830 3197
rect 1929 3192 2174 3197
rect 2193 3192 2230 3197
rect 2313 3192 2398 3197
rect 2457 3192 2526 3197
rect 2665 3197 2670 3202
rect 2745 3197 2750 3202
rect 2665 3192 2750 3197
rect 2833 3197 2838 3202
rect 3721 3197 3726 3202
rect 2833 3192 2934 3197
rect 2953 3192 2990 3197
rect 3201 3192 3726 3197
rect 3857 3197 3862 3202
rect 3857 3192 4190 3197
rect 4545 3192 4678 3197
rect 2313 3187 2318 3192
rect 737 3182 894 3187
rect 953 3182 982 3187
rect 1089 3182 1390 3187
rect 1545 3182 1798 3187
rect 2201 3182 2262 3187
rect 2289 3182 2318 3187
rect 2393 3187 2398 3192
rect 2545 3187 2646 3192
rect 2393 3182 2422 3187
rect 2457 3182 2550 3187
rect 2641 3182 2758 3187
rect 3009 3182 3158 3187
rect 3265 3182 3286 3187
rect 3377 3182 3494 3187
rect 3737 3182 3846 3187
rect 4489 3182 4598 3187
rect 449 3177 550 3182
rect 889 3177 958 3182
rect 1817 3177 1886 3182
rect 2001 3177 2182 3182
rect 2777 3177 3014 3182
rect 3153 3177 3158 3182
rect 4593 3177 4598 3182
rect 4761 3182 4806 3187
rect 4761 3177 4766 3182
rect 369 3172 454 3177
rect 545 3172 638 3177
rect 761 3172 798 3177
rect 1121 3172 1238 3177
rect 1505 3172 1822 3177
rect 1881 3172 2006 3177
rect 2177 3172 2454 3177
rect 2489 3172 2550 3177
rect 2609 3172 2782 3177
rect 3153 3172 3518 3177
rect 3537 3172 3638 3177
rect 3657 3172 3782 3177
rect 4593 3172 4766 3177
rect 3537 3167 3542 3172
rect 345 3162 526 3167
rect 737 3162 1398 3167
rect 1577 3162 1606 3167
rect 1793 3162 1870 3167
rect 2017 3162 2094 3167
rect 2113 3162 2406 3167
rect 2625 3162 2958 3167
rect 3049 3162 3078 3167
rect 3257 3162 3294 3167
rect 3385 3162 3542 3167
rect 3633 3167 3638 3172
rect 3633 3162 3734 3167
rect 1625 3157 1766 3162
rect 1889 3157 1998 3162
rect 2425 3157 2606 3162
rect 2953 3157 3054 3162
rect 3113 3157 3222 3162
rect 3753 3157 3838 3162
rect 297 3152 454 3157
rect 1081 3152 1134 3157
rect 1209 3152 1310 3157
rect 1305 3147 1310 3152
rect 1409 3152 1630 3157
rect 1761 3152 1894 3157
rect 1993 3152 2430 3157
rect 2601 3152 2934 3157
rect 1409 3147 1414 3152
rect 2929 3147 2934 3152
rect 3089 3152 3118 3157
rect 3217 3152 3246 3157
rect 3089 3147 3094 3152
rect 3241 3147 3246 3152
rect 3305 3152 3406 3157
rect 3417 3152 3718 3157
rect 3729 3152 3758 3157
rect 3833 3152 3958 3157
rect 4193 3152 4262 3157
rect 4313 3152 4358 3157
rect 4465 3152 4574 3157
rect 3305 3147 3310 3152
rect 4193 3147 4198 3152
rect 321 3142 390 3147
rect 505 3142 590 3147
rect 505 3137 510 3142
rect 305 3132 510 3137
rect 585 3137 590 3142
rect 657 3137 662 3147
rect 961 3142 1030 3147
rect 1049 3142 1230 3147
rect 1249 3142 1286 3147
rect 1305 3142 1414 3147
rect 1569 3142 1630 3147
rect 1689 3142 1750 3147
rect 1873 3142 2118 3147
rect 2217 3142 2462 3147
rect 2473 3142 2622 3147
rect 2633 3142 2910 3147
rect 2929 3142 3094 3147
rect 3145 3142 3190 3147
rect 3241 3142 3310 3147
rect 3425 3142 3510 3147
rect 3617 3142 3822 3147
rect 3953 3142 4014 3147
rect 4065 3142 4198 3147
rect 4257 3147 4262 3152
rect 4465 3147 4470 3152
rect 4257 3142 4470 3147
rect 4489 3142 4542 3147
rect 961 3137 966 3142
rect 585 3132 662 3137
rect 681 3132 910 3137
rect 937 3132 966 3137
rect 1025 3137 1030 3142
rect 1025 3132 1078 3137
rect 1673 3132 1702 3137
rect 1721 3132 1806 3137
rect 1969 3132 1990 3137
rect 2073 3132 2198 3137
rect 2241 3132 2310 3137
rect 2577 3132 2750 3137
rect 3353 3132 3702 3137
rect 3841 3132 3934 3137
rect 4617 3132 4662 3137
rect 681 3127 686 3132
rect 241 3122 382 3127
rect 441 3122 686 3127
rect 905 3127 910 3132
rect 1097 3127 1310 3132
rect 2385 3127 2558 3132
rect 3721 3127 3846 3132
rect 3929 3127 4038 3132
rect 905 3122 1102 3127
rect 1305 3122 1422 3127
rect 1449 3122 1654 3127
rect 1825 3122 1918 3127
rect 2081 3122 2390 3127
rect 2553 3122 2646 3127
rect 2833 3122 2918 3127
rect 2937 3122 3270 3127
rect 3289 3122 3454 3127
rect 3601 3122 3726 3127
rect 4033 3122 4246 3127
rect 4345 3122 4390 3127
rect 4537 3122 4574 3127
rect 1449 3117 1454 3122
rect 1649 3117 1830 3122
rect 1913 3117 1918 3122
rect 1985 3117 2054 3122
rect 2937 3117 2942 3122
rect 233 3112 286 3117
rect 329 3112 358 3117
rect 353 3107 358 3112
rect 433 3112 758 3117
rect 433 3107 438 3112
rect 753 3107 758 3112
rect 865 3112 894 3117
rect 961 3112 1006 3117
rect 1033 3112 1118 3117
rect 1137 3112 1254 3117
rect 1265 3112 1294 3117
rect 865 3107 870 3112
rect 217 3102 278 3107
rect 353 3102 438 3107
rect 457 3102 518 3107
rect 633 3102 734 3107
rect 753 3102 870 3107
rect 1265 3092 1270 3112
rect 1289 3097 1294 3112
rect 1433 3112 1454 3117
rect 1913 3112 1990 3117
rect 2049 3112 2302 3117
rect 2401 3112 2942 3117
rect 3265 3117 3270 3122
rect 3473 3117 3582 3122
rect 3265 3112 3478 3117
rect 3577 3112 3918 3117
rect 3993 3112 4022 3117
rect 4289 3112 4446 3117
rect 1433 3097 1438 3112
rect 2297 3107 2406 3112
rect 2961 3107 3102 3112
rect 3913 3107 3998 3112
rect 1465 3102 1502 3107
rect 1521 3102 1798 3107
rect 1817 3102 1902 3107
rect 2001 3102 2038 3107
rect 2105 3102 2134 3107
rect 2201 3102 2278 3107
rect 2425 3102 2470 3107
rect 2561 3102 2630 3107
rect 2881 3102 2966 3107
rect 3097 3102 3126 3107
rect 3185 3102 3582 3107
rect 3697 3102 3782 3107
rect 4353 3102 4414 3107
rect 1289 3092 1438 3097
rect 1673 3092 1718 3097
rect 1801 3092 1910 3097
rect 2297 3092 2406 3097
rect 2913 3092 3134 3097
rect 3433 3092 3654 3097
rect 3673 3092 3718 3097
rect 3761 3092 4278 3097
rect 2297 3087 2302 3092
rect 2401 3087 2574 3092
rect 3153 3087 3334 3092
rect 4273 3087 4278 3092
rect 4457 3092 4814 3097
rect 4457 3087 4462 3092
rect 1657 3082 1790 3087
rect 1897 3082 2302 3087
rect 2569 3082 2598 3087
rect 2649 3082 2790 3087
rect 2809 3082 3102 3087
rect 3129 3082 3158 3087
rect 3329 3082 3422 3087
rect 3561 3082 3638 3087
rect 3713 3082 3830 3087
rect 4273 3082 4462 3087
rect 1785 3077 1902 3082
rect 2649 3077 2654 3082
rect 1497 3072 1646 3077
rect 1641 3067 1646 3072
rect 1929 3072 2334 3077
rect 2385 3072 2654 3077
rect 2785 3077 2790 3082
rect 2785 3072 3318 3077
rect 3441 3072 3542 3077
rect 1929 3067 1934 3072
rect 3337 3067 3446 3072
rect 3537 3067 3638 3072
rect 1001 3062 1038 3067
rect 1305 3062 1374 3067
rect 1393 3062 1534 3067
rect 1641 3062 1934 3067
rect 2241 3062 2550 3067
rect 2665 3062 2774 3067
rect 2921 3062 3342 3067
rect 3633 3062 4206 3067
rect 1305 3057 1310 3062
rect 89 3052 366 3057
rect 89 3037 94 3052
rect 65 3032 94 3037
rect 361 3037 366 3052
rect 833 3052 910 3057
rect 1241 3052 1310 3057
rect 1369 3057 1374 3062
rect 1369 3052 1414 3057
rect 833 3047 838 3052
rect 641 3042 838 3047
rect 905 3047 910 3052
rect 1529 3047 1534 3062
rect 1953 3057 2246 3062
rect 2545 3057 2670 3062
rect 2769 3057 2926 3062
rect 1953 3047 1958 3057
rect 2265 3052 2366 3057
rect 2385 3052 2526 3057
rect 2945 3052 3534 3057
rect 3545 3052 3622 3057
rect 4105 3052 4134 3057
rect 3705 3047 3782 3052
rect 4129 3047 4134 3052
rect 4217 3052 4582 3057
rect 4217 3047 4222 3052
rect 905 3042 1126 3047
rect 1321 3042 1374 3047
rect 1529 3042 1958 3047
rect 1977 3042 2254 3047
rect 2441 3042 2558 3047
rect 2577 3042 2742 3047
rect 2249 3037 2254 3042
rect 2329 3037 2446 3042
rect 2577 3037 2582 3042
rect 361 3032 446 3037
rect 1337 3032 1358 3037
rect 1393 3032 1446 3037
rect 2249 3032 2334 3037
rect 2465 3032 2582 3037
rect 2737 3037 2742 3042
rect 2785 3042 2870 3047
rect 2961 3042 3358 3047
rect 3633 3042 3710 3047
rect 3777 3042 3934 3047
rect 4129 3042 4222 3047
rect 2785 3037 2790 3042
rect 2737 3032 2790 3037
rect 2865 3037 2870 3042
rect 3353 3037 3358 3042
rect 3569 3037 3638 3042
rect 2865 3032 2894 3037
rect 2929 3032 2974 3037
rect 3041 3032 3086 3037
rect 3233 3032 3262 3037
rect 3353 3032 3574 3037
rect 3721 3032 3766 3037
rect 4705 3032 4766 3037
rect 1393 3027 1398 3032
rect 3081 3027 3238 3032
rect 4705 3027 4710 3032
rect 105 3022 350 3027
rect 537 3022 654 3027
rect 849 3022 894 3027
rect 969 3022 1270 3027
rect 1329 3022 1398 3027
rect 1417 3022 1510 3027
rect 1593 3022 1678 3027
rect 2353 3022 2406 3027
rect 2521 3022 2910 3027
rect 2993 3022 3062 3027
rect 3313 3022 3334 3027
rect 3593 3022 4190 3027
rect 4417 3022 4710 3027
rect 4729 3022 4758 3027
rect 1593 3017 1598 3022
rect 745 3012 774 3017
rect 1201 3012 1382 3017
rect 1409 3012 1518 3017
rect 1537 3012 1598 3017
rect 1673 3017 1678 3022
rect 2401 3017 2406 3022
rect 1673 3012 2166 3017
rect 2225 3007 2230 3017
rect 2401 3012 2534 3017
rect 2529 3007 2534 3012
rect 2673 3012 2750 3017
rect 2921 3012 2982 3017
rect 3073 3012 3214 3017
rect 2673 3007 2678 3012
rect 1257 3002 1350 3007
rect 1409 3002 1534 3007
rect 1609 3002 1686 3007
rect 2225 3002 2390 3007
rect 1529 2997 1614 3002
rect 2385 2997 2390 3002
rect 2481 3002 2510 3007
rect 2529 3002 2678 3007
rect 2745 3007 2750 3012
rect 2849 3007 2926 3012
rect 2977 3007 3078 3012
rect 2745 3002 2854 3007
rect 3313 3002 3318 3022
rect 3489 3012 3710 3017
rect 4257 3012 4310 3017
rect 3465 3002 3870 3007
rect 2481 2997 2486 3002
rect 81 2992 270 2997
rect 361 2992 438 2997
rect 505 2992 574 2997
rect 633 2992 662 2997
rect 865 2992 1022 2997
rect 1121 2992 1174 2997
rect 1265 2992 1318 2997
rect 1337 2992 1510 2997
rect 1665 2992 1726 2997
rect 1793 2992 1822 2997
rect 1817 2987 1822 2992
rect 1905 2992 1958 2997
rect 1905 2987 1910 2992
rect 329 2982 358 2987
rect 449 2982 502 2987
rect 1009 2982 1110 2987
rect 1361 2982 1446 2987
rect 1513 2982 1550 2987
rect 1617 2982 1694 2987
rect 1817 2982 1910 2987
rect 1953 2987 1958 2992
rect 2033 2992 2230 2997
rect 2385 2992 2486 2997
rect 2697 2992 2726 2997
rect 2873 2992 3038 2997
rect 3057 2992 3366 2997
rect 3425 2992 3478 2997
rect 3601 2992 3630 2997
rect 3689 2992 3726 2997
rect 3881 2992 4294 2997
rect 4321 2992 4326 3017
rect 4369 3012 4454 3017
rect 4657 3012 4726 3017
rect 4657 3007 4662 3012
rect 4545 3002 4662 3007
rect 4377 2992 4438 2997
rect 4561 2992 4654 2997
rect 2033 2987 2038 2992
rect 3881 2987 3886 2992
rect 1953 2982 2038 2987
rect 2057 2982 2102 2987
rect 1553 2972 1582 2977
rect 585 2962 782 2967
rect 801 2962 838 2967
rect 1673 2962 1718 2967
rect 2121 2962 2270 2967
rect 585 2957 590 2962
rect 241 2952 342 2957
rect 361 2952 502 2957
rect 561 2952 590 2957
rect 777 2957 782 2962
rect 2121 2957 2126 2962
rect 777 2952 894 2957
rect 1937 2952 2054 2957
rect 2089 2952 2126 2957
rect 2265 2957 2270 2962
rect 2289 2957 2294 2987
rect 3297 2982 3886 2987
rect 4057 2982 4086 2987
rect 4273 2982 4318 2987
rect 4385 2982 4662 2987
rect 2665 2977 2798 2982
rect 2449 2972 2670 2977
rect 2793 2972 2822 2977
rect 2905 2972 3030 2977
rect 3145 2972 3662 2977
rect 2681 2962 2798 2967
rect 2929 2962 2950 2967
rect 2969 2962 3134 2967
rect 3545 2962 3574 2967
rect 3977 2962 4046 2967
rect 2265 2952 2294 2957
rect 3129 2957 3134 2962
rect 3265 2957 3550 2962
rect 3129 2952 3270 2957
rect 4049 2952 4094 2957
rect 4113 2952 4398 2957
rect 361 2947 366 2952
rect 113 2942 182 2947
rect 265 2942 366 2947
rect 497 2947 502 2952
rect 1937 2947 1942 2952
rect 497 2942 702 2947
rect 697 2937 702 2942
rect 769 2942 846 2947
rect 897 2942 974 2947
rect 1081 2942 1126 2947
rect 1553 2942 1598 2947
rect 1617 2942 1766 2947
rect 1841 2942 1942 2947
rect 2049 2947 2054 2952
rect 2713 2947 2814 2952
rect 4049 2947 4054 2952
rect 4113 2947 4118 2952
rect 2049 2942 2078 2947
rect 2105 2942 2326 2947
rect 2473 2942 2526 2947
rect 2577 2942 2638 2947
rect 2689 2942 2718 2947
rect 2809 2942 2838 2947
rect 2865 2942 2958 2947
rect 3289 2942 3318 2947
rect 3425 2942 3462 2947
rect 3473 2942 3590 2947
rect 3649 2942 3702 2947
rect 3945 2942 4054 2947
rect 4073 2942 4118 2947
rect 4393 2947 4398 2952
rect 4585 2952 4734 2957
rect 4585 2947 4590 2952
rect 4393 2942 4590 2947
rect 4729 2947 4734 2952
rect 4729 2942 4790 2947
rect 769 2937 774 2942
rect 2689 2937 2694 2942
rect 3425 2937 3430 2942
rect 145 2932 190 2937
rect 313 2932 462 2937
rect 697 2932 774 2937
rect 953 2932 1126 2937
rect 1577 2932 1638 2937
rect 2257 2932 2294 2937
rect 2337 2932 2358 2937
rect 2489 2932 2518 2937
rect 2545 2932 2694 2937
rect 2705 2932 2902 2937
rect 3073 2932 3430 2937
rect 3745 2932 3790 2937
rect 3865 2932 3966 2937
rect 4201 2932 4382 2937
rect 3609 2927 3726 2932
rect 193 2922 222 2927
rect 193 2917 198 2922
rect 177 2912 198 2917
rect 217 2907 222 2922
rect 457 2922 486 2927
rect 953 2922 998 2927
rect 1457 2922 1526 2927
rect 1545 2922 1750 2927
rect 1769 2922 1934 2927
rect 1953 2922 2126 2927
rect 2145 2922 2238 2927
rect 2281 2922 2310 2927
rect 2321 2922 2398 2927
rect 2633 2922 2718 2927
rect 3297 2922 3358 2927
rect 3585 2922 3614 2927
rect 3721 2922 3838 2927
rect 4089 2922 4142 2927
rect 4601 2922 4718 2927
rect 457 2907 462 2922
rect 1457 2917 1462 2922
rect 881 2912 926 2917
rect 1025 2912 1142 2917
rect 1257 2912 1462 2917
rect 1521 2917 1526 2922
rect 1769 2917 1774 2922
rect 1521 2912 1774 2917
rect 1929 2917 1934 2922
rect 2145 2917 2150 2922
rect 1929 2912 2150 2917
rect 2233 2917 2238 2922
rect 2473 2917 2614 2922
rect 2897 2917 2966 2922
rect 2233 2912 2278 2917
rect 2369 2912 2478 2917
rect 2609 2912 2670 2917
rect 2729 2912 2902 2917
rect 2961 2912 3286 2917
rect 2273 2907 2374 2912
rect 2665 2907 2734 2912
rect 3281 2907 3286 2912
rect 3441 2912 3574 2917
rect 3441 2907 3446 2912
rect 217 2902 462 2907
rect 1105 2902 1158 2907
rect 1185 2902 1286 2907
rect 1473 2902 1510 2907
rect 1561 2902 1590 2907
rect 1585 2897 1590 2902
rect 1673 2902 1702 2907
rect 1713 2902 1918 2907
rect 1985 2902 2038 2907
rect 2161 2902 2254 2907
rect 2489 2902 2646 2907
rect 2913 2902 2950 2907
rect 3281 2902 3446 2907
rect 3569 2907 3574 2912
rect 3649 2912 4078 2917
rect 3649 2907 3654 2912
rect 4073 2907 4078 2912
rect 4153 2912 4278 2917
rect 4377 2912 4558 2917
rect 4697 2912 4758 2917
rect 4153 2907 4158 2912
rect 3569 2902 3654 2907
rect 3673 2902 3758 2907
rect 3841 2902 3870 2907
rect 4073 2902 4158 2907
rect 4217 2902 4246 2907
rect 4361 2902 4422 2907
rect 1673 2897 1678 2902
rect 1913 2897 1990 2902
rect 2033 2897 2166 2902
rect 2393 2897 2470 2902
rect 97 2892 118 2897
rect 1585 2892 1678 2897
rect 1705 2892 1734 2897
rect 1729 2887 1734 2892
rect 2233 2892 2398 2897
rect 2465 2892 2686 2897
rect 2233 2887 2238 2892
rect 3865 2887 3870 2902
rect 4217 2887 4222 2902
rect 4417 2897 4422 2902
rect 4545 2902 4590 2907
rect 4545 2897 4550 2902
rect 4417 2892 4550 2897
rect 1729 2882 2238 2887
rect 2409 2882 2470 2887
rect 2705 2882 2894 2887
rect 2553 2877 2710 2882
rect 2889 2877 2894 2882
rect 2969 2882 3062 2887
rect 3081 2882 3134 2887
rect 3153 2882 3326 2887
rect 3865 2882 4222 2887
rect 2969 2877 2974 2882
rect 785 2872 814 2877
rect 1401 2872 1686 2877
rect 2257 2872 2558 2877
rect 2889 2872 2974 2877
rect 3057 2877 3062 2882
rect 3153 2877 3158 2882
rect 3057 2872 3158 2877
rect 3321 2877 3326 2882
rect 3321 2872 3382 2877
rect 1401 2867 1406 2872
rect 1377 2862 1406 2867
rect 1681 2867 1686 2872
rect 1681 2862 1718 2867
rect 1737 2862 1990 2867
rect 2393 2862 2438 2867
rect 2569 2862 3198 2867
rect 1737 2857 1742 2862
rect 1257 2852 1342 2857
rect 1577 2852 1742 2857
rect 1985 2857 1990 2862
rect 2433 2857 2574 2862
rect 3193 2857 3198 2862
rect 3281 2862 3310 2867
rect 3281 2857 3286 2862
rect 1985 2852 2414 2857
rect 2593 2852 2622 2857
rect 2673 2852 2702 2857
rect 2873 2852 2990 2857
rect 3009 2852 3054 2857
rect 2697 2847 2878 2852
rect 3049 2847 3054 2852
rect 3145 2852 3174 2857
rect 3193 2852 3286 2857
rect 4281 2852 4398 2857
rect 3145 2847 3150 2852
rect 4281 2847 4286 2852
rect 185 2842 262 2847
rect 1345 2842 1558 2847
rect 1857 2842 1950 2847
rect 1857 2837 1862 2842
rect 257 2832 326 2837
rect 345 2832 422 2837
rect 649 2832 694 2837
rect 1281 2832 1350 2837
rect 345 2827 350 2832
rect 273 2822 302 2827
rect 313 2822 350 2827
rect 417 2827 422 2832
rect 1345 2827 1350 2832
rect 1545 2832 1710 2837
rect 1745 2832 1862 2837
rect 1945 2837 1950 2842
rect 2433 2842 2510 2847
rect 2897 2842 2934 2847
rect 2945 2842 3014 2847
rect 3049 2842 3150 2847
rect 4257 2842 4286 2847
rect 4393 2847 4398 2852
rect 4441 2852 4606 2857
rect 4393 2842 4422 2847
rect 2433 2837 2438 2842
rect 1945 2832 1974 2837
rect 2377 2832 2406 2837
rect 2417 2832 2438 2837
rect 2505 2837 2510 2842
rect 4441 2837 4446 2852
rect 4601 2837 4606 2852
rect 4625 2842 4718 2847
rect 2505 2832 2662 2837
rect 2713 2832 2790 2837
rect 2809 2832 2910 2837
rect 2945 2832 3030 2837
rect 3577 2832 3662 2837
rect 3833 2832 4334 2837
rect 4401 2832 4446 2837
rect 4465 2832 4582 2837
rect 4601 2832 4662 2837
rect 1545 2827 1550 2832
rect 1745 2827 1750 2832
rect 2417 2827 2422 2832
rect 2713 2827 2718 2832
rect 417 2822 446 2827
rect 585 2822 622 2827
rect 713 2822 742 2827
rect 801 2822 846 2827
rect 913 2822 1014 2827
rect 1297 2822 1326 2827
rect 1345 2822 1550 2827
rect 1697 2822 1750 2827
rect 1873 2822 1910 2827
rect 1953 2822 1982 2827
rect 2057 2822 2102 2827
rect 2265 2822 2302 2827
rect 2345 2822 2422 2827
rect 2433 2822 2494 2827
rect 2689 2822 2718 2827
rect 2785 2827 2790 2832
rect 2945 2827 2950 2832
rect 4465 2827 4470 2832
rect 2785 2822 2822 2827
rect 2833 2822 2950 2827
rect 3065 2822 3326 2827
rect 3345 2822 3374 2827
rect 3649 2822 3670 2827
rect 3689 2822 3798 2827
rect 3993 2822 4038 2827
rect 4129 2822 4470 2827
rect 4577 2827 4582 2832
rect 4577 2822 4870 2827
rect 617 2817 718 2822
rect 249 2812 598 2817
rect 753 2812 822 2817
rect 961 2812 998 2817
rect 177 2802 262 2807
rect 569 2802 638 2807
rect 681 2802 734 2807
rect 753 2797 758 2812
rect 777 2802 918 2807
rect 225 2792 294 2797
rect 737 2792 758 2797
rect 913 2792 966 2797
rect 121 2782 198 2787
rect 409 2782 446 2787
rect 593 2782 622 2787
rect 617 2777 622 2782
rect 729 2782 878 2787
rect 993 2782 998 2812
rect 1009 2797 1014 2822
rect 3065 2817 3070 2822
rect 1713 2812 1750 2817
rect 1865 2812 1894 2817
rect 2153 2812 2262 2817
rect 2553 2812 2886 2817
rect 3041 2812 3070 2817
rect 3321 2817 3326 2822
rect 3689 2817 3694 2822
rect 3321 2812 3366 2817
rect 3417 2812 3558 2817
rect 3585 2812 3694 2817
rect 3793 2817 3798 2822
rect 3793 2812 3862 2817
rect 3961 2812 4006 2817
rect 4129 2812 4286 2817
rect 1217 2802 1310 2807
rect 1569 2802 1614 2807
rect 1745 2802 1750 2812
rect 1889 2807 2038 2812
rect 2033 2802 2158 2807
rect 2177 2802 2222 2807
rect 2625 2802 2694 2807
rect 2833 2802 3102 2807
rect 3217 2802 3262 2807
rect 2625 2797 2630 2802
rect 3417 2797 3422 2812
rect 1009 2792 1102 2797
rect 1369 2792 1414 2797
rect 1609 2792 2054 2797
rect 2121 2792 2182 2797
rect 2521 2792 2630 2797
rect 2649 2792 2846 2797
rect 3145 2792 3182 2797
rect 3241 2792 3350 2797
rect 3393 2792 3422 2797
rect 3553 2797 3558 2812
rect 4281 2807 4286 2812
rect 4385 2812 4638 2817
rect 4385 2807 4390 2812
rect 3657 2802 3902 2807
rect 4025 2802 4070 2807
rect 4137 2802 4262 2807
rect 4281 2802 4390 2807
rect 4465 2802 4510 2807
rect 3553 2792 3670 2797
rect 3801 2792 3894 2797
rect 3985 2792 4062 2797
rect 4209 2792 4230 2797
rect 4409 2792 4446 2797
rect 4625 2792 4654 2797
rect 3689 2787 3782 2792
rect 1121 2782 1198 2787
rect 1537 2782 1638 2787
rect 1897 2782 1982 2787
rect 2393 2782 2510 2787
rect 729 2777 734 2782
rect 1793 2777 1878 2782
rect 2505 2777 2510 2782
rect 2737 2782 3694 2787
rect 3777 2782 4182 2787
rect 4281 2782 4374 2787
rect 4393 2782 4566 2787
rect 2737 2777 2742 2782
rect 4281 2777 4286 2782
rect 441 2772 478 2777
rect 617 2772 734 2777
rect 1529 2772 1558 2777
rect 1649 2772 1798 2777
rect 1873 2772 1966 2777
rect 2201 2772 2374 2777
rect 2505 2772 2742 2777
rect 2809 2772 2854 2777
rect 3233 2772 3270 2777
rect 3353 2772 3406 2777
rect 3633 2772 3854 2777
rect 4177 2772 4286 2777
rect 4369 2777 4374 2782
rect 4369 2772 4446 2777
rect 4753 2772 4782 2777
rect 1553 2767 1654 2772
rect 2201 2767 2206 2772
rect 753 2762 958 2767
rect 1225 2762 1302 2767
rect 1321 2762 1486 2767
rect 1809 2762 1910 2767
rect 1225 2757 1230 2762
rect 817 2752 862 2757
rect 1201 2752 1230 2757
rect 1297 2757 1302 2762
rect 1905 2757 1910 2762
rect 1985 2762 2206 2767
rect 2369 2767 2374 2772
rect 3849 2767 4022 2772
rect 4177 2767 4182 2772
rect 2369 2762 2438 2767
rect 2761 2762 2846 2767
rect 2937 2762 3214 2767
rect 3601 2762 3694 2767
rect 3801 2762 3830 2767
rect 4017 2762 4182 2767
rect 4201 2762 4390 2767
rect 1985 2757 1990 2762
rect 2937 2757 2942 2762
rect 3209 2757 3278 2762
rect 3689 2757 3806 2762
rect 1297 2752 1382 2757
rect 1473 2752 1678 2757
rect 1473 2747 1478 2752
rect 1673 2747 1678 2752
rect 1801 2752 1854 2757
rect 1905 2752 1990 2757
rect 2113 2752 2294 2757
rect 2353 2752 2382 2757
rect 2449 2752 2614 2757
rect 2633 2752 2742 2757
rect 2913 2752 2942 2757
rect 3273 2752 3598 2757
rect 3609 2752 3670 2757
rect 3913 2752 3998 2757
rect 4241 2752 4294 2757
rect 1801 2747 1806 2752
rect 2377 2747 2454 2752
rect 2633 2747 2638 2752
rect 89 2742 134 2747
rect 337 2742 374 2747
rect 393 2742 502 2747
rect 585 2742 646 2747
rect 833 2742 958 2747
rect 1177 2742 1478 2747
rect 1497 2742 1526 2747
rect 393 2737 398 2742
rect 329 2732 398 2737
rect 497 2737 502 2742
rect 1521 2737 1526 2742
rect 1625 2742 1654 2747
rect 1673 2742 1806 2747
rect 2009 2742 2046 2747
rect 2225 2742 2342 2747
rect 1625 2737 1630 2742
rect 2337 2737 2342 2742
rect 2553 2742 2638 2747
rect 2737 2747 2742 2752
rect 3097 2747 3182 2752
rect 3913 2747 3918 2752
rect 2737 2742 3102 2747
rect 3177 2742 3262 2747
rect 3601 2742 3630 2747
rect 3729 2742 3790 2747
rect 3889 2742 3918 2747
rect 3993 2747 3998 2752
rect 3993 2742 4230 2747
rect 2553 2737 2558 2742
rect 4225 2737 4230 2742
rect 4297 2742 4318 2747
rect 4297 2737 4302 2742
rect 497 2732 526 2737
rect 625 2732 670 2737
rect 745 2732 942 2737
rect 1225 2732 1350 2737
rect 1393 2732 1454 2737
rect 1521 2732 1630 2737
rect 1825 2732 1862 2737
rect 2073 2732 2134 2737
rect 2289 2732 2318 2737
rect 2337 2732 2558 2737
rect 2593 2732 2630 2737
rect 3017 2732 3046 2737
rect 409 2722 454 2727
rect 513 2722 534 2727
rect 433 2712 462 2717
rect 513 2707 518 2722
rect 561 2712 606 2717
rect 185 2702 366 2707
rect 513 2702 542 2707
rect 625 2702 630 2732
rect 2737 2727 2910 2732
rect 3041 2727 3046 2732
rect 3113 2732 3166 2737
rect 3385 2732 3926 2737
rect 3937 2732 3982 2737
rect 4225 2732 4302 2737
rect 4313 2737 4318 2742
rect 4401 2742 4526 2747
rect 4641 2742 4758 2747
rect 4401 2737 4406 2742
rect 4313 2732 4406 2737
rect 4617 2732 4646 2737
rect 3113 2727 3118 2732
rect 889 2722 966 2727
rect 985 2722 1030 2727
rect 1305 2722 1374 2727
rect 2577 2722 2614 2727
rect 2625 2722 2742 2727
rect 2905 2722 2934 2727
rect 3041 2722 3118 2727
rect 3137 2722 3174 2727
rect 3681 2722 3774 2727
rect 3857 2722 3926 2727
rect 2625 2717 2630 2722
rect 3553 2717 3622 2722
rect 3937 2717 3942 2732
rect 4161 2722 4198 2727
rect 705 2712 806 2717
rect 1337 2712 1358 2717
rect 1505 2712 1582 2717
rect 1857 2712 1926 2717
rect 1961 2712 2006 2717
rect 2041 2712 2086 2717
rect 2273 2712 2334 2717
rect 2409 2712 2630 2717
rect 2641 2712 2670 2717
rect 2753 2712 2886 2717
rect 3153 2712 3206 2717
rect 3489 2712 3558 2717
rect 3617 2712 3646 2717
rect 3857 2712 3942 2717
rect 4241 2712 4294 2717
rect 2665 2707 2758 2712
rect 3665 2707 3806 2712
rect 3857 2707 3862 2712
rect 689 2702 758 2707
rect 793 2702 886 2707
rect 1257 2702 1350 2707
rect 1857 2702 1958 2707
rect 2033 2702 2062 2707
rect 2433 2702 2518 2707
rect 2809 2702 2846 2707
rect 3161 2702 3214 2707
rect 3281 2702 3470 2707
rect 3569 2702 3670 2707
rect 3801 2702 3862 2707
rect 3873 2702 3918 2707
rect 4377 2702 4430 2707
rect 3281 2697 3286 2702
rect 3465 2697 3550 2702
rect 4273 2697 4342 2702
rect 321 2692 358 2697
rect 569 2692 622 2697
rect 617 2687 622 2692
rect 713 2692 742 2697
rect 1313 2692 1350 2697
rect 1969 2692 2078 2697
rect 2593 2692 2622 2697
rect 2665 2692 2710 2697
rect 2809 2692 2878 2697
rect 3089 2692 3174 2697
rect 3257 2692 3286 2697
rect 3545 2692 3638 2697
rect 713 2687 718 2692
rect 3633 2687 3638 2692
rect 3929 2692 4278 2697
rect 4337 2692 4366 2697
rect 545 2682 598 2687
rect 617 2682 718 2687
rect 1185 2682 1278 2687
rect 1673 2682 2046 2687
rect 2057 2682 2110 2687
rect 2121 2682 2470 2687
rect 3153 2682 3454 2687
rect 3449 2677 3454 2682
rect 3521 2682 3550 2687
rect 3633 2682 3662 2687
rect 3521 2677 3526 2682
rect 3657 2677 3790 2682
rect 3929 2677 3934 2692
rect 4361 2687 4366 2692
rect 4441 2692 4614 2697
rect 4441 2687 4446 2692
rect 4169 2682 4198 2687
rect 129 2672 286 2677
rect 1641 2672 1742 2677
rect 1921 2672 2030 2677
rect 3225 2672 3270 2677
rect 3449 2672 3526 2677
rect 3785 2672 3934 2677
rect 4193 2677 4198 2682
rect 4289 2682 4318 2687
rect 4361 2682 4446 2687
rect 4289 2677 4294 2682
rect 4193 2672 4294 2677
rect 1897 2662 2422 2667
rect 3569 2662 3766 2667
rect 4385 2662 4438 2667
rect 3569 2657 3574 2662
rect 433 2652 462 2657
rect 1057 2652 1214 2657
rect 1593 2652 1638 2657
rect 1761 2652 1878 2657
rect 1961 2652 1990 2657
rect 2169 2652 2198 2657
rect 2281 2652 2310 2657
rect 2617 2652 3158 2657
rect 1057 2647 1062 2652
rect 609 2642 638 2647
rect 833 2642 934 2647
rect 1033 2642 1062 2647
rect 1209 2647 1214 2652
rect 1761 2647 1766 2652
rect 1209 2642 1286 2647
rect 1633 2642 1766 2647
rect 1873 2647 1878 2652
rect 1985 2647 2174 2652
rect 2617 2647 2622 2652
rect 1873 2642 1926 2647
rect 2297 2642 2318 2647
rect 2337 2642 2622 2647
rect 305 2632 342 2637
rect 609 2632 702 2637
rect 953 2632 1198 2637
rect 1361 2632 1446 2637
rect 1769 2632 1854 2637
rect 121 2612 214 2617
rect 233 2612 310 2617
rect 121 2607 126 2612
rect 97 2602 126 2607
rect 209 2607 214 2612
rect 337 2607 342 2632
rect 1361 2627 1366 2632
rect 593 2622 718 2627
rect 1017 2622 1110 2627
rect 1289 2622 1366 2627
rect 1441 2627 1446 2632
rect 1921 2627 1926 2642
rect 2337 2637 2342 2642
rect 3153 2637 3158 2652
rect 3289 2652 3574 2657
rect 3289 2647 3294 2652
rect 3177 2642 3294 2647
rect 3761 2647 3766 2662
rect 4321 2652 4422 2657
rect 3761 2642 3790 2647
rect 3881 2642 4110 2647
rect 4129 2642 4294 2647
rect 3881 2637 3886 2642
rect 2017 2632 2342 2637
rect 2897 2632 3030 2637
rect 3153 2632 3358 2637
rect 2017 2627 2022 2632
rect 2897 2627 2902 2632
rect 1441 2622 1470 2627
rect 1489 2622 1566 2627
rect 1713 2622 1790 2627
rect 1841 2622 1886 2627
rect 1921 2622 2022 2627
rect 2345 2622 2454 2627
rect 2513 2622 2598 2627
rect 2633 2622 2702 2627
rect 2793 2622 2902 2627
rect 3025 2627 3030 2632
rect 3353 2627 3358 2632
rect 3481 2632 3886 2637
rect 4105 2637 4110 2642
rect 4105 2632 4190 2637
rect 4577 2632 4710 2637
rect 3481 2627 3486 2632
rect 3025 2622 3158 2627
rect 3241 2622 3286 2627
rect 3353 2622 3486 2627
rect 3897 2622 3934 2627
rect 4097 2622 4158 2627
rect 4585 2622 4614 2627
rect 1489 2617 1494 2622
rect 785 2612 806 2617
rect 977 2612 1006 2617
rect 1001 2607 1006 2612
rect 1105 2612 1494 2617
rect 1561 2617 1566 2622
rect 2513 2617 2518 2622
rect 1561 2612 1630 2617
rect 2177 2612 2230 2617
rect 2457 2612 2518 2617
rect 2593 2617 2598 2622
rect 2593 2612 2790 2617
rect 2913 2612 3014 2617
rect 3169 2612 3198 2617
rect 3505 2612 3526 2617
rect 3929 2612 3982 2617
rect 4001 2612 4126 2617
rect 4257 2612 4286 2617
rect 1105 2607 1110 2612
rect 3049 2607 3150 2612
rect 3217 2607 3310 2612
rect 209 2602 246 2607
rect 313 2602 342 2607
rect 377 2602 486 2607
rect 585 2602 718 2607
rect 1001 2602 1110 2607
rect 1289 2602 1390 2607
rect 1481 2602 1550 2607
rect 1849 2602 1886 2607
rect 2041 2602 2110 2607
rect 2161 2602 2206 2607
rect 2529 2602 2902 2607
rect 2529 2597 2534 2602
rect 2897 2597 2902 2602
rect 3025 2602 3054 2607
rect 3145 2602 3222 2607
rect 3305 2602 3334 2607
rect 3025 2597 3030 2602
rect 4257 2597 4262 2612
rect 4345 2602 4390 2607
rect 217 2592 390 2597
rect 489 2592 662 2597
rect 657 2587 662 2592
rect 729 2592 958 2597
rect 1129 2592 1246 2597
rect 1329 2592 1366 2597
rect 1801 2592 1918 2597
rect 2177 2592 2222 2597
rect 2249 2592 2438 2597
rect 2505 2592 2534 2597
rect 2569 2592 2630 2597
rect 2641 2592 2742 2597
rect 2897 2592 3030 2597
rect 3073 2592 3158 2597
rect 3193 2592 3310 2597
rect 3609 2592 3790 2597
rect 3809 2592 3942 2597
rect 4089 2592 4238 2597
rect 4257 2592 4286 2597
rect 4369 2592 4406 2597
rect 4441 2592 4486 2597
rect 729 2587 734 2592
rect 1417 2587 1582 2592
rect 89 2582 302 2587
rect 337 2582 478 2587
rect 513 2582 638 2587
rect 657 2582 734 2587
rect 1345 2582 1382 2587
rect 1393 2582 1422 2587
rect 1577 2582 1606 2587
rect 1625 2582 1782 2587
rect 2249 2582 2254 2592
rect 1393 2577 1398 2582
rect 1625 2577 1630 2582
rect 225 2572 294 2577
rect 345 2572 438 2577
rect 1305 2572 1398 2577
rect 1417 2572 1630 2577
rect 1777 2577 1782 2582
rect 2145 2577 2254 2582
rect 2433 2577 2438 2592
rect 2465 2582 2614 2587
rect 3265 2582 3414 2587
rect 3513 2582 3590 2587
rect 3113 2577 3190 2582
rect 3609 2577 3614 2592
rect 1777 2572 1846 2577
rect 1857 2572 2150 2577
rect 2433 2572 3118 2577
rect 3185 2572 3614 2577
rect 3785 2577 3790 2592
rect 4345 2582 4478 2587
rect 4513 2582 4782 2587
rect 3785 2572 3822 2577
rect 3961 2572 4070 2577
rect 3961 2567 3966 2572
rect 49 2562 78 2567
rect 113 2562 1014 2567
rect 1265 2562 1510 2567
rect 1689 2562 1862 2567
rect 2065 2562 2094 2567
rect 49 2527 54 2562
rect 2089 2557 2094 2562
rect 2161 2562 2550 2567
rect 3129 2562 3174 2567
rect 3281 2562 3494 2567
rect 3593 2562 3774 2567
rect 3833 2562 3966 2567
rect 4065 2567 4070 2572
rect 4065 2562 4414 2567
rect 2161 2557 2166 2562
rect 3769 2557 3838 2562
rect 73 2552 198 2557
rect 1249 2552 1502 2557
rect 1601 2552 1806 2557
rect 2089 2552 2166 2557
rect 2593 2552 2654 2557
rect 3089 2552 3542 2557
rect 4249 2552 4278 2557
rect 4481 2552 4518 2557
rect 4561 2552 4638 2557
rect 2593 2547 2598 2552
rect 3561 2547 3630 2552
rect 4337 2547 4414 2552
rect 4561 2547 4566 2552
rect 177 2542 334 2547
rect 409 2542 438 2547
rect 729 2542 862 2547
rect 1001 2542 1038 2547
rect 1465 2542 1614 2547
rect 2353 2542 2462 2547
rect 2489 2542 2622 2547
rect 2633 2542 2790 2547
rect 3057 2542 3134 2547
rect 3201 2542 3566 2547
rect 3625 2542 3726 2547
rect 3785 2542 3886 2547
rect 3913 2542 4230 2547
rect 4265 2542 4342 2547
rect 4409 2542 4470 2547
rect 4537 2542 4566 2547
rect 4577 2542 4614 2547
rect 1281 2537 1414 2542
rect 4465 2537 4542 2542
rect 97 2532 190 2537
rect 281 2532 342 2537
rect 609 2532 782 2537
rect 817 2532 1110 2537
rect 1257 2532 1286 2537
rect 1409 2532 1590 2537
rect 1825 2532 1990 2537
rect 3105 2532 3246 2537
rect 3273 2532 3302 2537
rect 3537 2532 3614 2537
rect 4233 2532 4310 2537
rect 4369 2532 4398 2537
rect 1825 2527 1830 2532
rect 0 2522 54 2527
rect 81 2522 110 2527
rect 49 2517 54 2522
rect 49 2512 86 2517
rect 105 2507 110 2522
rect 297 2522 326 2527
rect 961 2522 1086 2527
rect 1249 2522 1398 2527
rect 1481 2522 1510 2527
rect 1545 2522 1830 2527
rect 1985 2527 1990 2532
rect 3321 2527 3518 2532
rect 3633 2527 4054 2532
rect 4369 2527 4374 2532
rect 1985 2522 2014 2527
rect 2145 2522 2262 2527
rect 2513 2522 2758 2527
rect 2865 2522 2918 2527
rect 3049 2522 3326 2527
rect 3513 2522 3558 2527
rect 3585 2522 3638 2527
rect 4049 2522 4206 2527
rect 4313 2522 4374 2527
rect 4497 2522 4518 2527
rect 4633 2522 4686 2527
rect 297 2507 302 2522
rect 1249 2517 1254 2522
rect 353 2512 430 2517
rect 609 2512 638 2517
rect 633 2507 638 2512
rect 785 2512 814 2517
rect 857 2512 942 2517
rect 953 2512 1014 2517
rect 1177 2512 1254 2517
rect 1281 2512 1334 2517
rect 1681 2512 1766 2517
rect 2153 2512 2190 2517
rect 2497 2512 2542 2517
rect 2673 2512 2886 2517
rect 2937 2512 3030 2517
rect 3097 2512 3230 2517
rect 3329 2512 3590 2517
rect 3609 2512 3734 2517
rect 3745 2512 3782 2517
rect 3809 2512 4038 2517
rect 4217 2512 4246 2517
rect 4305 2512 4342 2517
rect 4393 2512 4438 2517
rect 4561 2512 4678 2517
rect 785 2507 790 2512
rect 2937 2507 2942 2512
rect 105 2502 302 2507
rect 433 2502 542 2507
rect 633 2502 790 2507
rect 1001 2502 1046 2507
rect 1145 2502 1198 2507
rect 1305 2502 1334 2507
rect 1329 2497 1334 2502
rect 1409 2502 1518 2507
rect 1841 2502 2134 2507
rect 1409 2497 1414 2502
rect 2129 2497 2134 2502
rect 2201 2502 2486 2507
rect 2553 2502 2654 2507
rect 2665 2502 2702 2507
rect 2873 2502 2942 2507
rect 3025 2507 3030 2512
rect 3585 2507 3590 2512
rect 4305 2507 4310 2512
rect 3025 2502 3446 2507
rect 3545 2502 3574 2507
rect 3585 2502 3718 2507
rect 3873 2502 3918 2507
rect 4105 2502 4166 2507
rect 2201 2497 2206 2502
rect 2481 2497 2558 2502
rect 3441 2497 3550 2502
rect 3713 2497 3878 2502
rect 4161 2497 4166 2502
rect 4249 2502 4310 2507
rect 4329 2502 4406 2507
rect 4641 2502 4710 2507
rect 4249 2497 4254 2502
rect 1329 2492 1414 2497
rect 1721 2492 1758 2497
rect 2129 2492 2206 2497
rect 3121 2492 3222 2497
rect 3377 2492 3422 2497
rect 3625 2492 3694 2497
rect 4081 2492 4142 2497
rect 4161 2492 4254 2497
rect 4337 2492 4582 2497
rect 4617 2492 4662 2497
rect 2833 2487 2974 2492
rect 1737 2482 2022 2487
rect 2433 2482 2838 2487
rect 2969 2482 3158 2487
rect 3153 2477 3158 2482
rect 3241 2482 3358 2487
rect 3417 2482 3838 2487
rect 3241 2477 3246 2482
rect 1449 2472 1702 2477
rect 2225 2472 2318 2477
rect 2849 2472 2958 2477
rect 3153 2472 3246 2477
rect 3353 2477 3358 2482
rect 3833 2477 3838 2482
rect 3913 2482 4030 2487
rect 4289 2482 4326 2487
rect 3913 2477 3918 2482
rect 3353 2472 3614 2477
rect 3633 2472 3814 2477
rect 3833 2472 3918 2477
rect 4321 2477 4326 2482
rect 4401 2482 4430 2487
rect 4401 2477 4406 2482
rect 4321 2472 4406 2477
rect 1449 2457 1454 2472
rect 201 2452 366 2457
rect 481 2452 598 2457
rect 297 2442 438 2447
rect 481 2437 486 2452
rect 593 2447 598 2452
rect 1185 2452 1406 2457
rect 1425 2452 1454 2457
rect 1697 2457 1702 2472
rect 1961 2462 2214 2467
rect 2329 2462 3526 2467
rect 2209 2457 2334 2462
rect 3521 2457 3526 2462
rect 3681 2462 3814 2467
rect 4449 2462 4606 2467
rect 3681 2457 3686 2462
rect 4449 2457 4454 2462
rect 1697 2452 1886 2457
rect 2873 2452 2934 2457
rect 3169 2452 3430 2457
rect 3449 2452 3502 2457
rect 3521 2452 3686 2457
rect 3705 2452 3790 2457
rect 4353 2452 4454 2457
rect 4601 2457 4606 2462
rect 4601 2452 4758 2457
rect 1185 2447 1190 2452
rect 593 2442 1070 2447
rect 1161 2442 1190 2447
rect 1401 2447 1406 2452
rect 2633 2447 2822 2452
rect 1401 2442 1734 2447
rect 1841 2442 1934 2447
rect 2049 2442 2086 2447
rect 2105 2442 2174 2447
rect 2249 2442 2414 2447
rect 2489 2442 2518 2447
rect 2609 2442 2638 2447
rect 2817 2442 2950 2447
rect 4121 2442 4174 2447
rect 4409 2442 4590 2447
rect 1729 2437 1734 2442
rect 2105 2437 2110 2442
rect 321 2432 486 2437
rect 497 2432 526 2437
rect 1041 2432 1174 2437
rect 1433 2432 1502 2437
rect 1729 2432 1878 2437
rect 1873 2427 1878 2432
rect 1945 2432 2110 2437
rect 2169 2437 2174 2442
rect 3193 2437 3342 2442
rect 3449 2437 3526 2442
rect 4289 2437 4390 2442
rect 2169 2432 2238 2437
rect 2313 2432 2366 2437
rect 1945 2427 1950 2432
rect 2233 2427 2318 2432
rect 2361 2427 2366 2432
rect 2425 2432 2806 2437
rect 2961 2432 3198 2437
rect 3337 2432 3454 2437
rect 3521 2432 3694 2437
rect 2425 2427 2430 2432
rect 2801 2427 2966 2432
rect 3689 2427 3694 2432
rect 3777 2432 4294 2437
rect 4385 2432 4502 2437
rect 3777 2427 3782 2432
rect 377 2422 438 2427
rect 521 2422 582 2427
rect 1009 2422 1062 2427
rect 1217 2422 1374 2427
rect 1417 2422 1614 2427
rect 1873 2422 1950 2427
rect 2057 2422 2158 2427
rect 2337 2417 2342 2427
rect 2361 2422 2430 2427
rect 2505 2422 2614 2427
rect 2625 2422 2694 2427
rect 2721 2422 2782 2427
rect 3209 2422 3326 2427
rect 3465 2422 3510 2427
rect 3689 2422 3782 2427
rect 3801 2422 3838 2427
rect 4113 2422 4158 2427
rect 4305 2422 4438 2427
rect 4561 2422 4710 2427
rect 4729 2422 4758 2427
rect 1441 2412 1478 2417
rect 1825 2412 1854 2417
rect 2001 2412 2070 2417
rect 2241 2412 2342 2417
rect 2617 2412 2686 2417
rect 2737 2412 2934 2417
rect 3033 2412 3190 2417
rect 3265 2412 3310 2417
rect 3489 2412 3614 2417
rect 313 2402 342 2407
rect 561 2402 638 2407
rect 825 2402 862 2407
rect 1345 2402 1390 2407
rect 1465 2402 1566 2407
rect 1777 2402 1862 2407
rect 1977 2402 2006 2407
rect 2041 2402 2102 2407
rect 2217 2402 2254 2407
rect 2361 2402 2438 2407
rect 2273 2397 2366 2402
rect 2433 2397 2438 2402
rect 2633 2397 2766 2402
rect 3113 2397 3190 2402
rect 3265 2397 3270 2412
rect 3401 2402 3598 2407
rect 3937 2397 3942 2417
rect 4041 2407 4046 2417
rect 4393 2412 4446 2417
rect 4545 2412 4630 2417
rect 4705 2407 4710 2422
rect 4737 2412 4758 2417
rect 4017 2402 4046 2407
rect 4289 2402 4310 2407
rect 4377 2402 4406 2407
rect 4425 2402 4574 2407
rect 4585 2402 4606 2407
rect 4657 2402 4686 2407
rect 4705 2402 4734 2407
rect 4753 2397 4758 2412
rect 201 2392 270 2397
rect 345 2392 366 2397
rect 625 2392 742 2397
rect 873 2392 1006 2397
rect 1233 2392 1254 2397
rect 1273 2392 1358 2397
rect 1497 2392 1582 2397
rect 1785 2392 1814 2397
rect 1377 2387 1470 2392
rect 1809 2387 1814 2392
rect 1873 2392 2278 2397
rect 2433 2392 2638 2397
rect 2761 2392 2806 2397
rect 3049 2392 3118 2397
rect 3185 2392 3270 2397
rect 3305 2392 3342 2397
rect 3433 2392 3462 2397
rect 3553 2392 3606 2397
rect 3841 2392 3902 2397
rect 3937 2392 4142 2397
rect 4353 2392 4422 2397
rect 4625 2392 4654 2397
rect 4673 2392 4710 2397
rect 4737 2392 4758 2397
rect 1873 2387 1878 2392
rect 489 2382 622 2387
rect 1209 2382 1382 2387
rect 1465 2382 1670 2387
rect 1809 2382 1878 2387
rect 1977 2382 2054 2387
rect 2265 2382 2318 2387
rect 2313 2377 2318 2382
rect 2377 2382 2422 2387
rect 2649 2382 2758 2387
rect 3153 2382 3174 2387
rect 3329 2382 3358 2387
rect 2377 2377 2382 2382
rect 3353 2377 3358 2382
rect 3505 2382 3534 2387
rect 3553 2382 3670 2387
rect 3873 2382 3926 2387
rect 4345 2382 4414 2387
rect 4545 2382 4574 2387
rect 3505 2377 3510 2382
rect 4569 2377 4574 2382
rect 4649 2382 4702 2387
rect 4721 2382 4766 2387
rect 4649 2377 4654 2382
rect 1233 2372 1454 2377
rect 1609 2372 1646 2377
rect 2073 2372 2294 2377
rect 2313 2372 2382 2377
rect 2681 2372 2814 2377
rect 3353 2372 3510 2377
rect 4081 2372 4198 2377
rect 4289 2372 4318 2377
rect 4489 2372 4542 2377
rect 4569 2372 4654 2377
rect 4673 2372 4718 2377
rect 1449 2367 1614 2372
rect 641 2362 726 2367
rect 1249 2362 1430 2367
rect 1633 2362 1710 2367
rect 2233 2362 2262 2367
rect 2441 2362 2582 2367
rect 4065 2362 4342 2367
rect 4449 2362 4486 2367
rect 641 2357 646 2362
rect 577 2352 646 2357
rect 721 2357 726 2362
rect 1633 2357 1638 2362
rect 2113 2357 2214 2362
rect 2441 2357 2446 2362
rect 721 2352 750 2357
rect 1529 2352 1638 2357
rect 1705 2352 1814 2357
rect 1905 2352 1974 2357
rect 2089 2352 2118 2357
rect 2209 2352 2318 2357
rect 2417 2352 2446 2357
rect 2577 2357 2582 2362
rect 2577 2352 2606 2357
rect 2689 2352 2766 2357
rect 3241 2352 3318 2357
rect 3529 2352 3590 2357
rect 3609 2352 3726 2357
rect 3801 2352 3838 2357
rect 3961 2352 3990 2357
rect 4233 2352 4334 2357
rect 1377 2347 1470 2352
rect 3241 2347 3246 2352
rect 193 2342 278 2347
rect 321 2342 374 2347
rect 393 2342 462 2347
rect 569 2342 638 2347
rect 769 2342 950 2347
rect 985 2342 1070 2347
rect 1089 2342 1382 2347
rect 1465 2342 1518 2347
rect 1649 2342 1742 2347
rect 393 2337 398 2342
rect 297 2332 398 2337
rect 457 2337 462 2342
rect 769 2337 774 2342
rect 1513 2337 1654 2342
rect 1737 2337 1742 2342
rect 1825 2342 2270 2347
rect 2329 2342 2678 2347
rect 1825 2337 1830 2342
rect 2265 2337 2334 2342
rect 2673 2337 2678 2342
rect 2777 2342 3246 2347
rect 3313 2347 3318 2352
rect 3609 2347 3614 2352
rect 3313 2342 3614 2347
rect 3721 2347 3726 2352
rect 4009 2347 4150 2352
rect 3721 2342 3790 2347
rect 3849 2342 4014 2347
rect 4145 2342 4222 2347
rect 4321 2342 4350 2347
rect 2777 2337 2782 2342
rect 3785 2337 3854 2342
rect 4217 2337 4326 2342
rect 457 2332 774 2337
rect 873 2332 998 2337
rect 1393 2332 1454 2337
rect 1737 2332 1830 2337
rect 1865 2332 2006 2337
rect 2089 2332 2118 2337
rect 2137 2332 2246 2337
rect 2609 2332 2630 2337
rect 2673 2332 2782 2337
rect 3113 2332 3142 2337
rect 3481 2332 3630 2337
rect 3889 2332 4134 2337
rect 4425 2332 4446 2337
rect 2001 2327 2094 2332
rect 121 2322 158 2327
rect 513 2322 550 2327
rect 849 2322 878 2327
rect 969 2322 1070 2327
rect 1089 2322 1262 2327
rect 1321 2322 1462 2327
rect 1569 2322 1638 2327
rect 1945 2322 1982 2327
rect 2161 2322 2270 2327
rect 297 2317 494 2322
rect 569 2317 654 2322
rect 873 2317 974 2322
rect 1089 2317 1094 2322
rect 273 2312 302 2317
rect 489 2312 574 2317
rect 649 2312 790 2317
rect 273 2307 278 2312
rect 785 2307 790 2312
rect 993 2312 1094 2317
rect 1257 2317 1262 2322
rect 1569 2317 1574 2322
rect 1257 2312 1374 2317
rect 993 2307 998 2312
rect 1369 2307 1374 2312
rect 1473 2312 1574 2317
rect 1633 2317 1638 2322
rect 2265 2317 2270 2322
rect 2385 2322 2566 2327
rect 3257 2322 3302 2327
rect 3529 2322 3710 2327
rect 3825 2322 3894 2327
rect 3905 2322 3966 2327
rect 4001 2322 4022 2327
rect 4249 2322 4334 2327
rect 4585 2322 4718 2327
rect 2385 2317 2390 2322
rect 1633 2312 1718 2317
rect 1857 2312 2150 2317
rect 1473 2307 1478 2312
rect 137 2302 278 2307
rect 297 2302 358 2307
rect 377 2302 438 2307
rect 473 2302 638 2307
rect 737 2302 766 2307
rect 785 2302 998 2307
rect 1017 2302 1110 2307
rect 1145 2302 1246 2307
rect 1369 2302 1478 2307
rect 1585 2302 1622 2307
rect 1713 2302 1718 2312
rect 2145 2307 2150 2312
rect 2217 2312 2246 2317
rect 2265 2312 2390 2317
rect 2489 2312 2534 2317
rect 2609 2312 2638 2317
rect 2849 2312 2910 2317
rect 3113 2312 3318 2317
rect 3441 2312 3494 2317
rect 3649 2312 3958 2317
rect 3977 2312 4198 2317
rect 4217 2312 4254 2317
rect 4353 2312 4470 2317
rect 4697 2312 4758 2317
rect 2217 2307 2222 2312
rect 2145 2302 2222 2307
rect 2505 2302 2558 2307
rect 2977 2302 3094 2307
rect 3313 2302 3358 2307
rect 3481 2302 3694 2307
rect 3705 2302 3734 2307
rect 3753 2302 4390 2307
rect 2977 2297 2982 2302
rect 113 2292 262 2297
rect 321 2292 366 2297
rect 417 2292 558 2297
rect 697 2292 758 2297
rect 1265 2292 1350 2297
rect 2025 2292 2110 2297
rect 2729 2292 2830 2297
rect 2953 2292 2982 2297
rect 3089 2297 3094 2302
rect 4385 2297 4390 2302
rect 4481 2302 4638 2307
rect 4481 2297 4486 2302
rect 3089 2292 3390 2297
rect 3665 2292 3718 2297
rect 3953 2292 4030 2297
rect 4041 2292 4366 2297
rect 4385 2292 4486 2297
rect 1265 2287 1270 2292
rect 297 2282 510 2287
rect 1225 2282 1270 2287
rect 1345 2287 1350 2292
rect 2729 2287 2734 2292
rect 1345 2282 2014 2287
rect 2009 2277 2014 2282
rect 2121 2282 2734 2287
rect 2825 2287 2830 2292
rect 3737 2287 3934 2292
rect 2825 2282 3126 2287
rect 3257 2282 3310 2287
rect 3401 2282 3742 2287
rect 3929 2282 4246 2287
rect 2121 2277 2126 2282
rect 3121 2277 3262 2282
rect 3305 2277 3406 2282
rect 81 2272 110 2277
rect 521 2272 694 2277
rect 777 2272 1054 2277
rect 1217 2272 1334 2277
rect 2009 2272 2126 2277
rect 2745 2272 2798 2277
rect 105 2267 110 2272
rect 241 2267 526 2272
rect 105 2262 246 2267
rect 777 2262 782 2272
rect 625 2257 782 2262
rect 1049 2257 1054 2272
rect 2793 2267 2798 2272
rect 2921 2272 3102 2277
rect 2921 2267 2926 2272
rect 3097 2267 3102 2272
rect 3633 2272 3686 2277
rect 3633 2267 3638 2272
rect 1553 2262 1774 2267
rect 1553 2257 1558 2262
rect 265 2252 454 2257
rect 449 2247 454 2252
rect 601 2252 630 2257
rect 929 2252 1014 2257
rect 1049 2252 1558 2257
rect 1769 2257 1774 2262
rect 2153 2262 2246 2267
rect 2153 2257 2158 2262
rect 1769 2252 1798 2257
rect 1817 2252 2102 2257
rect 2129 2252 2158 2257
rect 2241 2257 2246 2262
rect 2441 2262 2686 2267
rect 2793 2262 2926 2267
rect 2945 2262 3006 2267
rect 3097 2262 3638 2267
rect 2441 2257 2446 2262
rect 2241 2252 2270 2257
rect 2385 2252 2446 2257
rect 2681 2257 2686 2262
rect 3681 2257 3686 2272
rect 4153 2272 4206 2277
rect 4153 2257 4158 2272
rect 2681 2252 2710 2257
rect 3681 2252 4158 2257
rect 4201 2257 4206 2272
rect 4377 2272 4630 2277
rect 4377 2257 4382 2272
rect 4529 2257 4622 2262
rect 4201 2252 4382 2257
rect 4505 2252 4534 2257
rect 4617 2252 4790 2257
rect 601 2247 606 2252
rect 929 2247 934 2252
rect 449 2242 606 2247
rect 625 2242 934 2247
rect 1009 2247 1014 2252
rect 1593 2247 1750 2252
rect 1817 2247 1822 2252
rect 1009 2242 1038 2247
rect 1569 2242 1598 2247
rect 1745 2242 1822 2247
rect 2097 2247 2102 2252
rect 2385 2247 2390 2252
rect 2097 2242 2126 2247
rect 2153 2242 2390 2247
rect 2457 2242 2670 2247
rect 2745 2242 2774 2247
rect 2953 2242 3078 2247
rect 3305 2242 3502 2247
rect 4553 2242 4606 2247
rect 1841 2237 2078 2242
rect 2665 2237 2750 2242
rect 3305 2237 3310 2242
rect 217 2232 310 2237
rect 361 2232 430 2237
rect 713 2232 782 2237
rect 945 2232 1078 2237
rect 1449 2232 1550 2237
rect 1577 2232 1846 2237
rect 2073 2232 2286 2237
rect 3049 2232 3126 2237
rect 3281 2232 3310 2237
rect 3497 2237 3502 2242
rect 3497 2232 3526 2237
rect 3593 2232 3662 2237
rect 3713 2232 3742 2237
rect 3761 2232 3806 2237
rect 3945 2232 4030 2237
rect 4297 2232 4318 2237
rect 4337 2232 4486 2237
rect 217 2227 222 2232
rect 193 2222 222 2227
rect 305 2227 310 2232
rect 1449 2227 1454 2232
rect 305 2222 374 2227
rect 905 2222 966 2227
rect 1145 2222 1334 2227
rect 1425 2222 1454 2227
rect 1545 2227 1550 2232
rect 4337 2227 4342 2232
rect 1545 2222 1614 2227
rect 1705 2222 1750 2227
rect 1809 2222 1942 2227
rect 1985 2222 2094 2227
rect 2185 2222 2262 2227
rect 2553 2222 2870 2227
rect 3033 2222 3062 2227
rect 3105 2222 3214 2227
rect 3241 2222 3278 2227
rect 3473 2222 3534 2227
rect 3585 2222 3758 2227
rect 3785 2222 3830 2227
rect 4017 2222 4062 2227
rect 4081 2222 4270 2227
rect 4289 2222 4342 2227
rect 4481 2227 4486 2232
rect 4481 2222 4510 2227
rect 4081 2217 4086 2222
rect 105 2212 294 2217
rect 425 2212 486 2217
rect 881 2212 958 2217
rect 1057 2212 1134 2217
rect 481 2207 486 2212
rect 113 2202 262 2207
rect 481 2202 558 2207
rect 1033 2202 1094 2207
rect 1129 2197 1134 2212
rect 1321 2212 1534 2217
rect 1625 2212 1694 2217
rect 1793 2212 1862 2217
rect 2073 2212 2542 2217
rect 2881 2212 3022 2217
rect 3289 2212 3678 2217
rect 3841 2212 4086 2217
rect 4265 2217 4270 2222
rect 4265 2212 4294 2217
rect 4353 2212 4470 2217
rect 4569 2212 4710 2217
rect 1321 2197 1326 2212
rect 1529 2207 1630 2212
rect 1689 2207 1798 2212
rect 1857 2207 2078 2212
rect 1817 2202 1838 2207
rect 2097 2202 2262 2207
rect 2537 2197 2542 2212
rect 2713 2207 2886 2212
rect 3017 2207 3294 2212
rect 3673 2207 3846 2212
rect 4289 2207 4358 2212
rect 2713 2197 2718 2207
rect 3505 2202 3534 2207
rect 3609 2202 3654 2207
rect 4033 2202 4126 2207
rect 4409 2202 4486 2207
rect 4529 2202 4566 2207
rect 817 2192 854 2197
rect 1129 2192 1326 2197
rect 1409 2192 1438 2197
rect 1561 2192 2086 2197
rect 2193 2192 2414 2197
rect 2537 2192 2718 2197
rect 2737 2192 3286 2197
rect 3457 2192 3502 2197
rect 3737 2192 3830 2197
rect 2081 2187 2198 2192
rect 3825 2187 3830 2192
rect 4081 2192 4294 2197
rect 4337 2192 4366 2197
rect 4481 2192 4590 2197
rect 4081 2187 4086 2192
rect 4481 2187 4486 2192
rect 145 2182 326 2187
rect 361 2182 462 2187
rect 361 2177 366 2182
rect 97 2172 134 2177
rect 337 2172 366 2177
rect 457 2177 462 2182
rect 577 2182 678 2187
rect 833 2182 878 2187
rect 2817 2182 2846 2187
rect 3297 2182 3382 2187
rect 3825 2182 4086 2187
rect 4329 2182 4358 2187
rect 4409 2182 4486 2187
rect 577 2177 582 2182
rect 457 2172 582 2177
rect 673 2177 678 2182
rect 1833 2177 1950 2182
rect 2841 2177 2846 2182
rect 2945 2177 3142 2182
rect 3297 2177 3302 2182
rect 673 2172 702 2177
rect 1345 2172 1838 2177
rect 1945 2172 2094 2177
rect 2153 2172 2318 2177
rect 2841 2172 2950 2177
rect 3137 2172 3302 2177
rect 4345 2172 4414 2177
rect 129 2167 134 2172
rect 209 2167 342 2172
rect 129 2162 214 2167
rect 1441 2162 1470 2167
rect 1761 2162 1934 2167
rect 2969 2162 3118 2167
rect 4185 2162 4310 2167
rect 4345 2162 4374 2167
rect 4433 2162 4478 2167
rect 1465 2157 1766 2162
rect 4185 2157 4190 2162
rect 233 2152 254 2157
rect 377 2152 518 2157
rect 561 2152 590 2157
rect 625 2152 678 2157
rect 945 2152 974 2157
rect 1785 2152 1814 2157
rect 1929 2152 2118 2157
rect 2297 2152 2318 2157
rect 3217 2152 3302 2157
rect 4161 2152 4190 2157
rect 4305 2157 4310 2162
rect 4305 2152 4510 2157
rect 4521 2152 4582 2157
rect 1809 2147 1934 2152
rect 3217 2147 3222 2152
rect 113 2142 206 2147
rect 297 2142 422 2147
rect 569 2142 630 2147
rect 1305 2142 1366 2147
rect 1377 2142 1534 2147
rect 1641 2142 1678 2147
rect 1953 2142 1974 2147
rect 2089 2142 2406 2147
rect 313 2132 366 2137
rect 409 2132 462 2137
rect 801 2132 862 2137
rect 1097 2132 1142 2137
rect 1337 2132 1358 2137
rect 1593 2132 1686 2137
rect 1801 2132 1886 2137
rect 241 2122 302 2127
rect 393 2122 526 2127
rect 649 2122 742 2127
rect 793 2122 870 2127
rect 1113 2122 1238 2127
rect 1329 2122 1382 2127
rect 1449 2122 1574 2127
rect 1953 2122 1958 2142
rect 2001 2132 2102 2137
rect 2241 2132 2550 2137
rect 2577 2127 2582 2147
rect 2801 2142 2846 2147
rect 3049 2142 3094 2147
rect 3193 2142 3222 2147
rect 3297 2147 3302 2152
rect 3297 2142 3326 2147
rect 3353 2142 3414 2147
rect 3441 2142 3614 2147
rect 3641 2142 4238 2147
rect 4233 2137 4238 2142
rect 4353 2142 4382 2147
rect 4465 2142 4502 2147
rect 4353 2137 4358 2142
rect 2601 2132 2782 2137
rect 3129 2132 3158 2137
rect 3257 2132 3422 2137
rect 3969 2132 3998 2137
rect 4233 2132 4358 2137
rect 4673 2132 4766 2137
rect 2601 2127 2606 2132
rect 2089 2122 2222 2127
rect 2577 2122 2606 2127
rect 2777 2127 2782 2132
rect 4673 2127 4678 2132
rect 2777 2122 3302 2127
rect 3593 2122 3646 2127
rect 4617 2122 4678 2127
rect 4761 2127 4766 2132
rect 4761 2122 4790 2127
rect 297 2117 398 2122
rect 649 2117 654 2122
rect 177 2112 270 2117
rect 417 2112 446 2117
rect 441 2107 446 2112
rect 505 2112 654 2117
rect 737 2117 742 2122
rect 1449 2117 1454 2122
rect 737 2112 766 2117
rect 809 2112 942 2117
rect 961 2112 1062 2117
rect 1297 2112 1358 2117
rect 1385 2112 1454 2117
rect 1569 2117 1574 2122
rect 3297 2117 3302 2122
rect 1569 2112 1718 2117
rect 2081 2112 2134 2117
rect 2201 2112 2350 2117
rect 2513 2112 2694 2117
rect 3185 2112 3278 2117
rect 3297 2112 3558 2117
rect 3721 2112 3766 2117
rect 4425 2112 4470 2117
rect 4697 2112 4758 2117
rect 505 2107 510 2112
rect 961 2107 966 2112
rect 281 2102 350 2107
rect 441 2102 510 2107
rect 561 2102 590 2107
rect 665 2102 966 2107
rect 1057 2107 1062 2112
rect 1177 2107 1262 2112
rect 1057 2102 1182 2107
rect 1257 2102 1286 2107
rect 585 2097 670 2102
rect 289 2092 350 2097
rect 945 2092 1022 2097
rect 1193 2092 1230 2097
rect 793 2087 926 2092
rect 1281 2087 1286 2102
rect 1465 2102 1590 2107
rect 1729 2102 2070 2107
rect 1465 2087 1470 2102
rect 1585 2097 1734 2102
rect 2065 2097 2070 2102
rect 2249 2102 2502 2107
rect 2585 2102 2646 2107
rect 2737 2102 2854 2107
rect 3497 2102 3550 2107
rect 3625 2102 3734 2107
rect 4617 2102 4678 2107
rect 2249 2097 2254 2102
rect 1489 2092 1566 2097
rect 2065 2092 2254 2097
rect 2273 2092 2350 2097
rect 2537 2092 2726 2097
rect 2721 2087 2726 2092
rect 2865 2092 3486 2097
rect 3561 2092 3670 2097
rect 4457 2092 4494 2097
rect 2865 2087 2870 2092
rect 3481 2087 3566 2092
rect 529 2082 566 2087
rect 585 2082 750 2087
rect 769 2082 798 2087
rect 921 2082 990 2087
rect 1001 2082 1046 2087
rect 1281 2082 1470 2087
rect 1505 2082 1662 2087
rect 1681 2082 1830 2087
rect 1849 2082 1878 2087
rect 1889 2082 1926 2087
rect 2409 2082 2686 2087
rect 2721 2082 2870 2087
rect 4073 2082 4158 2087
rect 585 2077 590 2082
rect 561 2072 590 2077
rect 745 2077 750 2082
rect 1681 2077 1686 2082
rect 745 2072 1086 2077
rect 1545 2072 1686 2077
rect 1825 2077 1830 2082
rect 3177 2077 3246 2082
rect 1825 2072 2006 2077
rect 2569 2072 2638 2077
rect 2921 2072 3134 2077
rect 3153 2072 3182 2077
rect 3241 2072 4126 2077
rect 609 2067 726 2072
rect 1705 2067 1806 2072
rect 2921 2067 2926 2072
rect 457 2062 614 2067
rect 721 2062 998 2067
rect 1105 2062 1190 2067
rect 1633 2062 1710 2067
rect 1801 2062 1886 2067
rect 2017 2062 2102 2067
rect 2177 2062 2254 2067
rect 2297 2062 2430 2067
rect 2513 2062 2590 2067
rect 2753 2062 2878 2067
rect 2897 2062 2926 2067
rect 3129 2067 3134 2072
rect 3129 2062 3230 2067
rect 4449 2062 4478 2067
rect 1025 2057 1110 2062
rect 1185 2057 1190 2062
rect 1553 2057 1638 2062
rect 1881 2057 2022 2062
rect 2177 2057 2182 2062
rect 505 2052 534 2057
rect 625 2052 886 2057
rect 1009 2052 1030 2057
rect 1185 2052 1558 2057
rect 1657 2052 1862 2057
rect 529 2047 630 2052
rect 881 2047 1014 2052
rect 1857 2047 1862 2052
rect 2113 2052 2182 2057
rect 2249 2057 2254 2062
rect 2753 2057 2758 2062
rect 2249 2052 2350 2057
rect 2113 2047 2118 2052
rect 2345 2047 2350 2052
rect 2441 2052 2502 2057
rect 2441 2047 2446 2052
rect 793 2042 862 2047
rect 1041 2042 1126 2047
rect 1569 2042 1814 2047
rect 1857 2042 2118 2047
rect 2193 2042 2238 2047
rect 2345 2042 2446 2047
rect 2497 2047 2502 2052
rect 2601 2052 2758 2057
rect 2873 2057 2878 2062
rect 2945 2057 3110 2062
rect 2873 2052 2950 2057
rect 3105 2052 3390 2057
rect 2601 2047 2606 2052
rect 3385 2047 3390 2052
rect 3489 2052 3646 2057
rect 3489 2047 3494 2052
rect 2497 2042 2606 2047
rect 2769 2042 3166 2047
rect 3385 2042 3494 2047
rect 3641 2047 3646 2052
rect 3745 2052 3774 2057
rect 4073 2052 4142 2057
rect 3745 2047 3750 2052
rect 4073 2047 4078 2052
rect 3641 2042 3750 2047
rect 3969 2042 4078 2047
rect 4137 2047 4142 2052
rect 4137 2042 4246 2047
rect 4297 2042 4382 2047
rect 649 2037 758 2042
rect 4297 2037 4302 2042
rect 289 2032 382 2037
rect 513 2032 582 2037
rect 321 2022 462 2027
rect 545 2012 574 2017
rect 593 2007 598 2037
rect 577 2002 598 2007
rect 625 2032 654 2037
rect 753 2032 782 2037
rect 801 2032 854 2037
rect 873 2032 974 2037
rect 1129 2032 1174 2037
rect 1361 2032 1446 2037
rect 1665 2032 1702 2037
rect 2257 2032 2326 2037
rect 3105 2032 3166 2037
rect 4089 2032 4302 2037
rect 4377 2037 4382 2042
rect 4377 2032 4694 2037
rect 625 2002 630 2032
rect 2257 2027 2262 2032
rect 665 2022 710 2027
rect 769 2022 830 2027
rect 769 2002 774 2022
rect 1009 2017 1014 2027
rect 1057 2022 1150 2027
rect 1377 2022 1406 2027
rect 1737 2022 1766 2027
rect 1801 2022 1838 2027
rect 2065 2022 2262 2027
rect 2321 2027 2326 2032
rect 2865 2027 3006 2032
rect 2321 2022 2870 2027
rect 3001 2022 3366 2027
rect 3513 2022 3534 2027
rect 3577 2022 3622 2027
rect 3881 2022 3990 2027
rect 4105 2022 4174 2027
rect 4225 2022 4366 2027
rect 1761 2017 1766 2022
rect 1009 2012 1126 2017
rect 1761 2012 1854 2017
rect 1929 2012 2134 2017
rect 2273 2012 2310 2017
rect 2881 2012 2990 2017
rect 3113 2012 3134 2017
rect 3185 2012 3230 2017
rect 3905 2012 3982 2017
rect 4217 2012 4326 2017
rect 2489 2007 2846 2012
rect 3281 2007 3390 2012
rect 865 2002 1006 2007
rect 1937 2002 1990 2007
rect 2089 2002 2118 2007
rect 2113 1997 2118 2002
rect 2313 2002 2494 2007
rect 2841 2002 3286 2007
rect 3385 2002 3414 2007
rect 3489 2002 3526 2007
rect 4337 2002 4654 2007
rect 4697 2002 4758 2007
rect 2313 1997 2318 2002
rect 4337 1997 4342 2002
rect 481 1992 550 1997
rect 1273 1992 1526 1997
rect 1681 1992 1718 1997
rect 1801 1992 1870 1997
rect 2113 1992 2318 1997
rect 2505 1992 2830 1997
rect 2905 1992 3134 1997
rect 3297 1992 3430 1997
rect 3569 1992 3622 1997
rect 4057 1992 4182 1997
rect 4193 1992 4214 1997
rect 3153 1987 3278 1992
rect 4193 1987 4198 1992
rect 609 1982 862 1987
rect 1129 1982 1254 1987
rect 1289 1982 1366 1987
rect 1769 1982 1846 1987
rect 1865 1982 1918 1987
rect 1937 1982 2022 1987
rect 1129 1977 1134 1982
rect 321 1972 358 1977
rect 897 1972 1086 1977
rect 1105 1972 1134 1977
rect 1249 1977 1254 1982
rect 1937 1977 1942 1982
rect 1249 1972 1358 1977
rect 1377 1972 1446 1977
rect 1457 1972 1534 1977
rect 1617 1972 1782 1977
rect 1881 1972 1942 1977
rect 2017 1977 2022 1982
rect 2361 1982 2486 1987
rect 2601 1982 3158 1987
rect 3273 1982 3486 1987
rect 3753 1982 3886 1987
rect 4145 1982 4198 1987
rect 4209 1987 4214 1992
rect 4305 1992 4342 1997
rect 4305 1987 4310 1992
rect 4209 1982 4310 1987
rect 4329 1982 4406 1987
rect 2361 1977 2366 1982
rect 2481 1977 2582 1982
rect 2017 1972 2062 1977
rect 2337 1972 2366 1977
rect 2577 1972 3310 1977
rect 3649 1972 3710 1977
rect 897 1967 902 1972
rect 529 1962 566 1967
rect 769 1962 854 1967
rect 873 1962 902 1967
rect 1081 1967 1086 1972
rect 1081 1962 1430 1967
rect 1537 1962 1566 1967
rect 1649 1962 1678 1967
rect 769 1957 774 1962
rect 97 1952 254 1957
rect 401 1952 558 1957
rect 649 1952 678 1957
rect 745 1952 774 1957
rect 849 1957 854 1962
rect 1425 1957 1542 1962
rect 1673 1957 1678 1962
rect 1753 1962 2006 1967
rect 1753 1957 1758 1962
rect 2001 1957 2006 1962
rect 2073 1962 2694 1967
rect 2801 1962 2862 1967
rect 2889 1962 3166 1967
rect 3273 1962 3302 1967
rect 3425 1962 3582 1967
rect 3601 1962 3630 1967
rect 2073 1957 2078 1962
rect 2689 1957 2806 1962
rect 3161 1957 3278 1962
rect 3425 1957 3430 1962
rect 849 1952 878 1957
rect 945 1952 1014 1957
rect 1033 1952 1078 1957
rect 1305 1952 1326 1957
rect 1337 1952 1406 1957
rect 1673 1952 1758 1957
rect 1777 1952 1894 1957
rect 1937 1952 1974 1957
rect 2001 1952 2078 1957
rect 2441 1952 2486 1957
rect 2497 1952 2542 1957
rect 2577 1952 2598 1957
rect 2617 1952 2670 1957
rect 2825 1952 2870 1957
rect 3097 1952 3142 1957
rect 3401 1952 3430 1957
rect 3577 1957 3582 1962
rect 3577 1952 3686 1957
rect 3729 1952 3878 1957
rect 4137 1952 4254 1957
rect 4377 1952 4462 1957
rect 4529 1952 4590 1957
rect 945 1947 950 1952
rect 233 1942 278 1947
rect 329 1942 390 1947
rect 169 1932 222 1937
rect 385 1927 390 1942
rect 521 1942 950 1947
rect 1009 1947 1014 1952
rect 2929 1947 2998 1952
rect 1009 1942 1334 1947
rect 521 1927 526 1942
rect 1329 1937 1334 1942
rect 1417 1942 1638 1947
rect 1881 1942 1982 1947
rect 2401 1942 2558 1947
rect 2681 1942 2814 1947
rect 2881 1942 2934 1947
rect 2993 1942 3334 1947
rect 3353 1942 3614 1947
rect 4257 1942 4526 1947
rect 4641 1942 4798 1947
rect 1417 1937 1422 1942
rect 689 1927 694 1937
rect 961 1932 1078 1937
rect 265 1922 334 1927
rect 385 1922 526 1927
rect 545 1922 894 1927
rect 913 1922 1006 1927
rect 1081 1922 1118 1927
rect 633 1912 694 1917
rect 825 1912 918 1917
rect 1065 1912 1150 1917
rect 1201 1912 1206 1937
rect 1329 1932 1422 1937
rect 1633 1937 1638 1942
rect 1793 1937 1886 1942
rect 2553 1937 2686 1942
rect 2809 1937 2886 1942
rect 3329 1937 3334 1942
rect 3673 1937 3758 1942
rect 1633 1932 1798 1937
rect 1905 1932 1998 1937
rect 2089 1932 2118 1937
rect 2321 1932 2390 1937
rect 2489 1932 2518 1937
rect 2945 1932 2982 1937
rect 3161 1932 3206 1937
rect 3329 1932 3678 1937
rect 3753 1932 3782 1937
rect 2321 1927 2326 1932
rect 2385 1927 2494 1932
rect 3777 1927 3782 1932
rect 3881 1932 3942 1937
rect 4137 1932 4182 1937
rect 4377 1932 4438 1937
rect 4465 1932 4606 1937
rect 3881 1927 3886 1932
rect 1241 1922 1310 1927
rect 1441 1922 1558 1927
rect 1849 1922 1942 1927
rect 2009 1922 2326 1927
rect 2561 1922 2606 1927
rect 2809 1922 2878 1927
rect 3057 1922 3118 1927
rect 3137 1922 3582 1927
rect 3689 1922 3718 1927
rect 3777 1922 3886 1927
rect 3985 1922 4046 1927
rect 1241 1917 1246 1922
rect 1217 1912 1246 1917
rect 1305 1917 1310 1922
rect 3577 1917 3694 1922
rect 1305 1912 1454 1917
rect 1817 1912 1854 1917
rect 2425 1912 2494 1917
rect 2537 1912 2646 1917
rect 2713 1912 2798 1917
rect 2969 1912 2998 1917
rect 3033 1912 3078 1917
rect 3097 1912 3558 1917
rect 4257 1912 4486 1917
rect 4569 1912 4662 1917
rect 4481 1907 4486 1912
rect 1257 1902 1294 1907
rect 1473 1902 1622 1907
rect 1641 1902 1734 1907
rect 2937 1902 3182 1907
rect 1313 1897 1478 1902
rect 1617 1897 1622 1902
rect 3177 1897 3182 1902
rect 3257 1902 3286 1907
rect 3409 1902 3758 1907
rect 4481 1902 4582 1907
rect 4625 1902 4678 1907
rect 3257 1897 3262 1902
rect 1185 1892 1318 1897
rect 1617 1892 1670 1897
rect 1729 1892 1758 1897
rect 1777 1892 2038 1897
rect 2057 1892 2158 1897
rect 2177 1892 2262 1897
rect 1497 1887 1598 1892
rect 1777 1887 1782 1892
rect 697 1882 1502 1887
rect 1593 1882 1782 1887
rect 2033 1887 2038 1892
rect 2177 1887 2182 1892
rect 2033 1882 2182 1887
rect 2257 1887 2262 1892
rect 2313 1892 2382 1897
rect 2529 1892 2894 1897
rect 2913 1892 3102 1897
rect 3177 1892 3262 1897
rect 3289 1892 3518 1897
rect 3777 1892 4006 1897
rect 2313 1887 2318 1892
rect 2257 1882 2318 1887
rect 2377 1887 2382 1892
rect 3777 1887 3782 1892
rect 2377 1882 2518 1887
rect 2601 1882 2630 1887
rect 3001 1882 3022 1887
rect 3041 1882 3158 1887
rect 3537 1882 3782 1887
rect 2513 1877 2606 1882
rect 2873 1877 2982 1882
rect 3041 1877 3046 1882
rect 3233 1877 3334 1882
rect 3377 1877 3542 1882
rect 4001 1877 4006 1892
rect 4025 1882 4118 1887
rect 4137 1882 4366 1887
rect 4137 1877 4142 1882
rect 1241 1872 1486 1877
rect 1545 1872 1662 1877
rect 1753 1872 1862 1877
rect 1977 1872 2038 1877
rect 2161 1872 2246 1877
rect 2329 1872 2366 1877
rect 2849 1872 2878 1877
rect 2977 1872 3046 1877
rect 3081 1872 3110 1877
rect 3209 1872 3238 1877
rect 3329 1872 3382 1877
rect 4001 1872 4142 1877
rect 4361 1877 4366 1882
rect 4361 1872 4750 1877
rect 1273 1862 1446 1867
rect 1841 1862 2102 1867
rect 2433 1862 3318 1867
rect 3393 1862 3486 1867
rect 3553 1862 4094 1867
rect 2129 1857 2246 1862
rect 3393 1857 3398 1862
rect 3481 1857 3558 1862
rect 4089 1857 4094 1862
rect 4201 1862 4278 1867
rect 4201 1857 4206 1862
rect 601 1852 670 1857
rect 601 1847 606 1852
rect 465 1842 606 1847
rect 665 1847 670 1852
rect 889 1852 1126 1857
rect 1145 1852 1174 1857
rect 1465 1852 1726 1857
rect 1745 1852 1774 1857
rect 1873 1852 2134 1857
rect 2241 1852 2374 1857
rect 2865 1852 3398 1857
rect 3417 1852 3462 1857
rect 3729 1852 3846 1857
rect 3977 1852 4006 1857
rect 4089 1852 4206 1857
rect 4281 1852 4350 1857
rect 4545 1852 4590 1857
rect 889 1847 894 1852
rect 665 1842 894 1847
rect 1121 1847 1126 1852
rect 1193 1847 1374 1852
rect 1465 1847 1470 1852
rect 1121 1842 1198 1847
rect 1369 1842 1470 1847
rect 1721 1847 1726 1852
rect 1721 1842 2414 1847
rect 2513 1842 2542 1847
rect 2569 1842 2590 1847
rect 2617 1842 2686 1847
rect 2617 1837 2622 1842
rect 121 1832 158 1837
rect 937 1832 1246 1837
rect 1265 1832 1358 1837
rect 1473 1832 2502 1837
rect 2593 1832 2622 1837
rect 2681 1837 2686 1842
rect 2705 1842 2990 1847
rect 3017 1842 3718 1847
rect 2705 1837 2710 1842
rect 3713 1837 3718 1842
rect 3857 1842 4038 1847
rect 4681 1842 4774 1847
rect 3857 1837 3862 1842
rect 4681 1837 4686 1842
rect 2681 1832 2710 1837
rect 2881 1832 2918 1837
rect 2937 1832 3358 1837
rect 3713 1832 3862 1837
rect 3921 1832 4014 1837
rect 4657 1832 4686 1837
rect 4769 1837 4774 1842
rect 4769 1832 4798 1837
rect 2497 1827 2598 1832
rect 3457 1827 3670 1832
rect 617 1822 654 1827
rect 673 1822 886 1827
rect 905 1822 1158 1827
rect 1249 1822 1334 1827
rect 1657 1822 1742 1827
rect 1857 1822 1894 1827
rect 1929 1822 2046 1827
rect 2097 1822 2230 1827
rect 2281 1822 2318 1827
rect 673 1817 678 1822
rect 337 1812 358 1817
rect 369 1812 678 1817
rect 881 1817 886 1822
rect 1353 1817 1494 1822
rect 2313 1817 2318 1822
rect 2385 1822 2414 1827
rect 2633 1822 2670 1827
rect 2777 1822 2822 1827
rect 2833 1822 2910 1827
rect 3025 1822 3158 1827
rect 3433 1822 3462 1827
rect 3665 1822 3694 1827
rect 3929 1822 3998 1827
rect 4105 1822 4150 1827
rect 4217 1822 4510 1827
rect 4529 1822 4582 1827
rect 4649 1822 4678 1827
rect 4697 1822 4750 1827
rect 2385 1817 2390 1822
rect 881 1812 1358 1817
rect 1489 1812 2206 1817
rect 2265 1812 2294 1817
rect 2313 1812 2390 1817
rect 2465 1812 2694 1817
rect 2921 1812 3078 1817
rect 3201 1812 3366 1817
rect 3385 1812 3614 1817
rect 3673 1812 3718 1817
rect 3737 1812 3902 1817
rect 4121 1812 4198 1817
rect 97 1802 222 1807
rect 289 1802 318 1807
rect 369 1797 374 1812
rect 521 1802 550 1807
rect 689 1802 1478 1807
rect 1809 1802 1966 1807
rect 2041 1802 2158 1807
rect 2633 1802 2734 1807
rect 2961 1802 3014 1807
rect 3065 1802 3150 1807
rect 241 1792 374 1797
rect 545 1797 550 1802
rect 625 1797 694 1802
rect 1553 1797 1622 1802
rect 1689 1797 1782 1802
rect 3201 1797 3206 1812
rect 3361 1807 3366 1812
rect 3737 1807 3742 1812
rect 3897 1807 4038 1812
rect 4217 1807 4222 1822
rect 4505 1812 4510 1822
rect 4505 1807 4646 1812
rect 4713 1807 4718 1817
rect 4777 1812 4814 1817
rect 3361 1802 3742 1807
rect 4033 1802 4222 1807
rect 4241 1802 4318 1807
rect 4641 1802 4670 1807
rect 4697 1802 4718 1807
rect 4241 1797 4246 1802
rect 545 1792 630 1797
rect 945 1792 1110 1797
rect 1233 1792 1286 1797
rect 1393 1792 1558 1797
rect 1617 1792 1694 1797
rect 1777 1792 1806 1797
rect 2017 1792 2094 1797
rect 2273 1792 2342 1797
rect 2449 1792 2558 1797
rect 2665 1792 2782 1797
rect 2953 1792 2982 1797
rect 3153 1792 3206 1797
rect 3217 1792 3246 1797
rect 3257 1792 3694 1797
rect 3761 1792 3878 1797
rect 3913 1792 4022 1797
rect 4089 1792 4126 1797
rect 4217 1792 4246 1797
rect 4313 1797 4318 1802
rect 4313 1792 4718 1797
rect 1825 1787 1998 1792
rect 4017 1787 4022 1792
rect 153 1782 270 1787
rect 409 1782 518 1787
rect 513 1777 518 1782
rect 649 1782 934 1787
rect 649 1777 654 1782
rect 513 1772 654 1777
rect 929 1777 934 1782
rect 993 1782 1094 1787
rect 993 1777 998 1782
rect 1089 1777 1094 1782
rect 1305 1782 1606 1787
rect 1305 1777 1310 1782
rect 1601 1777 1606 1782
rect 1705 1782 1830 1787
rect 1993 1782 2406 1787
rect 2657 1782 2822 1787
rect 3049 1782 3942 1787
rect 4017 1782 4310 1787
rect 1705 1777 1710 1782
rect 4305 1777 4310 1782
rect 4609 1782 4742 1787
rect 4609 1777 4614 1782
rect 929 1772 998 1777
rect 1049 1772 1070 1777
rect 1089 1772 1310 1777
rect 1425 1772 1582 1777
rect 1601 1772 1710 1777
rect 1809 1772 2070 1777
rect 2337 1772 2646 1777
rect 2761 1772 2934 1777
rect 2969 1772 3630 1777
rect 3737 1772 4022 1777
rect 4161 1772 4214 1777
rect 4305 1772 4614 1777
rect 4633 1772 4662 1777
rect 377 1762 494 1767
rect 785 1762 814 1767
rect 1017 1762 1054 1767
rect 1329 1762 1390 1767
rect 1505 1762 1526 1767
rect 1577 1757 1582 1772
rect 1809 1767 1814 1772
rect 2137 1767 2238 1772
rect 2641 1767 2766 1772
rect 3625 1767 3742 1772
rect 4657 1767 4662 1772
rect 4737 1772 4766 1777
rect 4737 1767 4742 1772
rect 1729 1762 1814 1767
rect 1841 1762 1918 1767
rect 2081 1762 2142 1767
rect 2233 1762 2318 1767
rect 2785 1762 2838 1767
rect 2945 1762 3062 1767
rect 3161 1762 3502 1767
rect 1729 1757 1734 1762
rect 1913 1757 2086 1762
rect 3057 1757 3166 1762
rect 3497 1757 3502 1762
rect 3761 1762 4286 1767
rect 4657 1762 4742 1767
rect 3761 1757 3766 1762
rect 673 1752 702 1757
rect 881 1752 990 1757
rect 1441 1752 1534 1757
rect 1577 1752 1734 1757
rect 1833 1752 1894 1757
rect 2153 1752 2278 1757
rect 2289 1752 2358 1757
rect 2425 1752 2446 1757
rect 2649 1752 2718 1757
rect 3185 1752 3262 1757
rect 3353 1752 3470 1757
rect 3497 1752 3766 1757
rect 3785 1752 4222 1757
rect 4465 1752 4534 1757
rect 881 1747 886 1752
rect 2745 1747 3038 1752
rect 4529 1747 4534 1752
rect 345 1742 510 1747
rect 769 1742 886 1747
rect 1089 1742 1158 1747
rect 1281 1742 1382 1747
rect 1777 1742 1846 1747
rect 1993 1742 2110 1747
rect 2553 1742 2654 1747
rect 2721 1742 2750 1747
rect 3033 1742 3350 1747
rect 3369 1742 3398 1747
rect 3881 1742 3918 1747
rect 3953 1742 3990 1747
rect 3985 1737 3990 1742
rect 4065 1742 4206 1747
rect 4225 1742 4270 1747
rect 4441 1742 4486 1747
rect 4529 1742 4606 1747
rect 4065 1737 4070 1742
rect 1305 1732 1326 1737
rect 1473 1732 1558 1737
rect 1753 1732 1782 1737
rect 1841 1732 1878 1737
rect 2169 1732 2310 1737
rect 2561 1732 3022 1737
rect 3233 1732 3390 1737
rect 3417 1732 3478 1737
rect 3625 1732 3766 1737
rect 3849 1732 3894 1737
rect 3945 1732 3966 1737
rect 3985 1732 4070 1737
rect 4169 1732 4222 1737
rect 4289 1732 4374 1737
rect 281 1722 382 1727
rect 489 1722 566 1727
rect 625 1722 678 1727
rect 961 1722 998 1727
rect 1361 1722 1398 1727
rect 1513 1722 1566 1727
rect 1841 1722 1846 1732
rect 3625 1727 3630 1732
rect 2249 1722 2286 1727
rect 2393 1722 2758 1727
rect 2889 1722 3230 1727
rect 3257 1722 3366 1727
rect 3393 1722 3502 1727
rect 3601 1722 3630 1727
rect 3761 1727 3766 1732
rect 4289 1727 4294 1732
rect 3761 1722 3894 1727
rect 4129 1722 4166 1727
rect 4201 1722 4294 1727
rect 4369 1727 4374 1732
rect 4369 1722 4446 1727
rect 4561 1722 4694 1727
rect 2753 1717 2894 1722
rect 3393 1717 3398 1722
rect 1009 1712 1118 1717
rect 1225 1712 1350 1717
rect 1545 1712 1590 1717
rect 1657 1712 1758 1717
rect 1801 1712 1878 1717
rect 2153 1712 2198 1717
rect 2217 1712 2302 1717
rect 2345 1712 2390 1717
rect 2497 1712 2734 1717
rect 2913 1712 3030 1717
rect 3233 1712 3278 1717
rect 3369 1712 3398 1717
rect 3425 1712 3494 1717
rect 3649 1712 3742 1717
rect 3801 1712 3878 1717
rect 3889 1712 3894 1722
rect 3937 1712 3966 1717
rect 4081 1712 4214 1717
rect 4233 1712 4294 1717
rect 4649 1712 4718 1717
rect 3049 1707 3150 1712
rect 3649 1707 3654 1712
rect 1097 1702 1198 1707
rect 1569 1702 1630 1707
rect 1753 1702 1910 1707
rect 2481 1702 2726 1707
rect 2761 1702 2870 1707
rect 2905 1702 3054 1707
rect 3145 1702 3222 1707
rect 3217 1697 3222 1702
rect 3289 1702 3358 1707
rect 3289 1697 3294 1702
rect 593 1692 646 1697
rect 1857 1692 1894 1697
rect 2625 1692 2742 1697
rect 2945 1692 3134 1697
rect 3217 1692 3294 1697
rect 3353 1697 3358 1702
rect 3425 1702 3454 1707
rect 3473 1702 3654 1707
rect 3737 1707 3742 1712
rect 4081 1707 4086 1712
rect 3737 1702 4086 1707
rect 4209 1707 4214 1712
rect 4209 1702 4422 1707
rect 4489 1702 4670 1707
rect 3425 1697 3430 1702
rect 3353 1692 3430 1697
rect 3497 1692 3526 1697
rect 3649 1692 3958 1697
rect 3521 1687 3654 1692
rect 1793 1682 1822 1687
rect 1849 1682 1886 1687
rect 2001 1682 2046 1687
rect 2305 1682 2462 1687
rect 2649 1682 2862 1687
rect 3673 1682 3734 1687
rect 4545 1682 4598 1687
rect 2305 1677 2310 1682
rect 1633 1672 1774 1677
rect 1873 1672 1918 1677
rect 2065 1672 2262 1677
rect 2281 1672 2310 1677
rect 2457 1677 2462 1682
rect 2881 1677 3022 1682
rect 2457 1672 2638 1677
rect 1633 1667 1638 1672
rect 1097 1662 1182 1667
rect 1097 1657 1102 1662
rect 985 1652 1102 1657
rect 1177 1657 1182 1662
rect 1537 1662 1638 1667
rect 1769 1667 1774 1672
rect 2065 1667 2070 1672
rect 1769 1662 1854 1667
rect 1537 1657 1542 1662
rect 1849 1657 1854 1662
rect 1937 1662 2070 1667
rect 1937 1657 1942 1662
rect 1177 1652 1542 1657
rect 1673 1652 1750 1657
rect 1849 1652 1942 1657
rect 2257 1657 2262 1672
rect 2633 1667 2638 1672
rect 2705 1672 2886 1677
rect 3017 1672 3102 1677
rect 3177 1672 3926 1677
rect 3977 1672 4334 1677
rect 2705 1667 2710 1672
rect 3977 1667 3982 1672
rect 2633 1662 2710 1667
rect 2729 1662 2814 1667
rect 2841 1662 3006 1667
rect 3001 1657 3006 1662
rect 3113 1662 3166 1667
rect 3113 1657 3118 1662
rect 2257 1652 2454 1657
rect 2809 1652 2918 1657
rect 3001 1652 3118 1657
rect 3161 1657 3166 1662
rect 3289 1662 3318 1667
rect 3657 1662 3734 1667
rect 3937 1662 3982 1667
rect 4329 1667 4334 1672
rect 4329 1662 4534 1667
rect 3289 1657 3294 1662
rect 3849 1657 3942 1662
rect 4057 1657 4174 1662
rect 4529 1657 4534 1662
rect 4609 1662 4870 1667
rect 4609 1657 4614 1662
rect 3161 1652 3294 1657
rect 3313 1652 3646 1657
rect 3745 1652 3854 1657
rect 3953 1652 4014 1657
rect 4033 1652 4062 1657
rect 4169 1652 4198 1657
rect 4529 1652 4614 1657
rect 1673 1647 1678 1652
rect 1649 1642 1678 1647
rect 1745 1647 1750 1652
rect 3641 1647 3750 1652
rect 1745 1642 2142 1647
rect 2265 1642 2294 1647
rect 2673 1642 2950 1647
rect 3865 1642 4150 1647
rect 4289 1642 4318 1647
rect 3401 1637 3494 1642
rect 4145 1637 4230 1642
rect 4289 1637 4294 1642
rect 385 1632 414 1637
rect 521 1632 566 1637
rect 137 1622 222 1627
rect 337 1622 358 1627
rect 385 1612 390 1632
rect 561 1612 566 1632
rect 577 1612 582 1637
rect 657 1632 742 1637
rect 1017 1632 1038 1637
rect 1113 1632 1166 1637
rect 1289 1632 1390 1637
rect 1553 1632 1750 1637
rect 1897 1632 1950 1637
rect 2177 1632 2246 1637
rect 2473 1632 2646 1637
rect 2745 1632 2790 1637
rect 2857 1632 2886 1637
rect 1289 1627 1294 1632
rect 593 1622 654 1627
rect 817 1622 918 1627
rect 977 1622 1102 1627
rect 1177 1622 1294 1627
rect 1385 1627 1390 1632
rect 2473 1627 2478 1632
rect 1385 1622 1542 1627
rect 1097 1617 1182 1622
rect 1537 1617 1542 1622
rect 1641 1622 1886 1627
rect 2097 1622 2166 1627
rect 2257 1622 2478 1627
rect 2641 1627 2646 1632
rect 2881 1627 2886 1632
rect 2953 1632 2982 1637
rect 3337 1632 3406 1637
rect 3489 1632 3614 1637
rect 3689 1632 3718 1637
rect 2953 1627 2958 1632
rect 3713 1627 3718 1632
rect 3809 1632 3870 1637
rect 3977 1632 3998 1637
rect 4049 1632 4126 1637
rect 4225 1632 4294 1637
rect 4425 1632 4502 1637
rect 4633 1632 4694 1637
rect 3809 1627 3814 1632
rect 4049 1627 4054 1632
rect 2641 1622 2766 1627
rect 2817 1622 2854 1627
rect 2881 1622 2958 1627
rect 3129 1622 3166 1627
rect 3345 1622 3374 1627
rect 3401 1622 3478 1627
rect 3713 1622 3814 1627
rect 3849 1622 4054 1627
rect 4081 1622 4206 1627
rect 4393 1622 4438 1627
rect 4561 1622 4614 1627
rect 4657 1622 4798 1627
rect 1641 1617 1646 1622
rect 1881 1617 1950 1622
rect 2097 1617 2102 1622
rect 2161 1617 2262 1622
rect 593 1612 614 1617
rect 1305 1612 1374 1617
rect 1537 1612 1646 1617
rect 1673 1612 1702 1617
rect 1945 1612 2102 1617
rect 3185 1612 3318 1617
rect 593 1602 598 1612
rect 897 1602 918 1607
rect 1033 1602 1166 1607
rect 1209 1602 1502 1607
rect 1665 1602 1686 1607
rect 281 1592 470 1597
rect 913 1592 918 1602
rect 1697 1597 1702 1612
rect 3185 1607 3190 1612
rect 1809 1602 1918 1607
rect 2121 1602 2230 1607
rect 2425 1602 2470 1607
rect 2481 1602 2518 1607
rect 2553 1602 2630 1607
rect 3121 1602 3190 1607
rect 3313 1607 3318 1612
rect 3601 1607 3606 1617
rect 3833 1612 3862 1617
rect 4153 1612 4174 1617
rect 4617 1612 4750 1617
rect 3857 1607 3862 1612
rect 3313 1602 3438 1607
rect 3577 1602 3606 1607
rect 3841 1602 3862 1607
rect 4113 1602 4150 1607
rect 4529 1602 4654 1607
rect 4529 1597 4534 1602
rect 1353 1592 1438 1597
rect 1577 1592 1678 1597
rect 1697 1592 1758 1597
rect 1833 1592 1926 1597
rect 2169 1592 2222 1597
rect 2249 1592 2278 1597
rect 2297 1592 2398 1597
rect 2441 1592 2494 1597
rect 2969 1592 3078 1597
rect 3113 1592 3142 1597
rect 2297 1587 2302 1592
rect 1137 1582 1510 1587
rect 1585 1582 1822 1587
rect 1945 1582 2022 1587
rect 2129 1582 2302 1587
rect 2393 1587 2398 1592
rect 3137 1587 3142 1592
rect 3201 1592 3302 1597
rect 3201 1587 3206 1592
rect 2393 1582 2422 1587
rect 2489 1582 2534 1587
rect 3137 1582 3206 1587
rect 3297 1587 3302 1592
rect 3401 1592 3718 1597
rect 3865 1592 4038 1597
rect 4289 1592 4534 1597
rect 4545 1592 4718 1597
rect 3401 1587 3406 1592
rect 4545 1587 4550 1592
rect 3297 1582 3406 1587
rect 3545 1582 3614 1587
rect 3705 1582 3790 1587
rect 4241 1582 4374 1587
rect 1945 1577 1950 1582
rect 1673 1572 1950 1577
rect 2017 1577 2022 1582
rect 4369 1577 4374 1582
rect 4449 1582 4550 1587
rect 4569 1582 4638 1587
rect 4449 1577 4454 1582
rect 2017 1572 2134 1577
rect 2145 1572 2198 1577
rect 2377 1572 2614 1577
rect 3425 1572 3502 1577
rect 3785 1572 3854 1577
rect 4369 1572 4454 1577
rect 4473 1572 4638 1577
rect 2217 1567 2342 1572
rect 585 1562 614 1567
rect 1265 1562 1398 1567
rect 1641 1562 2006 1567
rect 2113 1562 2222 1567
rect 2337 1562 2478 1567
rect 2577 1562 2606 1567
rect 3169 1562 3294 1567
rect 3393 1562 3542 1567
rect 617 1552 646 1557
rect 737 1552 870 1557
rect 1009 1552 1222 1557
rect 1009 1547 1014 1552
rect 521 1542 726 1547
rect 825 1542 854 1547
rect 985 1542 1014 1547
rect 1217 1547 1222 1552
rect 1265 1547 1270 1562
rect 1217 1542 1270 1547
rect 1393 1547 1398 1562
rect 2001 1557 2118 1562
rect 2473 1557 2582 1562
rect 3169 1557 3174 1562
rect 1505 1552 1590 1557
rect 1649 1552 1694 1557
rect 1761 1552 1806 1557
rect 1889 1552 1926 1557
rect 2137 1552 2326 1557
rect 2409 1552 2454 1557
rect 3145 1552 3174 1557
rect 3289 1557 3294 1562
rect 3537 1557 3542 1562
rect 3625 1562 3702 1567
rect 3761 1562 3838 1567
rect 4601 1562 4646 1567
rect 3625 1557 3630 1562
rect 3289 1552 3318 1557
rect 3361 1552 3494 1557
rect 3537 1552 3630 1557
rect 3689 1552 3782 1557
rect 4337 1552 4374 1557
rect 4529 1552 4598 1557
rect 4641 1552 4790 1557
rect 1393 1542 1486 1547
rect 1553 1542 1606 1547
rect 2057 1542 2206 1547
rect 2529 1542 2566 1547
rect 2961 1542 3006 1547
rect 3249 1542 3278 1547
rect 3409 1542 3510 1547
rect 4513 1542 4590 1547
rect 4657 1542 4678 1547
rect 721 1537 830 1542
rect 361 1532 462 1537
rect 865 1532 974 1537
rect 969 1527 974 1532
rect 1105 1532 1206 1537
rect 1617 1532 1750 1537
rect 1105 1527 1110 1532
rect 1201 1527 1422 1532
rect 1497 1527 1622 1532
rect 1745 1527 1750 1532
rect 1817 1532 2046 1537
rect 2185 1532 2382 1537
rect 2417 1532 2478 1537
rect 2585 1532 2750 1537
rect 2817 1532 2942 1537
rect 2985 1532 3222 1537
rect 3449 1532 3518 1537
rect 3737 1532 3806 1537
rect 4281 1532 4358 1537
rect 4465 1532 4486 1537
rect 4497 1532 4566 1537
rect 4585 1532 4630 1537
rect 1817 1527 1822 1532
rect 2041 1527 2190 1532
rect 89 1522 270 1527
rect 385 1507 390 1527
rect 545 1522 574 1527
rect 569 1517 574 1522
rect 737 1522 774 1527
rect 969 1522 1110 1527
rect 1417 1522 1502 1527
rect 1745 1522 1822 1527
rect 2657 1522 2702 1527
rect 2873 1522 2902 1527
rect 3073 1522 3102 1527
rect 737 1517 742 1522
rect 2209 1517 2358 1522
rect 2433 1517 2502 1522
rect 3097 1517 3102 1522
rect 3225 1522 3302 1527
rect 3425 1522 3494 1527
rect 3529 1522 3606 1527
rect 4465 1522 4470 1532
rect 4689 1527 4694 1537
rect 4649 1522 4694 1527
rect 3225 1517 3230 1522
rect 569 1512 742 1517
rect 761 1512 846 1517
rect 1225 1512 1270 1517
rect 1329 1512 1398 1517
rect 1577 1512 1686 1517
rect 1881 1512 2214 1517
rect 2353 1512 2438 1517
rect 2497 1512 2646 1517
rect 2713 1512 2806 1517
rect 2641 1507 2718 1512
rect 2801 1507 2806 1512
rect 2881 1512 2910 1517
rect 3097 1512 3230 1517
rect 3465 1512 3502 1517
rect 3585 1512 3630 1517
rect 3753 1512 3814 1517
rect 4113 1512 4134 1517
rect 4329 1512 4606 1517
rect 4689 1512 4734 1517
rect 2881 1507 2886 1512
rect 385 1502 462 1507
rect 1129 1502 1206 1507
rect 1305 1502 1334 1507
rect 1457 1502 1622 1507
rect 1665 1502 1702 1507
rect 2225 1502 2262 1507
rect 2313 1502 2342 1507
rect 2449 1502 2486 1507
rect 2801 1502 2886 1507
rect 3561 1502 3590 1507
rect 1129 1497 1134 1502
rect 1201 1497 1278 1502
rect 2337 1497 2454 1502
rect 785 1492 1134 1497
rect 1273 1492 1446 1497
rect 1441 1487 1446 1492
rect 1713 1492 2214 1497
rect 1713 1487 1718 1492
rect 1145 1482 1262 1487
rect 1441 1482 1718 1487
rect 2209 1487 2214 1492
rect 2473 1492 2502 1497
rect 2625 1492 2710 1497
rect 3833 1492 3958 1497
rect 4193 1492 4318 1497
rect 2473 1487 2478 1492
rect 3833 1487 3838 1492
rect 2209 1482 2478 1487
rect 3489 1482 3838 1487
rect 3953 1487 3958 1492
rect 4313 1487 4318 1492
rect 4417 1492 4590 1497
rect 4417 1487 4422 1492
rect 3953 1482 3982 1487
rect 4313 1482 4422 1487
rect 4481 1482 4502 1487
rect 4537 1482 4630 1487
rect 4441 1472 4470 1477
rect 3785 1467 3934 1472
rect 969 1462 1062 1467
rect 969 1457 974 1462
rect 801 1452 974 1457
rect 1057 1457 1062 1462
rect 1345 1462 2598 1467
rect 1345 1457 1350 1462
rect 1057 1452 1350 1457
rect 2593 1457 2598 1462
rect 3201 1462 3430 1467
rect 3473 1462 3494 1467
rect 3761 1462 3790 1467
rect 3929 1462 4182 1467
rect 2593 1452 2622 1457
rect 1785 1447 2094 1452
rect 3201 1447 3206 1462
rect 241 1442 358 1447
rect 241 1437 246 1442
rect 217 1432 246 1437
rect 353 1437 358 1442
rect 409 1442 502 1447
rect 409 1437 414 1442
rect 353 1432 414 1437
rect 497 1437 502 1442
rect 1577 1442 1718 1447
rect 1577 1437 1582 1442
rect 497 1432 526 1437
rect 601 1432 814 1437
rect 985 1432 1046 1437
rect 1361 1432 1582 1437
rect 1713 1437 1718 1442
rect 1761 1442 1790 1447
rect 2089 1442 2118 1447
rect 2137 1442 2206 1447
rect 2489 1442 2574 1447
rect 2601 1442 2662 1447
rect 2681 1442 2758 1447
rect 1761 1437 1766 1442
rect 1713 1432 1766 1437
rect 2113 1437 2118 1442
rect 2489 1437 2494 1442
rect 2113 1432 2310 1437
rect 2353 1432 2494 1437
rect 2569 1437 2574 1442
rect 2681 1437 2686 1442
rect 2569 1432 2686 1437
rect 2753 1437 2758 1442
rect 2849 1442 2926 1447
rect 2849 1437 2854 1442
rect 2753 1432 2854 1437
rect 2921 1437 2926 1442
rect 3073 1442 3206 1447
rect 3425 1447 3430 1462
rect 4465 1457 4470 1472
rect 4641 1472 4678 1477
rect 4641 1457 4646 1472
rect 3473 1452 3542 1457
rect 3585 1452 3670 1457
rect 3769 1452 3918 1457
rect 4465 1452 4646 1457
rect 3585 1447 3590 1452
rect 3425 1442 3454 1447
rect 3561 1442 3590 1447
rect 3665 1447 3670 1452
rect 3665 1442 3766 1447
rect 3785 1442 3822 1447
rect 4313 1442 4422 1447
rect 3073 1437 3078 1442
rect 4313 1437 4318 1442
rect 2921 1432 3078 1437
rect 3217 1432 3278 1437
rect 3329 1432 3414 1437
rect 3409 1427 3414 1432
rect 3489 1432 3654 1437
rect 3753 1432 3830 1437
rect 3977 1432 4022 1437
rect 4177 1432 4318 1437
rect 4417 1437 4422 1442
rect 4417 1432 4446 1437
rect 3489 1427 3494 1432
rect 193 1422 254 1427
rect 777 1422 878 1427
rect 1033 1422 1150 1427
rect 1593 1422 1718 1427
rect 1969 1422 2278 1427
rect 2433 1422 2470 1427
rect 2505 1422 2638 1427
rect 2865 1422 2910 1427
rect 3097 1422 3134 1427
rect 3281 1422 3374 1427
rect 3409 1422 3494 1427
rect 3577 1422 3638 1427
rect 3817 1422 3862 1427
rect 4225 1422 4278 1427
rect 4337 1422 4550 1427
rect 4673 1422 4798 1427
rect 1713 1417 1718 1422
rect 1777 1417 1974 1422
rect 193 1412 350 1417
rect 345 1407 350 1412
rect 425 1412 550 1417
rect 833 1412 886 1417
rect 1025 1412 1174 1417
rect 1417 1412 1550 1417
rect 1713 1412 1782 1417
rect 1993 1412 2022 1417
rect 2153 1412 2222 1417
rect 425 1407 430 1412
rect 2017 1407 2158 1412
rect 2217 1407 2222 1412
rect 2345 1412 2390 1417
rect 2441 1412 2742 1417
rect 3089 1412 3190 1417
rect 4473 1412 4534 1417
rect 2345 1407 2350 1412
rect 345 1402 430 1407
rect 489 1402 526 1407
rect 681 1402 734 1407
rect 953 1402 1166 1407
rect 1801 1402 1910 1407
rect 2177 1402 2198 1407
rect 2217 1402 2350 1407
rect 2465 1402 2654 1407
rect 2785 1402 2830 1407
rect 2841 1402 2886 1407
rect 3297 1402 3366 1407
rect 3713 1402 3822 1407
rect 3929 1402 4006 1407
rect 3929 1397 3934 1402
rect 449 1392 574 1397
rect 625 1392 678 1397
rect 673 1387 678 1392
rect 745 1392 790 1397
rect 1049 1392 1102 1397
rect 1137 1392 1246 1397
rect 1321 1392 1454 1397
rect 1729 1392 1758 1397
rect 1953 1392 2078 1397
rect 2097 1392 2190 1397
rect 2369 1392 2454 1397
rect 2577 1392 2614 1397
rect 2961 1392 3070 1397
rect 3481 1392 3558 1397
rect 3681 1392 3750 1397
rect 3833 1392 3934 1397
rect 4001 1397 4006 1402
rect 4081 1402 4206 1407
rect 4081 1397 4086 1402
rect 4001 1392 4086 1397
rect 4201 1397 4206 1402
rect 4201 1392 4246 1397
rect 4257 1392 4382 1397
rect 4529 1392 4598 1397
rect 745 1387 750 1392
rect 2961 1387 2966 1392
rect 233 1382 262 1387
rect 673 1382 750 1387
rect 1041 1382 1094 1387
rect 1209 1382 1254 1387
rect 2041 1382 2158 1387
rect 2409 1382 2566 1387
rect 2625 1382 2966 1387
rect 3065 1387 3070 1392
rect 3745 1387 3838 1392
rect 3065 1382 3110 1387
rect 3537 1382 3726 1387
rect 2561 1377 2630 1382
rect 3721 1377 3726 1382
rect 3857 1382 3990 1387
rect 3857 1377 3862 1382
rect 137 1372 206 1377
rect 225 1372 310 1377
rect 2209 1372 2318 1377
rect 2977 1372 3222 1377
rect 3721 1372 3862 1377
rect 3985 1377 3990 1382
rect 4097 1382 4254 1387
rect 4537 1382 4606 1387
rect 4097 1377 4102 1382
rect 3985 1372 4102 1377
rect 4569 1372 4694 1377
rect 137 1367 142 1372
rect 105 1362 142 1367
rect 201 1367 206 1372
rect 2209 1367 2214 1372
rect 201 1362 230 1367
rect 329 1362 454 1367
rect 1489 1362 1606 1367
rect 2105 1362 2214 1367
rect 2313 1367 2318 1372
rect 2313 1362 2342 1367
rect 2377 1362 2414 1367
rect 2521 1362 2798 1367
rect 225 1357 334 1362
rect 1489 1357 1494 1362
rect 409 1352 438 1357
rect 1033 1352 1190 1357
rect 1465 1352 1494 1357
rect 1601 1357 1606 1362
rect 2521 1357 2526 1362
rect 1601 1352 1958 1357
rect 2057 1352 2142 1357
rect 2441 1352 2526 1357
rect 2793 1357 2798 1362
rect 2881 1362 2958 1367
rect 2993 1362 3126 1367
rect 3137 1362 3166 1367
rect 3305 1362 3342 1367
rect 3881 1362 3918 1367
rect 4449 1362 4518 1367
rect 2881 1357 2886 1362
rect 2793 1352 2886 1357
rect 2953 1357 2958 1362
rect 4449 1357 4454 1362
rect 2953 1352 2990 1357
rect 3153 1352 3190 1357
rect 3257 1352 3286 1357
rect 3905 1352 4454 1357
rect 4513 1357 4518 1362
rect 4513 1352 4566 1357
rect 2161 1347 2398 1352
rect 2561 1347 2758 1352
rect 3905 1347 3910 1352
rect 4561 1347 4566 1352
rect 4633 1352 4718 1357
rect 4633 1347 4638 1352
rect 153 1342 182 1347
rect 209 1342 246 1347
rect 385 1342 478 1347
rect 497 1342 582 1347
rect 841 1342 862 1347
rect 1145 1342 1198 1347
rect 1481 1342 1590 1347
rect 2017 1342 2166 1347
rect 2393 1342 2422 1347
rect 2537 1342 2566 1347
rect 2753 1342 2782 1347
rect 2897 1342 2926 1347
rect 2961 1342 3006 1347
rect 3361 1342 3398 1347
rect 3441 1342 3534 1347
rect 3705 1342 3910 1347
rect 3937 1342 3974 1347
rect 4393 1342 4422 1347
rect 4417 1337 4422 1342
rect 4489 1342 4542 1347
rect 4561 1342 4638 1347
rect 4489 1337 4494 1342
rect 129 1332 262 1337
rect 1097 1332 1374 1337
rect 2049 1332 2286 1337
rect 2321 1332 2374 1337
rect 2369 1327 2374 1332
rect 2433 1332 3206 1337
rect 4417 1332 4494 1337
rect 4513 1332 4542 1337
rect 2433 1327 2438 1332
rect 681 1322 822 1327
rect 1393 1322 1470 1327
rect 2289 1322 2350 1327
rect 2369 1322 2438 1327
rect 2481 1322 2630 1327
rect 2729 1322 2942 1327
rect 3049 1322 3078 1327
rect 3329 1322 3366 1327
rect 185 1312 302 1317
rect 393 1312 446 1317
rect 505 1312 550 1317
rect 1009 1312 1078 1317
rect 1201 1312 1334 1317
rect 1345 1312 1422 1317
rect 1577 1312 1694 1317
rect 1809 1312 1846 1317
rect 2097 1312 2166 1317
rect 2601 1312 2686 1317
rect 2777 1312 2822 1317
rect 2889 1312 2950 1317
rect 3577 1312 3702 1317
rect 3793 1312 3838 1317
rect 3881 1312 3934 1317
rect 3969 1312 4022 1317
rect 4249 1312 4294 1317
rect 4465 1312 4518 1317
rect 4665 1312 4718 1317
rect 1329 1307 1334 1312
rect 97 1302 182 1307
rect 401 1302 438 1307
rect 513 1302 542 1307
rect 697 1302 718 1307
rect 1057 1302 1078 1307
rect 1329 1302 1598 1307
rect 1721 1302 1766 1307
rect 1977 1302 2118 1307
rect 2137 1302 2286 1307
rect 2473 1302 2702 1307
rect 2921 1302 2966 1307
rect 3057 1302 3102 1307
rect 3121 1302 3206 1307
rect 3273 1302 3326 1307
rect 433 1292 462 1297
rect 1081 1292 1102 1297
rect 2665 1292 2886 1297
rect 3097 1292 3182 1297
rect 2185 1287 2294 1292
rect 1833 1282 2078 1287
rect 2161 1282 2190 1287
rect 2289 1282 2318 1287
rect 2529 1282 3094 1287
rect 3697 1282 3702 1312
rect 4281 1302 4390 1307
rect 4489 1302 4510 1307
rect 1833 1277 1838 1282
rect 1809 1272 1838 1277
rect 2073 1277 2078 1282
rect 2073 1272 2150 1277
rect 2217 1272 2310 1277
rect 2337 1272 2510 1277
rect 2801 1272 2942 1277
rect 3057 1272 3086 1277
rect 3241 1272 3478 1277
rect 3505 1272 3526 1277
rect 2145 1267 2222 1272
rect 2337 1267 2342 1272
rect 2505 1267 2686 1272
rect 2937 1267 3062 1272
rect 3241 1267 3246 1272
rect 1305 1262 2062 1267
rect 2057 1257 2062 1262
rect 2241 1262 2342 1267
rect 2681 1262 2710 1267
rect 3113 1262 3246 1267
rect 2241 1257 2246 1262
rect 3113 1257 3118 1262
rect 3473 1257 3478 1272
rect 185 1252 214 1257
rect 809 1252 910 1257
rect 1057 1252 1174 1257
rect 1761 1252 1982 1257
rect 2057 1252 2246 1257
rect 2369 1252 2406 1257
rect 2425 1252 3118 1257
rect 3369 1252 3454 1257
rect 3473 1252 3566 1257
rect 3585 1252 3830 1257
rect 809 1247 814 1252
rect 177 1242 222 1247
rect 785 1242 814 1247
rect 905 1247 910 1252
rect 3369 1247 3374 1252
rect 905 1242 942 1247
rect 1073 1242 1102 1247
rect 1201 1242 1294 1247
rect 2297 1242 2366 1247
rect 2393 1242 2518 1247
rect 1097 1237 1206 1242
rect 1721 1237 1822 1242
rect 2513 1237 2518 1242
rect 2657 1242 2702 1247
rect 3257 1242 3374 1247
rect 3449 1247 3454 1252
rect 3585 1247 3590 1252
rect 3449 1242 3590 1247
rect 3825 1247 3830 1252
rect 3969 1252 4150 1257
rect 4649 1252 4718 1257
rect 3825 1242 3950 1247
rect 2657 1237 2662 1242
rect 2841 1237 2910 1242
rect 3969 1237 3974 1252
rect 337 1232 374 1237
rect 689 1232 766 1237
rect 969 1232 1070 1237
rect 1297 1232 1342 1237
rect 1697 1232 1726 1237
rect 1817 1232 2038 1237
rect 2265 1232 2318 1237
rect 2361 1232 2430 1237
rect 2441 1232 2478 1237
rect 2513 1232 2662 1237
rect 2681 1232 2846 1237
rect 2905 1232 3318 1237
rect 3313 1227 3318 1232
rect 3385 1232 3438 1237
rect 3385 1227 3390 1232
rect 289 1222 382 1227
rect 817 1222 894 1227
rect 1065 1222 1094 1227
rect 1201 1222 1334 1227
rect 1385 1222 1518 1227
rect 1385 1217 1390 1222
rect 1097 1212 1190 1217
rect 1257 1212 1390 1217
rect 1513 1217 1518 1222
rect 1561 1222 1678 1227
rect 1745 1222 1806 1227
rect 1969 1222 2006 1227
rect 2073 1222 2102 1227
rect 2233 1222 2278 1227
rect 2321 1222 2470 1227
rect 2857 1222 3030 1227
rect 3089 1222 3118 1227
rect 3313 1222 3390 1227
rect 3433 1227 3438 1232
rect 3513 1232 3558 1237
rect 3937 1232 3974 1237
rect 4145 1237 4150 1252
rect 4433 1242 4478 1247
rect 4145 1232 4174 1237
rect 4449 1232 4526 1237
rect 3513 1227 3518 1232
rect 3937 1227 3942 1232
rect 3433 1222 3518 1227
rect 3537 1222 3686 1227
rect 3721 1222 3782 1227
rect 3825 1222 3942 1227
rect 3953 1222 3998 1227
rect 4089 1222 4158 1227
rect 4257 1222 4302 1227
rect 4417 1222 4462 1227
rect 4497 1222 4534 1227
rect 4561 1222 4598 1227
rect 4609 1222 4630 1227
rect 4689 1222 4742 1227
rect 1561 1217 1566 1222
rect 1513 1212 1566 1217
rect 1673 1217 1678 1222
rect 3113 1217 3294 1222
rect 1673 1212 1822 1217
rect 1993 1212 2014 1217
rect 2385 1212 2414 1217
rect 2497 1212 2774 1217
rect 2793 1212 3054 1217
rect 1185 1207 1262 1212
rect 2497 1207 2502 1212
rect 337 1202 622 1207
rect 945 1202 1046 1207
rect 1401 1202 1550 1207
rect 1833 1202 2046 1207
rect 945 1197 950 1202
rect 89 1192 278 1197
rect 369 1192 414 1197
rect 457 1192 494 1197
rect 921 1192 950 1197
rect 1041 1197 1046 1202
rect 1313 1197 1406 1202
rect 1545 1197 1550 1202
rect 1721 1197 1838 1202
rect 2041 1197 2046 1202
rect 2113 1202 2502 1207
rect 2769 1207 2774 1212
rect 3289 1207 3294 1217
rect 3537 1207 3542 1222
rect 3825 1217 3830 1222
rect 3657 1212 3830 1217
rect 3865 1212 3974 1217
rect 4065 1212 4150 1217
rect 4193 1212 4238 1217
rect 4529 1212 4534 1222
rect 4609 1217 4614 1222
rect 4577 1212 4614 1217
rect 4625 1212 4678 1217
rect 4425 1207 4510 1212
rect 2769 1202 2870 1207
rect 2977 1202 3270 1207
rect 3289 1202 3542 1207
rect 3569 1202 3590 1207
rect 3801 1202 3878 1207
rect 4073 1202 4142 1207
rect 4225 1202 4430 1207
rect 4505 1202 4566 1207
rect 4577 1202 4582 1212
rect 4689 1202 4734 1207
rect 2113 1197 2118 1202
rect 2537 1197 2638 1202
rect 2865 1197 2982 1202
rect 1041 1192 1142 1197
rect 1185 1192 1270 1197
rect 1313 1187 1318 1197
rect 1441 1192 1526 1197
rect 1545 1192 1726 1197
rect 1929 1192 2014 1197
rect 2041 1192 2118 1197
rect 2433 1192 2494 1197
rect 2513 1192 2542 1197
rect 2633 1192 2774 1197
rect 2809 1192 2846 1197
rect 3561 1192 3694 1197
rect 3689 1187 3694 1192
rect 3809 1192 3918 1197
rect 3809 1187 3814 1192
rect 3913 1187 3918 1192
rect 3985 1192 4110 1197
rect 4145 1192 4190 1197
rect 4233 1192 4270 1197
rect 4441 1192 4558 1197
rect 4569 1192 4702 1197
rect 3985 1187 3990 1192
rect 81 1182 198 1187
rect 737 1182 1318 1187
rect 1337 1182 1446 1187
rect 1745 1182 1862 1187
rect 2305 1182 2470 1187
rect 2481 1182 3118 1187
rect 3113 1177 3118 1182
rect 3217 1182 3246 1187
rect 3689 1182 3814 1187
rect 3857 1182 3894 1187
rect 3913 1182 3990 1187
rect 4345 1182 4374 1187
rect 3217 1177 3222 1182
rect 4369 1177 4374 1182
rect 4481 1182 4598 1187
rect 4481 1177 4486 1182
rect 4593 1177 4598 1182
rect 4745 1182 4782 1187
rect 4745 1177 4750 1182
rect 873 1172 902 1177
rect 897 1167 902 1172
rect 993 1172 1046 1177
rect 1137 1172 1166 1177
rect 1369 1172 1398 1177
rect 1545 1172 1806 1177
rect 993 1167 998 1172
rect 897 1162 998 1167
rect 1161 1167 1166 1172
rect 1257 1167 1374 1172
rect 1801 1167 1806 1172
rect 1873 1172 2022 1177
rect 2193 1172 2222 1177
rect 2313 1172 2446 1177
rect 2577 1172 2646 1177
rect 2841 1172 2902 1177
rect 3113 1172 3222 1177
rect 3441 1172 3526 1177
rect 3545 1172 3566 1177
rect 4369 1172 4486 1177
rect 4505 1172 4574 1177
rect 4593 1172 4750 1177
rect 1873 1167 1878 1172
rect 2665 1167 2734 1172
rect 3441 1167 3446 1172
rect 1161 1162 1262 1167
rect 1633 1162 1766 1167
rect 1801 1162 1878 1167
rect 2417 1162 2486 1167
rect 2561 1162 2670 1167
rect 2729 1162 3094 1167
rect 3417 1162 3446 1167
rect 3521 1167 3526 1172
rect 3521 1162 3582 1167
rect 0 1152 118 1157
rect 401 1152 542 1157
rect 1017 1152 1046 1157
rect 1113 1152 1134 1157
rect 1281 1152 1318 1157
rect 1313 1147 1318 1152
rect 1409 1152 1534 1157
rect 1409 1147 1414 1152
rect 329 1142 358 1147
rect 881 1142 1038 1147
rect 1065 1142 1158 1147
rect 1177 1142 1230 1147
rect 1313 1142 1414 1147
rect 1529 1147 1534 1152
rect 1681 1152 1758 1157
rect 2225 1152 2718 1157
rect 2793 1152 2910 1157
rect 3345 1152 3542 1157
rect 3561 1152 3694 1157
rect 3849 1152 3974 1157
rect 1681 1147 1686 1152
rect 2225 1147 2230 1152
rect 1529 1142 1686 1147
rect 1705 1142 2230 1147
rect 2369 1142 2590 1147
rect 2929 1142 3150 1147
rect 3529 1142 3598 1147
rect 3961 1142 3982 1147
rect 4153 1142 4614 1147
rect 345 1132 462 1137
rect 969 1132 1086 1137
rect 2697 1132 2822 1137
rect 3169 1132 3254 1137
rect 3521 1132 3574 1137
rect 3945 1132 4102 1137
rect 4169 1132 4222 1137
rect 1913 1127 2006 1132
rect 2377 1127 2702 1132
rect 2817 1127 2822 1132
rect 625 1122 702 1127
rect 1137 1122 1182 1127
rect 1193 1122 1294 1127
rect 1889 1122 1918 1127
rect 2001 1122 2030 1127
rect 2057 1122 2102 1127
rect 2233 1122 2382 1127
rect 2817 1122 2918 1127
rect 2913 1117 2918 1122
rect 2985 1122 3022 1127
rect 3057 1122 3270 1127
rect 3465 1122 3542 1127
rect 3577 1122 3614 1127
rect 3769 1122 3886 1127
rect 4065 1122 4110 1127
rect 4177 1122 4294 1127
rect 4657 1122 4678 1127
rect 2985 1117 2990 1122
rect 3769 1117 3774 1122
rect 185 1112 358 1117
rect 1137 1112 1206 1117
rect 1233 1112 1302 1117
rect 1401 1112 1486 1117
rect 1665 1112 1726 1117
rect 1737 1112 1774 1117
rect 1913 1112 2030 1117
rect 2233 1112 2262 1117
rect 2393 1112 2470 1117
rect 2489 1112 2638 1117
rect 2713 1112 2750 1117
rect 2761 1112 2806 1117
rect 2913 1112 2990 1117
rect 3009 1112 3086 1117
rect 3225 1112 3302 1117
rect 3369 1112 3502 1117
rect 3585 1112 3630 1117
rect 3745 1112 3774 1117
rect 3881 1117 3886 1122
rect 3881 1112 3910 1117
rect 3953 1112 3990 1117
rect 4169 1112 4230 1117
rect 4625 1112 4654 1117
rect 345 1102 398 1107
rect 1169 1102 1238 1107
rect 1289 1102 1334 1107
rect 1817 1102 1846 1107
rect 2049 1102 2158 1107
rect 2177 1102 2406 1107
rect 2417 1102 2478 1107
rect 2049 1097 2054 1102
rect 1257 1092 1294 1097
rect 1441 1092 1646 1097
rect 1841 1092 2054 1097
rect 2153 1097 2158 1102
rect 2153 1092 2214 1097
rect 2401 1092 2406 1102
rect 2473 1097 2478 1102
rect 2577 1102 2606 1107
rect 3153 1102 3214 1107
rect 3481 1102 3550 1107
rect 3689 1102 3870 1107
rect 2577 1097 2582 1102
rect 3865 1097 3870 1102
rect 3953 1102 4118 1107
rect 4241 1102 4670 1107
rect 3953 1097 3958 1102
rect 2473 1092 2582 1097
rect 3025 1092 3102 1097
rect 3137 1092 3222 1097
rect 3641 1092 3686 1097
rect 3737 1092 3830 1097
rect 3865 1092 3958 1097
rect 473 1082 502 1087
rect 1233 1082 1262 1087
rect 1257 1077 1262 1082
rect 1345 1082 1454 1087
rect 2041 1082 2142 1087
rect 1345 1077 1350 1082
rect 2137 1077 2142 1082
rect 2241 1082 2382 1087
rect 2857 1082 2942 1087
rect 3521 1082 3750 1087
rect 4305 1082 4350 1087
rect 2241 1077 2246 1082
rect 2857 1077 2862 1082
rect 1257 1072 1350 1077
rect 1665 1072 1822 1077
rect 2137 1072 2246 1077
rect 2449 1072 2862 1077
rect 2937 1077 2942 1082
rect 2937 1072 3302 1077
rect 3673 1072 3774 1077
rect 1665 1067 1670 1072
rect 1641 1062 1670 1067
rect 1817 1067 1822 1072
rect 3769 1067 3774 1072
rect 3841 1072 4342 1077
rect 3841 1067 3846 1072
rect 1817 1062 2118 1067
rect 2873 1062 3014 1067
rect 3641 1062 3694 1067
rect 3769 1062 3846 1067
rect 4337 1062 4398 1067
rect 737 1052 926 1057
rect 1745 1052 1782 1057
rect 2265 1052 2374 1057
rect 2393 1052 2462 1057
rect 2585 1052 2646 1057
rect 2921 1052 3030 1057
rect 3585 1052 3678 1057
rect 4097 1052 4198 1057
rect 737 1037 742 1052
rect 273 1032 310 1037
rect 713 1032 742 1037
rect 921 1037 926 1052
rect 2265 1047 2270 1052
rect 1545 1042 1638 1047
rect 1657 1042 1702 1047
rect 1745 1042 1838 1047
rect 2105 1042 2270 1047
rect 2369 1047 2374 1052
rect 2369 1042 2438 1047
rect 2657 1042 2694 1047
rect 2809 1042 2974 1047
rect 3089 1042 3286 1047
rect 3089 1037 3094 1042
rect 921 1032 950 1037
rect 1401 1032 1470 1037
rect 1601 1032 1838 1037
rect 2281 1032 3094 1037
rect 3281 1037 3286 1042
rect 3281 1032 3366 1037
rect 3553 1032 3582 1037
rect 4289 1032 4374 1037
rect 4601 1032 4638 1037
rect 1401 1027 1406 1032
rect 249 1022 334 1027
rect 441 1022 558 1027
rect 665 1022 830 1027
rect 857 1022 926 1027
rect 1017 1022 1142 1027
rect 1185 1022 1406 1027
rect 1465 1027 1470 1032
rect 4289 1027 4294 1032
rect 1465 1022 1494 1027
rect 1561 1022 1638 1027
rect 1689 1022 1758 1027
rect 217 1012 246 1017
rect 473 1012 734 1017
rect 1017 1007 1022 1022
rect 449 1002 566 1007
rect 817 1002 846 1007
rect 993 1002 1022 1007
rect 1137 1007 1142 1022
rect 1753 1017 1758 1022
rect 1849 1022 2038 1027
rect 2441 1022 2494 1027
rect 2617 1022 2662 1027
rect 2801 1022 2846 1027
rect 2857 1022 2998 1027
rect 3129 1022 3230 1027
rect 3305 1022 3358 1027
rect 3425 1022 3462 1027
rect 3521 1022 3566 1027
rect 4057 1022 4102 1027
rect 4193 1022 4294 1027
rect 4369 1027 4374 1032
rect 4369 1022 4502 1027
rect 1849 1017 1854 1022
rect 2209 1017 2390 1022
rect 3129 1017 3134 1022
rect 1161 1012 1222 1017
rect 1465 1012 1510 1017
rect 1593 1012 1630 1017
rect 1705 1012 1734 1017
rect 1753 1012 1854 1017
rect 2185 1012 2214 1017
rect 2385 1012 2542 1017
rect 2537 1007 2542 1012
rect 2625 1012 2790 1017
rect 2625 1007 2630 1012
rect 1137 1002 1190 1007
rect 1417 1002 1566 1007
rect 2033 1002 2126 1007
rect 2241 1002 2374 1007
rect 265 992 294 997
rect 961 992 1022 997
rect 1065 992 1182 997
rect 1305 992 1326 997
rect 1481 992 1518 997
rect 1617 992 1710 997
rect 1801 992 2046 997
rect 2369 987 2374 1002
rect 2489 1002 2518 1007
rect 2537 1002 2630 1007
rect 2785 1007 2790 1012
rect 2857 1012 2886 1017
rect 3105 1012 3134 1017
rect 3225 1017 3230 1022
rect 4609 1017 4614 1027
rect 3225 1012 3334 1017
rect 3545 1012 4014 1017
rect 4129 1012 4174 1017
rect 4305 1012 4358 1017
rect 4473 1012 4750 1017
rect 2857 1007 2862 1012
rect 2785 1002 2862 1007
rect 2945 1002 3278 1007
rect 4193 1002 4286 1007
rect 4561 1002 4590 1007
rect 2489 987 2494 1002
rect 3481 997 3566 1002
rect 4193 997 4198 1002
rect 2889 992 2918 997
rect 3113 992 3238 997
rect 3457 992 3486 997
rect 3561 992 3638 997
rect 3841 992 3870 997
rect 4009 992 4198 997
rect 4281 997 4286 1002
rect 4281 992 4374 997
rect 4465 992 4486 997
rect 4633 992 4662 997
rect 2913 987 3118 992
rect 929 982 974 987
rect 1009 982 1054 987
rect 1161 982 1206 987
rect 1745 982 1782 987
rect 2185 982 2350 987
rect 2369 982 2494 987
rect 2649 982 2702 987
rect 2721 982 2878 987
rect 2873 977 2878 982
rect 3137 982 3206 987
rect 3433 982 3550 987
rect 4009 982 4038 987
rect 4169 982 4278 987
rect 4609 982 4646 987
rect 3137 977 3142 982
rect 969 972 1542 977
rect 1713 972 1742 977
rect 2873 972 3142 977
rect 3161 972 3190 977
rect 3201 967 3206 982
rect 3257 972 3358 977
rect 3401 972 3446 977
rect 3713 972 3742 977
rect 3993 972 4022 977
rect 3257 967 3262 972
rect 1017 962 1078 967
rect 1193 962 1270 967
rect 1721 962 1822 967
rect 2513 962 2630 967
rect 3201 962 3262 967
rect 3353 967 3358 972
rect 3353 962 3630 967
rect 4057 962 4150 967
rect 2513 957 2518 962
rect 633 952 774 957
rect 793 952 1006 957
rect 233 942 318 947
rect 417 942 518 947
rect 593 942 654 947
rect 729 942 758 947
rect 777 942 854 947
rect 1001 937 1006 952
rect 1145 952 1382 957
rect 1545 952 1654 957
rect 2137 952 2254 957
rect 2273 952 2470 957
rect 2489 952 2518 957
rect 2625 957 2630 962
rect 4057 957 4062 962
rect 2625 952 2790 957
rect 3817 952 4062 957
rect 4145 957 4150 962
rect 4145 952 4206 957
rect 1145 937 1150 952
rect 1169 942 1238 947
rect 1369 942 1462 947
rect 1561 942 1638 947
rect 1889 942 1942 947
rect 2025 942 2126 947
rect 2273 937 2278 952
rect 2465 937 2470 952
rect 2529 942 2646 947
rect 2881 942 3038 947
rect 3145 942 3174 947
rect 3265 942 3350 947
rect 3393 942 3430 947
rect 3465 942 3526 947
rect 3809 942 3974 947
rect 4041 942 4078 947
rect 4385 942 4494 947
rect 65 927 70 937
rect 209 932 270 937
rect 1001 932 1150 937
rect 1233 932 1262 937
rect 1593 932 1614 937
rect 1625 932 1694 937
rect 1785 932 1830 937
rect 305 927 398 932
rect 1433 927 1534 932
rect 65 922 198 927
rect 281 922 310 927
rect 393 922 422 927
rect 625 922 670 927
rect 1273 922 1438 927
rect 1529 922 1806 927
rect 193 917 286 922
rect 1825 917 1830 932
rect 2145 932 2278 937
rect 2329 932 2406 937
rect 2465 932 2742 937
rect 2145 927 2150 932
rect 2329 927 2334 932
rect 1889 922 2150 927
rect 2273 922 2334 927
rect 2401 927 2406 932
rect 2737 927 2742 932
rect 2793 932 2862 937
rect 3753 932 3782 937
rect 3857 932 4150 937
rect 2793 927 2798 932
rect 2857 927 2950 932
rect 3097 927 3214 932
rect 2401 922 2438 927
rect 2449 922 2478 927
rect 2577 922 2718 927
rect 2737 922 2798 927
rect 2945 922 3102 927
rect 3209 922 3238 927
rect 3249 922 3294 927
rect 3425 922 3446 927
rect 3713 922 4086 927
rect 4585 922 4710 927
rect 2473 917 2582 922
rect 321 912 374 917
rect 633 912 678 917
rect 1185 912 1262 917
rect 1257 907 1262 912
rect 1369 912 1518 917
rect 1609 912 1662 917
rect 1785 912 1830 917
rect 1873 912 1958 917
rect 2121 912 2230 917
rect 2345 912 2390 917
rect 2601 912 2934 917
rect 3081 912 3126 917
rect 3137 912 3174 917
rect 3337 912 3390 917
rect 3713 912 3718 922
rect 4081 917 4086 922
rect 3817 912 3846 917
rect 3857 912 3894 917
rect 4081 912 4134 917
rect 4353 912 4398 917
rect 4457 912 4486 917
rect 4617 912 4646 917
rect 4689 912 4734 917
rect 1369 907 1374 912
rect 257 902 334 907
rect 657 902 774 907
rect 953 902 990 907
rect 1065 902 1102 907
rect 1121 902 1182 907
rect 1257 902 1374 907
rect 1465 902 1894 907
rect 1889 897 1894 902
rect 1953 902 2014 907
rect 2369 902 2630 907
rect 3001 902 3702 907
rect 1953 897 1958 902
rect 2769 897 2902 902
rect 3697 897 3702 902
rect 3777 902 3846 907
rect 3929 902 3982 907
rect 4473 902 4598 907
rect 3777 897 3782 902
rect 281 892 398 897
rect 641 892 670 897
rect 1889 892 1958 897
rect 2089 892 2182 897
rect 2425 892 2454 897
rect 2537 892 2606 897
rect 2617 892 2774 897
rect 2897 892 2990 897
rect 3105 892 3134 897
rect 3361 892 3390 897
rect 3697 892 3782 897
rect 3801 892 3878 897
rect 4393 892 4422 897
rect 1177 887 1246 892
rect 2089 887 2094 892
rect 1 882 246 887
rect 241 877 246 882
rect 377 882 406 887
rect 505 882 550 887
rect 761 882 990 887
rect 1073 882 1182 887
rect 1241 882 1830 887
rect 1977 882 2094 887
rect 2177 887 2182 892
rect 2449 887 2542 892
rect 2985 887 3110 892
rect 4417 887 4422 892
rect 4537 892 4566 897
rect 4537 887 4542 892
rect 2177 882 2414 887
rect 377 877 382 882
rect 2409 877 2414 882
rect 2785 882 2886 887
rect 3329 882 3422 887
rect 4249 882 4318 887
rect 4417 882 4542 887
rect 241 872 382 877
rect 1193 872 1230 877
rect 2105 872 2166 877
rect 2409 872 2566 877
rect 2561 867 2566 872
rect 2785 867 2790 882
rect 3057 872 3086 877
rect 961 862 1038 867
rect 1817 862 1838 867
rect 2025 862 2094 867
rect 961 857 966 862
rect 777 852 886 857
rect 937 852 966 857
rect 1033 857 1038 862
rect 2089 857 2094 862
rect 2177 862 2238 867
rect 2313 862 2390 867
rect 2561 862 2790 867
rect 3081 867 3086 872
rect 3145 872 3382 877
rect 3145 867 3150 872
rect 3081 862 3150 867
rect 3473 862 3638 867
rect 2177 857 2182 862
rect 2313 857 2318 862
rect 1033 852 1062 857
rect 1097 852 1254 857
rect 1497 852 1686 857
rect 2089 852 2182 857
rect 2289 852 2318 857
rect 2385 857 2390 862
rect 2385 852 2542 857
rect 2809 852 2990 857
rect 3361 852 3430 857
rect 889 842 1086 847
rect 1081 837 1086 842
rect 1265 842 1486 847
rect 1777 842 1814 847
rect 1857 842 2070 847
rect 2233 842 2374 847
rect 1265 837 1270 842
rect 1481 837 1558 842
rect 1641 837 1758 842
rect 1857 837 1862 842
rect 737 832 1062 837
rect 1081 832 1270 837
rect 1553 832 1646 837
rect 1753 832 1862 837
rect 2065 837 2070 842
rect 2809 837 2814 852
rect 2065 832 2470 837
rect 2593 832 2686 837
rect 2785 832 2814 837
rect 2985 837 2990 852
rect 3473 847 3478 862
rect 3633 857 3638 862
rect 4009 862 4102 867
rect 4009 857 4014 862
rect 3633 852 4014 857
rect 4097 857 4102 862
rect 4097 852 4478 857
rect 3281 842 3478 847
rect 3497 842 3526 847
rect 3553 842 3582 847
rect 3281 837 3286 842
rect 2985 832 3094 837
rect 3129 832 3286 837
rect 3297 832 3326 837
rect 3497 832 3622 837
rect 4025 832 4086 837
rect 4665 832 4694 837
rect 2593 827 2598 832
rect 313 822 358 827
rect 809 822 886 827
rect 1489 822 1518 827
rect 1657 822 1734 827
rect 1761 822 1862 827
rect 2017 822 2054 827
rect 2209 822 2302 827
rect 2377 822 2454 827
rect 2569 822 2598 827
rect 2681 827 2686 832
rect 3321 827 3502 832
rect 2681 822 2710 827
rect 2793 822 2838 827
rect 2889 822 2982 827
rect 3121 822 3158 827
rect 3529 822 3606 827
rect 3633 822 3670 827
rect 3761 822 3854 827
rect 3873 822 3974 827
rect 3993 822 4038 827
rect 4281 822 4334 827
rect 4417 822 4462 827
rect 4625 822 4670 827
rect 4697 822 4742 827
rect 905 817 1126 822
rect 2977 817 3110 822
rect 3873 817 3878 822
rect 473 812 550 817
rect 697 812 774 817
rect 769 807 774 812
rect 881 812 910 817
rect 1121 812 1982 817
rect 2353 812 2390 817
rect 2465 812 2846 817
rect 2897 812 2926 817
rect 3105 812 3878 817
rect 3969 817 3974 822
rect 3969 812 4174 817
rect 4273 812 4406 817
rect 4473 812 4518 817
rect 4529 812 4574 817
rect 4601 812 4718 817
rect 881 807 886 812
rect 2193 807 2334 812
rect 2385 807 2470 812
rect 4401 807 4478 812
rect 4513 807 4518 812
rect 417 802 446 807
rect 769 802 886 807
rect 905 802 1110 807
rect 1617 802 1670 807
rect 1745 802 1766 807
rect 2041 802 2070 807
rect 2169 802 2198 807
rect 2329 802 2366 807
rect 2497 802 3102 807
rect 3537 802 4070 807
rect 4513 802 4638 807
rect 4673 802 4718 807
rect 3121 797 3302 802
rect 3385 797 3518 802
rect 393 792 502 797
rect 673 792 750 797
rect 985 792 1086 797
rect 1393 792 1510 797
rect 1569 792 1598 797
rect 1729 792 1806 797
rect 1833 792 1974 797
rect 1993 792 2054 797
rect 2113 792 2950 797
rect 3065 792 3126 797
rect 3297 792 3390 797
rect 3513 792 3614 797
rect 3905 792 4198 797
rect 4385 792 4414 797
rect 4449 792 4518 797
rect 4609 792 4630 797
rect 1833 787 1838 792
rect 1537 782 1694 787
rect 1809 782 1838 787
rect 1969 787 1974 792
rect 2945 787 3070 792
rect 3729 787 3806 792
rect 4193 787 4198 792
rect 1969 782 2254 787
rect 2369 782 2398 787
rect 2609 782 2702 787
rect 2825 782 2926 787
rect 3089 782 3286 787
rect 3401 782 3502 787
rect 3561 782 3734 787
rect 3801 782 3942 787
rect 4193 782 4302 787
rect 2473 777 2590 782
rect 3937 777 4062 782
rect 337 772 366 777
rect 617 772 686 777
rect 1241 772 1270 777
rect 1657 772 1798 777
rect 1793 767 1798 772
rect 1857 772 2094 777
rect 2129 772 2158 777
rect 2265 772 2478 777
rect 2585 772 2846 777
rect 2961 772 3222 777
rect 3521 772 3558 777
rect 3745 772 3830 777
rect 4057 772 4254 777
rect 4377 772 4454 777
rect 1857 767 1862 772
rect 2153 767 2270 772
rect 4449 767 4454 772
rect 4521 772 4550 777
rect 4521 767 4526 772
rect 337 762 358 767
rect 729 762 798 767
rect 1793 762 1862 767
rect 1977 762 2022 767
rect 2305 762 2422 767
rect 2489 762 2942 767
rect 3009 762 3118 767
rect 3153 762 3206 767
rect 3249 762 3334 767
rect 3401 762 3534 767
rect 3841 762 4126 767
rect 4281 762 4310 767
rect 4369 762 4430 767
rect 4449 762 4526 767
rect 729 757 734 762
rect 673 752 734 757
rect 793 757 798 762
rect 4121 757 4286 762
rect 793 752 878 757
rect 1001 752 1142 757
rect 1233 752 1630 757
rect 1881 752 2006 757
rect 2089 752 2190 757
rect 2265 752 2766 757
rect 2897 752 2982 757
rect 3033 752 3110 757
rect 3193 752 3230 757
rect 3241 752 3366 757
rect 3393 752 3470 757
rect 3529 752 3686 757
rect 3761 752 3830 757
rect 1001 747 1006 752
rect 89 742 478 747
rect 553 742 662 747
rect 745 742 782 747
rect 969 742 1006 747
rect 1137 747 1142 752
rect 2785 747 2878 752
rect 3825 747 3830 752
rect 3961 752 4102 757
rect 4337 752 4374 757
rect 4633 752 4686 757
rect 3961 747 3966 752
rect 1137 742 1166 747
rect 1305 742 1326 747
rect 1561 742 1750 747
rect 1793 742 1870 747
rect 233 732 270 737
rect 1081 732 1102 737
rect 1193 732 1270 737
rect 1193 727 1198 732
rect 89 722 126 727
rect 641 722 798 727
rect 897 722 926 727
rect 1017 722 1198 727
rect 1265 727 1270 732
rect 1393 732 1462 737
rect 1633 732 1678 737
rect 1393 727 1398 732
rect 1265 722 1398 727
rect 1457 727 1462 732
rect 1865 727 1870 742
rect 2009 742 2078 747
rect 2009 727 2014 742
rect 2073 737 2078 742
rect 2137 742 2318 747
rect 2729 742 2790 747
rect 2873 742 3182 747
rect 2137 737 2142 742
rect 2313 737 2734 742
rect 3177 737 3182 742
rect 3241 742 3414 747
rect 3481 742 3574 747
rect 3713 742 3782 747
rect 3825 742 3966 747
rect 3985 742 4030 747
rect 4145 742 4262 747
rect 4289 742 4406 747
rect 4593 742 4710 747
rect 3241 737 3246 742
rect 2073 732 2142 737
rect 2161 732 2190 737
rect 1457 722 1486 727
rect 1865 722 2014 727
rect 2185 727 2190 732
rect 2265 732 2294 737
rect 2753 732 2790 737
rect 2849 732 3006 737
rect 3017 732 3062 737
rect 3177 732 3246 737
rect 3265 732 3342 737
rect 3721 732 3766 737
rect 2265 727 2270 732
rect 3473 727 3566 732
rect 4025 727 4030 737
rect 4169 732 4326 737
rect 4697 732 4742 737
rect 2185 722 2270 727
rect 2289 722 2406 727
rect 2425 722 2486 727
rect 2601 722 2710 727
rect 2817 722 3038 727
rect 3449 722 3478 727
rect 3561 722 3622 727
rect 3713 722 3814 727
rect 3833 722 3950 727
rect 4025 722 4086 727
rect 4121 722 4238 727
rect 4433 722 4494 727
rect 753 712 878 717
rect 897 707 902 722
rect 3257 717 3350 722
rect 3833 717 3838 722
rect 969 712 998 717
rect 1025 712 1134 717
rect 1209 712 1326 717
rect 1409 712 1454 717
rect 1577 712 1654 717
rect 1713 712 1838 717
rect 2033 712 2054 717
rect 2377 712 2422 717
rect 2529 712 2566 717
rect 2601 712 2950 717
rect 2945 707 2950 712
rect 3073 712 3262 717
rect 3345 712 3838 717
rect 3945 717 3950 722
rect 3945 712 3974 717
rect 3993 712 4038 717
rect 4073 712 4174 717
rect 4561 712 4598 717
rect 4665 712 4694 717
rect 3073 707 3078 712
rect 785 702 902 707
rect 913 702 998 707
rect 1097 702 1566 707
rect 1561 697 1566 702
rect 1633 702 1702 707
rect 2201 702 2262 707
rect 2505 702 2542 707
rect 2745 702 2926 707
rect 2945 702 3078 707
rect 3273 702 3334 707
rect 3425 702 3518 707
rect 3553 702 3606 707
rect 3737 702 3766 707
rect 3849 702 3950 707
rect 4041 702 4070 707
rect 4177 702 4230 707
rect 4577 702 4630 707
rect 4641 702 4670 707
rect 1633 697 1638 702
rect 3761 697 3854 702
rect 1209 692 1318 697
rect 1561 692 1638 697
rect 1657 692 1806 697
rect 2305 692 2374 697
rect 2769 692 2846 697
rect 3377 692 3414 697
rect 3409 687 3414 692
rect 3537 692 3734 697
rect 4129 692 4158 697
rect 3537 687 3542 692
rect 4153 687 4158 692
rect 4233 692 4262 697
rect 4489 692 4550 697
rect 4233 687 4238 692
rect 1129 682 1254 687
rect 1777 682 1806 687
rect 2097 682 2294 687
rect 2385 682 2566 687
rect 3137 682 3182 687
rect 3297 682 3326 687
rect 3409 682 3542 687
rect 3561 682 3598 687
rect 3617 682 3814 687
rect 2289 677 2390 682
rect 1129 672 1238 677
rect 1409 672 1502 677
rect 1761 672 1782 677
rect 2057 672 2118 677
rect 2953 672 3126 677
rect 1409 667 1414 672
rect 3121 667 3126 672
rect 3193 672 3286 677
rect 3193 667 3198 672
rect 1161 662 1414 667
rect 2137 662 2238 667
rect 2257 662 2534 667
rect 2585 662 2934 667
rect 3121 662 3198 667
rect 3281 667 3286 672
rect 3617 667 3622 682
rect 3809 677 3814 682
rect 3961 682 4110 687
rect 4153 682 4238 687
rect 4545 687 4550 692
rect 4617 692 4654 697
rect 4617 687 4622 692
rect 4545 682 4622 687
rect 4641 682 4726 687
rect 3961 677 3966 682
rect 3633 672 3662 677
rect 3761 672 3790 677
rect 3809 672 3966 677
rect 3657 667 3766 672
rect 3281 662 3622 667
rect 2001 657 2142 662
rect 2233 657 2238 662
rect 2585 657 2590 662
rect 825 652 870 657
rect 1417 652 1462 657
rect 1521 652 1734 657
rect 1753 652 1798 657
rect 1977 652 2006 657
rect 2233 652 2366 657
rect 2401 652 2470 657
rect 2561 652 2590 657
rect 2929 657 2934 662
rect 2929 652 3014 657
rect 3665 652 3710 657
rect 4065 652 4230 657
rect 4249 652 4278 657
rect 4297 652 4390 657
rect 4409 652 4622 657
rect 1521 647 1526 652
rect 345 642 406 647
rect 1097 642 1118 647
rect 1297 642 1526 647
rect 1729 647 1734 652
rect 2465 647 2566 652
rect 4065 647 4070 652
rect 1729 642 1766 647
rect 1897 642 2238 647
rect 2321 642 2446 647
rect 2761 642 2838 647
rect 4041 642 4070 647
rect 4225 647 4230 652
rect 4297 647 4302 652
rect 4225 642 4302 647
rect 4385 647 4390 652
rect 4385 642 4414 647
rect 4473 642 4574 647
rect 1761 637 1878 642
rect 2761 637 2766 642
rect 337 632 406 637
rect 1321 632 1606 637
rect 1873 632 2766 637
rect 2833 637 2838 642
rect 2833 632 2862 637
rect 2889 632 3246 637
rect 3537 632 3558 637
rect 3913 632 4014 637
rect 4137 632 4182 637
rect 4193 632 4374 637
rect 3913 627 3918 632
rect 361 622 390 627
rect 1233 622 1294 627
rect 1409 622 1478 627
rect 1513 622 1590 627
rect 1601 622 2070 627
rect 2177 622 2230 627
rect 2241 622 2318 627
rect 2401 622 2438 627
rect 2449 617 2454 627
rect 2777 622 2902 627
rect 3289 622 3326 627
rect 3369 622 3430 627
rect 3521 622 3582 627
rect 3889 622 3918 627
rect 4009 627 4014 632
rect 4193 627 4198 632
rect 4369 627 4374 632
rect 4449 632 4478 637
rect 4553 632 4590 637
rect 4665 632 4702 637
rect 4449 627 4454 632
rect 4009 622 4198 627
rect 4289 622 4334 627
rect 4369 622 4454 627
rect 4545 622 4606 627
rect 4689 622 4734 627
rect 137 612 174 617
rect 609 612 646 617
rect 809 612 894 617
rect 1193 612 1262 617
rect 2145 612 2198 617
rect 2265 612 2454 617
rect 2513 612 2614 617
rect 2793 612 2830 617
rect 2913 612 2966 617
rect 3017 612 3206 617
rect 3305 612 3334 617
rect 3457 612 3486 617
rect 3593 612 3742 617
rect 3777 612 3918 617
rect 4089 612 4118 617
rect 4217 612 4246 617
rect 1321 607 1790 612
rect 1913 607 2126 612
rect 2513 607 2518 612
rect 3017 607 3022 612
rect 593 602 742 607
rect 1169 602 1326 607
rect 1785 602 1918 607
rect 2121 602 2518 607
rect 2681 602 2782 607
rect 2777 597 2782 602
rect 2841 602 2870 607
rect 2993 602 3022 607
rect 3201 607 3206 612
rect 3481 607 3598 612
rect 4113 607 4222 612
rect 3201 602 3350 607
rect 3945 602 3998 607
rect 4353 602 4526 607
rect 4601 602 4630 607
rect 2841 597 2846 602
rect 4353 597 4358 602
rect 297 592 342 597
rect 569 592 678 597
rect 761 592 1150 597
rect 1345 592 1534 597
rect 1577 592 1774 597
rect 1929 592 2262 597
rect 2305 592 2358 597
rect 2409 592 2510 597
rect 2705 592 2734 597
rect 2777 592 2846 597
rect 2929 592 3094 597
rect 3129 592 3222 597
rect 3497 592 3558 597
rect 3857 592 3910 597
rect 3969 592 4022 597
rect 4153 592 4358 597
rect 4521 597 4526 602
rect 4521 592 4870 597
rect 761 587 766 592
rect 193 582 278 587
rect 641 582 766 587
rect 1145 587 1150 592
rect 1145 582 1334 587
rect 193 577 198 582
rect 169 572 198 577
rect 273 577 278 582
rect 1329 577 1334 582
rect 1457 582 2454 587
rect 2865 582 2894 587
rect 2993 582 3150 587
rect 3177 582 3302 587
rect 3729 582 3846 587
rect 1457 577 1462 582
rect 2889 577 2998 582
rect 3841 577 3846 582
rect 3953 582 4054 587
rect 4425 582 4534 587
rect 3953 577 3958 582
rect 273 572 518 577
rect 657 572 1022 577
rect 1329 572 1462 577
rect 1481 572 1734 577
rect 1865 572 2110 577
rect 2233 572 2390 577
rect 2417 572 2446 577
rect 2825 572 2870 577
rect 3113 572 3142 577
rect 3169 572 3206 577
rect 3513 572 3550 577
rect 3841 572 3958 577
rect 3977 572 4070 577
rect 4233 572 4414 577
rect 4553 572 4582 577
rect 2865 567 2870 572
rect 3017 567 3118 572
rect 4409 567 4494 572
rect 4553 567 4558 572
rect 201 562 246 567
rect 521 562 694 567
rect 833 562 886 567
rect 689 557 838 562
rect 881 557 886 562
rect 1033 562 1134 567
rect 1593 562 1790 567
rect 1953 562 2006 567
rect 2321 562 2686 567
rect 2865 562 3022 567
rect 4489 562 4558 567
rect 1033 557 1038 562
rect 2137 557 2270 562
rect 289 552 334 557
rect 881 552 1038 557
rect 1241 552 1318 557
rect 1433 552 1502 557
rect 1689 552 1718 557
rect 1801 552 1886 557
rect 2113 552 2142 557
rect 2265 552 2310 557
rect 2417 552 2446 557
rect 2673 552 2710 557
rect 2809 552 2846 557
rect 1713 547 1806 552
rect 2305 547 2422 552
rect 2841 547 2846 552
rect 3041 552 3070 557
rect 3673 552 3870 557
rect 4281 552 4342 557
rect 4385 552 4470 557
rect 3041 547 3046 552
rect 3673 547 3678 552
rect 241 542 326 547
rect 361 542 470 547
rect 713 542 806 547
rect 1089 542 1126 547
rect 1169 542 1262 547
rect 1385 542 1462 547
rect 1641 542 1686 547
rect 2017 542 2070 547
rect 2161 542 2254 547
rect 2625 542 2702 547
rect 2801 542 2822 547
rect 2841 542 3046 547
rect 3153 542 3238 547
rect 3417 542 3462 547
rect 3569 542 3598 547
rect 3649 542 3678 547
rect 3865 547 3870 552
rect 3865 542 3958 547
rect 4145 542 4358 547
rect 4377 542 4430 547
rect 3233 537 3238 542
rect 4353 537 4358 542
rect 233 532 278 537
rect 753 532 1038 537
rect 1073 532 1238 537
rect 1481 532 1590 537
rect 1617 532 1790 537
rect 2209 532 2318 537
rect 1481 527 1486 532
rect 473 522 534 527
rect 601 522 710 527
rect 801 522 830 527
rect 1121 522 1150 527
rect 1257 522 1342 527
rect 1433 522 1486 527
rect 1585 527 1590 532
rect 2313 527 2318 532
rect 2385 532 2414 537
rect 3105 532 3150 537
rect 3233 532 3302 537
rect 3481 532 3518 537
rect 3649 532 3670 537
rect 4017 532 4238 537
rect 4353 532 4566 537
rect 2385 527 2390 532
rect 1585 522 1614 527
rect 1945 522 2094 527
rect 2313 522 2390 527
rect 3113 522 3158 527
rect 3153 517 3158 522
rect 3265 522 3406 527
rect 3673 522 3854 527
rect 4417 522 4446 527
rect 3265 517 3270 522
rect 4441 517 4446 522
rect 4569 522 4670 527
rect 4569 517 4574 522
rect 177 512 262 517
rect 329 512 398 517
rect 585 512 814 517
rect 873 512 902 517
rect 1321 512 1366 517
rect 1377 512 1406 517
rect 1497 512 1526 517
rect 1569 512 1718 517
rect 1777 512 1830 517
rect 1849 512 2030 517
rect 2105 512 2294 517
rect 2633 512 2798 517
rect 2841 512 2862 517
rect 3057 512 3134 517
rect 3153 512 3270 517
rect 3289 512 3334 517
rect 3625 512 3670 517
rect 3817 512 3870 517
rect 4025 512 4054 517
rect 1401 507 1502 512
rect 1713 507 1718 512
rect 2025 507 2110 512
rect 105 502 198 507
rect 649 502 694 507
rect 817 502 1206 507
rect 1345 502 1374 507
rect 1713 502 1910 507
rect 1945 502 2006 507
rect 2769 502 2774 512
rect 4049 507 4054 512
rect 4153 512 4206 517
rect 4441 512 4574 517
rect 4609 512 4638 517
rect 4673 512 4718 517
rect 4153 507 4158 512
rect 3545 502 3710 507
rect 3705 497 3710 502
rect 3777 502 3806 507
rect 3857 502 3902 507
rect 4049 502 4158 507
rect 4369 502 4406 507
rect 3777 497 3782 502
rect 121 492 150 497
rect 681 492 702 497
rect 889 492 918 497
rect 913 487 918 492
rect 1017 492 1046 497
rect 1409 492 1438 497
rect 1017 487 1022 492
rect 1433 487 1438 492
rect 1825 492 1878 497
rect 1825 487 1830 492
rect 641 482 678 487
rect 913 482 1022 487
rect 1057 482 1086 487
rect 1081 477 1086 482
rect 1153 482 1182 487
rect 1433 482 1830 487
rect 1873 487 1878 492
rect 2017 492 2182 497
rect 2017 487 2022 492
rect 1873 482 2022 487
rect 2177 487 2182 492
rect 2257 492 2286 497
rect 3569 492 3654 497
rect 3705 492 3782 497
rect 4401 497 4406 502
rect 4593 502 4622 507
rect 4593 497 4598 502
rect 4401 492 4598 497
rect 2257 487 2262 492
rect 2177 482 2262 487
rect 3377 482 3534 487
rect 1153 477 1158 482
rect 1081 472 1158 477
rect 1889 462 2158 467
rect 1889 457 1894 462
rect 801 452 886 457
rect 1545 452 1590 457
rect 1697 452 1894 457
rect 2153 457 2158 462
rect 2513 462 3182 467
rect 2153 452 2182 457
rect 2201 452 2358 457
rect 2377 452 2406 457
rect 801 447 806 452
rect 321 442 390 447
rect 689 442 758 447
rect 777 442 806 447
rect 881 447 886 452
rect 2201 447 2206 452
rect 881 442 1278 447
rect 1425 442 1526 447
rect 1561 442 1622 447
rect 1905 442 2062 447
rect 2097 442 2206 447
rect 2353 447 2358 452
rect 2513 447 2518 462
rect 2353 442 2518 447
rect 3177 447 3182 462
rect 3177 442 3342 447
rect 4425 442 4550 447
rect 689 437 694 442
rect 185 432 254 437
rect 665 432 694 437
rect 753 437 758 442
rect 1425 437 1430 442
rect 753 432 870 437
rect 1001 432 1070 437
rect 1401 432 1430 437
rect 1521 437 1526 442
rect 4425 437 4430 442
rect 1521 432 1598 437
rect 1609 432 1654 437
rect 1961 432 2102 437
rect 2129 432 2262 437
rect 2529 432 2798 437
rect 2921 432 3030 437
rect 3129 432 3166 437
rect 3401 432 3454 437
rect 3577 432 3598 437
rect 4201 432 4334 437
rect 4401 432 4430 437
rect 4545 437 4550 442
rect 4545 432 4574 437
rect 529 422 622 427
rect 649 422 798 427
rect 1209 422 1406 427
rect 1569 422 1638 427
rect 1649 422 1950 427
rect 1969 422 2046 427
rect 2145 422 2350 427
rect 2401 422 2510 427
rect 2937 422 2982 427
rect 2401 417 2406 422
rect 769 407 774 417
rect 1001 412 1094 417
rect 1185 412 1286 417
rect 1417 412 1662 417
rect 1897 412 1926 417
rect 2049 412 2142 417
rect 2329 412 2406 417
rect 2505 417 2510 422
rect 2505 412 2574 417
rect 2761 412 2838 417
rect 2913 412 2934 417
rect 1305 407 1398 412
rect 1681 407 1806 412
rect 2177 407 2286 412
rect 3025 407 3030 432
rect 3097 422 3142 427
rect 3273 422 3414 427
rect 3441 422 3486 427
rect 3569 422 3614 427
rect 3897 422 3942 427
rect 4201 417 4206 432
rect 3049 412 3118 417
rect 3561 412 3590 417
rect 3657 412 3718 417
rect 3737 412 3854 417
rect 4113 412 4206 417
rect 4329 417 4334 432
rect 4329 412 4558 417
rect 385 402 414 407
rect 689 402 734 407
rect 769 402 846 407
rect 1281 402 1310 407
rect 1393 402 1414 407
rect 1545 402 1686 407
rect 1801 402 2078 407
rect 2153 402 2182 407
rect 2281 402 2310 407
rect 1281 397 1286 402
rect 1409 397 1550 402
rect 2073 397 2158 402
rect 2305 397 2310 402
rect 2417 402 2614 407
rect 2737 402 2782 407
rect 3025 402 3262 407
rect 2417 397 2422 402
rect 3257 397 3262 402
rect 3337 402 3366 407
rect 3721 402 3766 407
rect 4217 402 4318 407
rect 3337 397 3342 402
rect 137 392 182 397
rect 769 392 830 397
rect 905 392 1286 397
rect 1305 392 1382 397
rect 1569 392 1710 397
rect 1721 392 1790 397
rect 1921 392 1990 397
rect 2001 392 2054 397
rect 2193 392 2286 397
rect 2305 392 2422 397
rect 2441 392 2678 397
rect 2897 392 2950 397
rect 3049 392 3086 397
rect 3257 392 3342 397
rect 3385 392 3542 397
rect 3681 392 3782 397
rect 3873 392 4030 397
rect 4273 392 4302 397
rect 4313 392 4358 397
rect 4425 392 4462 397
rect 3385 387 3390 392
rect 433 382 622 387
rect 801 382 950 387
rect 1401 382 1630 387
rect 1705 382 1870 387
rect 2049 382 2102 387
rect 2201 382 2238 387
rect 3361 382 3390 387
rect 3537 387 3542 392
rect 3873 387 3878 392
rect 3537 382 3878 387
rect 4025 387 4030 392
rect 4025 382 4054 387
rect 4233 382 4310 387
rect 4321 382 4598 387
rect 433 367 438 382
rect 353 362 438 367
rect 617 367 622 382
rect 4321 377 4326 382
rect 641 372 758 377
rect 753 367 758 372
rect 889 372 1342 377
rect 1353 372 1446 377
rect 2177 372 2222 377
rect 2641 372 2702 377
rect 2921 372 3094 377
rect 3713 372 3750 377
rect 3897 372 4006 377
rect 4105 372 4198 377
rect 4281 372 4326 377
rect 4337 372 4574 377
rect 889 367 894 372
rect 1465 367 1598 372
rect 2921 367 2926 372
rect 617 362 654 367
rect 753 362 894 367
rect 1017 362 1046 367
rect 1369 362 1422 367
rect 1433 362 1470 367
rect 1593 362 1694 367
rect 1777 362 2030 367
rect 2169 362 2214 367
rect 2537 362 2622 367
rect 1777 357 1782 362
rect 257 352 374 357
rect 481 352 662 357
rect 913 352 1198 357
rect 1193 347 1198 352
rect 1273 352 1390 357
rect 1481 352 1646 357
rect 1657 352 1782 357
rect 2025 357 2030 362
rect 2537 357 2542 362
rect 2025 352 2230 357
rect 2513 352 2542 357
rect 2617 357 2622 362
rect 2721 362 2878 367
rect 2897 362 2926 367
rect 3089 367 3094 372
rect 3769 367 3902 372
rect 4001 367 4006 372
rect 3089 362 3190 367
rect 3265 362 3774 367
rect 4001 362 4494 367
rect 4513 362 4550 367
rect 2721 357 2726 362
rect 2617 352 2726 357
rect 2873 357 2878 362
rect 2977 357 3070 362
rect 2873 352 2982 357
rect 3065 352 3102 357
rect 3673 352 3710 357
rect 3777 352 3990 357
rect 4217 352 4310 357
rect 4393 352 4542 357
rect 4553 352 4622 357
rect 1273 347 1278 352
rect 3209 347 3350 352
rect 3777 347 3782 352
rect 3985 347 4222 352
rect 4305 347 4398 352
rect 321 342 350 347
rect 593 342 710 347
rect 985 342 1038 347
rect 1193 342 1278 347
rect 1345 342 1406 347
rect 1513 342 1542 347
rect 1585 342 1662 347
rect 1793 342 2014 347
rect 2281 342 2334 347
rect 2497 342 2606 347
rect 2673 342 2702 347
rect 2769 342 2846 347
rect 2865 342 2918 347
rect 2993 342 3030 347
rect 3041 342 3214 347
rect 3345 342 3782 347
rect 3793 342 3830 347
rect 3849 342 3894 347
rect 4241 342 4286 347
rect 4417 342 4558 347
rect 4625 342 4710 347
rect 2161 337 2246 342
rect 2601 337 2678 342
rect 2769 337 2774 342
rect 81 332 142 337
rect 529 332 574 337
rect 633 332 734 337
rect 977 332 1110 337
rect 1297 332 1398 337
rect 1561 332 1654 337
rect 1665 332 1686 337
rect 1681 327 1686 332
rect 1985 332 2110 337
rect 2137 332 2166 337
rect 2241 332 2310 337
rect 2745 332 2774 337
rect 2841 337 2846 342
rect 3041 337 3046 342
rect 2841 332 3046 337
rect 3073 332 3334 337
rect 3457 332 3582 337
rect 3649 332 3894 337
rect 3945 332 4006 337
rect 4041 332 4174 337
rect 1985 327 1990 332
rect 4041 327 4046 332
rect 233 322 310 327
rect 345 322 382 327
rect 657 322 782 327
rect 1537 322 1614 327
rect 1657 322 1686 327
rect 1873 322 1990 327
rect 2169 322 2230 327
rect 2633 322 2662 327
rect 2721 322 2934 327
rect 3081 322 3478 327
rect 3721 322 3806 327
rect 3865 322 4046 327
rect 4169 327 4174 332
rect 4241 327 4246 342
rect 4625 337 4630 342
rect 4361 332 4630 337
rect 4649 327 4758 332
rect 4169 322 4270 327
rect 4409 322 4494 327
rect 4569 322 4654 327
rect 4753 322 4782 327
rect 785 312 1046 317
rect 1097 312 1158 317
rect 1417 312 1518 317
rect 1601 312 1654 317
rect 1705 312 1806 317
rect 1825 312 1854 317
rect 1969 312 2038 317
rect 2441 312 2486 317
rect 2577 312 2670 317
rect 2681 312 2710 317
rect 1041 307 1046 312
rect 1417 307 1422 312
rect 737 302 798 307
rect 1041 302 1214 307
rect 1233 302 1358 307
rect 1377 302 1422 307
rect 1513 307 1518 312
rect 1705 307 1710 312
rect 1513 302 1710 307
rect 1801 307 1806 312
rect 2705 307 2710 312
rect 2801 312 2830 317
rect 2905 312 2950 317
rect 3113 312 3254 317
rect 3265 312 3310 317
rect 3457 312 3502 317
rect 3569 312 3974 317
rect 3993 312 4030 317
rect 4049 312 4406 317
rect 4433 312 4438 322
rect 4537 312 4582 317
rect 4689 312 4734 317
rect 2801 307 2806 312
rect 3249 307 3254 312
rect 1801 302 1982 307
rect 2057 302 2150 307
rect 1233 297 1238 302
rect 1177 292 1238 297
rect 1353 297 1358 302
rect 2057 297 2062 302
rect 1353 292 1878 297
rect 1993 292 2062 297
rect 2145 297 2150 302
rect 2249 302 2422 307
rect 2473 302 2678 307
rect 2705 302 2806 307
rect 3145 302 3230 307
rect 3249 302 3366 307
rect 3617 302 3894 307
rect 4017 302 4342 307
rect 2249 297 2254 302
rect 2145 292 2254 297
rect 2417 297 2422 302
rect 3889 297 4022 302
rect 4337 297 4342 302
rect 4441 302 4494 307
rect 4441 297 4446 302
rect 2417 292 2446 297
rect 2585 292 2646 297
rect 3105 292 3326 297
rect 3697 292 3870 297
rect 4337 292 4446 297
rect 4489 297 4494 302
rect 4585 302 4638 307
rect 4585 297 4590 302
rect 4489 292 4590 297
rect 4609 292 4662 297
rect 1873 287 1998 292
rect 2441 287 2590 292
rect 953 282 1158 287
rect 2273 282 2398 287
rect 2609 282 2630 287
rect 2697 282 2990 287
rect 3089 282 3342 287
rect 3385 282 3598 287
rect 3633 282 3790 287
rect 3833 282 3878 287
rect 3953 282 4070 287
rect 953 277 958 282
rect 1153 277 1510 282
rect 1569 277 1854 282
rect 2057 277 2278 282
rect 2393 277 2398 282
rect 2697 277 2702 282
rect 849 272 958 277
rect 1505 272 1574 277
rect 1849 272 2062 277
rect 2393 272 2494 277
rect 2569 272 2702 277
rect 2985 277 2990 282
rect 3385 277 3390 282
rect 2985 272 3078 277
rect 3361 272 3390 277
rect 3593 277 3598 282
rect 3953 277 3958 282
rect 3593 272 3662 277
rect 3809 272 3838 277
rect 3929 272 3958 277
rect 4065 277 4070 282
rect 4065 272 4094 277
rect 4137 272 4318 277
rect 3073 267 3078 272
rect 3145 267 3366 272
rect 3657 267 3814 272
rect 4137 267 4142 272
rect 969 262 1494 267
rect 1585 262 1838 267
rect 2073 262 2382 267
rect 2473 262 2806 267
rect 3073 262 3150 267
rect 3409 262 3574 267
rect 3969 262 4142 267
rect 4313 267 4318 272
rect 4313 262 4342 267
rect 1489 257 1590 262
rect 1833 257 2078 262
rect 2377 257 2478 262
rect 3409 257 3414 262
rect 3569 257 3638 262
rect 705 252 830 257
rect 1777 252 1814 257
rect 2497 252 2974 257
rect 3169 252 3238 257
rect 3345 252 3414 257
rect 3633 252 3958 257
rect 4057 252 4254 257
rect 705 247 710 252
rect 681 242 710 247
rect 825 247 830 252
rect 1025 247 1470 252
rect 1609 247 1710 252
rect 2097 247 2230 252
rect 3169 247 3174 252
rect 825 242 1030 247
rect 1465 242 1614 247
rect 1705 242 2102 247
rect 2225 242 2574 247
rect 2593 242 2766 247
rect 2777 242 2798 247
rect 2961 242 3174 247
rect 3233 247 3238 252
rect 3953 247 4062 252
rect 4369 247 4374 257
rect 3233 242 3454 247
rect 3497 242 3566 247
rect 4265 242 4518 247
rect 4681 242 4758 247
rect 2825 237 2926 242
rect 4153 237 4270 242
rect 4681 237 4686 242
rect 473 232 654 237
rect 721 232 822 237
rect 1041 232 1374 237
rect 1385 232 1454 237
rect 1625 232 1694 237
rect 2113 232 2214 237
rect 2537 232 2782 237
rect 2801 232 2830 237
rect 2921 232 3006 237
rect 3185 232 3214 237
rect 3337 232 3398 237
rect 3553 232 3598 237
rect 3617 232 4158 237
rect 4337 232 4582 237
rect 4641 232 4686 237
rect 4753 237 4758 242
rect 4753 232 4798 237
rect 1473 227 1606 232
rect 1713 227 2094 232
rect 3209 227 3342 232
rect 3617 227 3622 232
rect 217 222 254 227
rect 593 222 750 227
rect 833 222 1478 227
rect 1601 222 1718 227
rect 2089 222 2526 227
rect 2593 222 2758 227
rect 2857 222 2910 227
rect 3105 222 3150 227
rect 3361 222 3422 227
rect 3449 222 3622 227
rect 4177 222 4390 227
rect 4409 222 4446 227
rect 4697 222 4742 227
rect 2521 217 2598 222
rect 4177 217 4182 222
rect 4385 217 4390 222
rect 169 212 206 217
rect 201 207 206 212
rect 265 212 326 217
rect 1057 212 1182 217
rect 1233 212 1614 217
rect 1633 212 1678 217
rect 1737 212 2238 217
rect 2617 212 2702 217
rect 2761 212 2838 217
rect 2889 212 2958 217
rect 2977 212 3086 217
rect 3233 212 3318 217
rect 3385 212 3446 217
rect 3785 212 3814 217
rect 3833 212 4070 217
rect 4089 212 4182 217
rect 4201 212 4366 217
rect 4385 212 4622 217
rect 265 207 270 212
rect 2337 207 2430 212
rect 2977 207 2982 212
rect 201 202 270 207
rect 1369 202 1558 207
rect 1649 202 2030 207
rect 2025 197 2030 202
rect 2121 202 2150 207
rect 2161 202 2342 207
rect 2425 202 2662 207
rect 2897 202 2982 207
rect 3081 207 3086 212
rect 3561 207 3638 212
rect 3833 207 3838 212
rect 3081 202 3158 207
rect 3273 202 3326 207
rect 3401 202 3566 207
rect 3633 202 3838 207
rect 4065 207 4070 212
rect 4065 202 4358 207
rect 2121 197 2126 202
rect 321 192 414 197
rect 537 192 662 197
rect 697 192 750 197
rect 809 192 942 197
rect 1017 192 1118 197
rect 1177 192 1974 197
rect 2025 192 2126 197
rect 2209 192 2278 197
rect 2353 192 2446 197
rect 2625 192 2726 197
rect 2753 192 2814 197
rect 2937 192 3078 197
rect 3193 192 3254 197
rect 3305 192 3358 197
rect 3577 192 3622 197
rect 3753 192 3782 197
rect 633 182 790 187
rect 513 177 614 182
rect 809 177 814 192
rect 489 172 518 177
rect 609 172 814 177
rect 937 177 942 192
rect 2481 187 2606 192
rect 3777 187 3782 192
rect 3953 192 4102 197
rect 3953 187 3958 192
rect 1201 182 1574 187
rect 1585 182 1646 187
rect 1689 182 1790 187
rect 1865 182 1918 187
rect 2185 182 2486 187
rect 2601 182 2686 187
rect 2825 182 2910 187
rect 2905 177 2910 182
rect 3033 182 3286 187
rect 3345 182 3478 187
rect 3777 182 3958 187
rect 4097 187 4102 192
rect 4177 192 4206 197
rect 4313 192 4334 197
rect 4177 187 4182 192
rect 4097 182 4182 187
rect 4353 187 4358 202
rect 4601 202 4678 207
rect 4601 187 4606 202
rect 4353 182 4606 187
rect 3033 177 3038 182
rect 937 172 1502 177
rect 1945 172 2006 177
rect 2481 172 2518 177
rect 2529 172 2710 177
rect 2905 172 3038 177
rect 3057 172 3126 177
rect 3201 172 3262 177
rect 2353 167 2486 172
rect 433 162 494 167
rect 553 162 1286 167
rect 1281 157 1286 162
rect 1393 162 1422 167
rect 1465 162 1550 167
rect 1641 162 1894 167
rect 1913 162 2030 167
rect 2065 162 2358 167
rect 2497 162 2566 167
rect 2841 162 2886 167
rect 1393 157 1398 162
rect 1641 157 1646 162
rect 481 152 510 157
rect 617 152 670 157
rect 721 152 1206 157
rect 1281 152 1398 157
rect 1617 152 1646 157
rect 1889 157 1894 162
rect 1889 152 2062 157
rect 2353 152 2606 157
rect 3457 152 3574 157
rect 3833 152 4502 157
rect 4585 152 4702 157
rect 505 147 622 152
rect 2057 147 2198 152
rect 401 142 438 147
rect 641 142 694 147
rect 705 142 758 147
rect 801 142 870 147
rect 1129 142 1222 147
rect 1417 142 1446 147
rect 1441 137 1446 142
rect 1561 142 1910 147
rect 1985 142 2038 147
rect 1561 137 1566 142
rect 2193 137 2198 147
rect 2353 137 2358 152
rect 4497 147 4502 152
rect 2417 142 2470 147
rect 2561 142 2622 147
rect 2673 142 2734 147
rect 2937 142 2998 147
rect 3121 142 3270 147
rect 3313 142 3350 147
rect 3489 142 3526 147
rect 3617 142 3902 147
rect 4497 142 4622 147
rect 529 132 598 137
rect 993 132 1030 137
rect 1305 132 1366 137
rect 1441 132 1566 137
rect 1601 132 1662 137
rect 1729 132 1758 137
rect 1841 132 1942 137
rect 2137 132 2174 137
rect 2193 132 2358 137
rect 681 122 766 127
rect 2617 122 2654 127
rect 593 112 742 117
rect 1945 112 2014 117
rect 2377 112 2446 117
rect 2681 112 2806 117
rect 2849 112 2894 117
rect 2977 112 3022 117
rect 3169 112 3214 117
rect 3249 112 3294 117
rect 4281 112 4326 117
rect 4417 112 4462 117
rect 4601 112 4646 117
rect 761 102 1934 107
rect 2025 102 2646 107
rect 1929 97 2030 102
rect 2385 87 2454 92
rect 1993 82 2390 87
rect 2449 82 2478 87
rect 753 72 1982 77
rect 2401 72 2430 77
rect 1977 67 2406 72
rect 1281 52 2790 57
rect 1065 32 1270 37
rect 1265 27 1270 32
rect 2801 32 3030 37
rect 2801 27 2806 32
rect 1265 22 2806 27
use top_level_VIA1  top_level_VIA1_0
timestamp 1680363874
transform 1 0 24 0 1 4717
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_1
timestamp 1680363874
transform 1 0 4851 0 1 4717
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_2
timestamp 1680363874
transform 1 0 48 0 1 4693
box -10 -10 10 10
use M3_M2  M3_M2_0
timestamp 1680363874
transform 1 0 2004 0 1 4685
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1680363874
transform 1 0 2316 0 1 4685
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_3
timestamp 1680363874
transform 1 0 4827 0 1 4693
box -10 -10 10 10
use top_level_VIA0  top_level_VIA0_0
timestamp 1680363874
transform 1 0 24 0 1 4670
box -10 -3 10 3
use M2_M1  M2_M1_0
timestamp 1680363874
transform 1 0 68 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1680363874
transform 1 0 140 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1680363874
transform 1 0 164 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_60
timestamp 1680363874
transform 1 0 164 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1680363874
transform 1 0 252 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1680363874
transform 1 0 284 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1680363874
transform 1 0 204 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_41
timestamp 1680363874
transform 1 0 252 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1680363874
transform 1 0 204 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1680363874
transform 1 0 292 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1680363874
transform 1 0 308 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1680363874
transform 1 0 316 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1680363874
transform 1 0 404 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1680363874
transform 1 0 356 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1680363874
transform 1 0 404 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1680363874
transform 1 0 436 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1680363874
transform 1 0 356 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1680363874
transform 1 0 460 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_4
timestamp 1680363874
transform 1 0 476 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1680363874
transform 1 0 492 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1680363874
transform 1 0 548 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1680363874
transform 1 0 588 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1680363874
transform 1 0 508 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1680363874
transform 1 0 532 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1680363874
transform 1 0 588 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1680363874
transform 1 0 508 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1680363874
transform 1 0 532 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1680363874
transform 1 0 596 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1680363874
transform 1 0 508 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1680363874
transform 1 0 620 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1680363874
transform 1 0 652 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1680363874
transform 1 0 668 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1680363874
transform 1 0 692 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1680363874
transform 1 0 748 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1680363874
transform 1 0 668 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1680363874
transform 1 0 660 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1680363874
transform 1 0 692 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1680363874
transform 1 0 764 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1680363874
transform 1 0 828 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1680363874
transform 1 0 780 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1680363874
transform 1 0 780 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1680363874
transform 1 0 828 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1680363874
transform 1 0 876 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1680363874
transform 1 0 908 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1680363874
transform 1 0 924 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1680363874
transform 1 0 900 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1680363874
transform 1 0 916 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1680363874
transform 1 0 924 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1680363874
transform 1 0 916 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1680363874
transform 1 0 956 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1680363874
transform 1 0 940 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1680363874
transform 1 0 1004 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1680363874
transform 1 0 940 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1680363874
transform 1 0 956 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_68
timestamp 1680363874
transform 1 0 1004 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1680363874
transform 1 0 1060 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_5
timestamp 1680363874
transform 1 0 1108 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_17
timestamp 1680363874
transform 1 0 1092 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1680363874
transform 1 0 1108 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1680363874
transform 1 0 1116 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1680363874
transform 1 0 1132 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1680363874
transform 1 0 1148 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1680363874
transform 1 0 1100 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1680363874
transform 1 0 1116 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1680363874
transform 1 0 1124 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1680363874
transform 1 0 1140 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1680363874
transform 1 0 1156 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1680363874
transform 1 0 1100 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1680363874
transform 1 0 1116 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1680363874
transform 1 0 1140 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1680363874
transform 1 0 1172 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1680363874
transform 1 0 1188 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1680363874
transform 1 0 1212 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1680363874
transform 1 0 1268 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1680363874
transform 1 0 1188 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1680363874
transform 1 0 1268 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1680363874
transform 1 0 1220 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1680363874
transform 1 0 1308 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1680363874
transform 1 0 1316 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1680363874
transform 1 0 1316 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_24
timestamp 1680363874
transform 1 0 1388 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1680363874
transform 1 0 1388 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_102
timestamp 1680363874
transform 1 0 1436 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1680363874
transform 1 0 1436 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_25
timestamp 1680363874
transform 1 0 1508 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1680363874
transform 1 0 1484 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1680363874
transform 1 0 1484 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1680363874
transform 1 0 1564 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1680363874
transform 1 0 1476 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1680363874
transform 1 0 1508 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_26
timestamp 1680363874
transform 1 0 1596 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1680363874
transform 1 0 1620 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1680363874
transform 1 0 1612 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1680363874
transform 1 0 1676 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1680363874
transform 1 0 1652 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1680363874
transform 1 0 1652 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1680363874
transform 1 0 1748 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1680363874
transform 1 0 1748 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_106
timestamp 1680363874
transform 1 0 1756 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_16
timestamp 1680363874
transform 1 0 1780 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1680363874
transform 1 0 1820 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_30
timestamp 1680363874
transform 1 0 1780 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1680363874
transform 1 0 1788 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1680363874
transform 1 0 1820 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_53
timestamp 1680363874
transform 1 0 1796 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_107
timestamp 1680363874
transform 1 0 1868 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1680363874
transform 1 0 1868 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_33
timestamp 1680363874
transform 1 0 1884 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_2
timestamp 1680363874
transform 1 0 1940 0 1 4645
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1680363874
transform 1 0 1948 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1680363874
transform 1 0 1988 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_34
timestamp 1680363874
transform 1 0 1948 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1680363874
transform 1 0 1988 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1680363874
transform 1 0 1972 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1680363874
transform 1 0 1988 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1680363874
transform 1 0 1956 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1680363874
transform 1 0 1988 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_36
timestamp 1680363874
transform 1 0 2020 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1680363874
transform 1 0 2060 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1680363874
transform 1 0 2100 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1680363874
transform 1 0 2100 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_38
timestamp 1680363874
transform 1 0 2164 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1680363874
transform 1 0 2220 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1680363874
transform 1 0 2140 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1680363874
transform 1 0 2140 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1680363874
transform 1 0 2252 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1680363874
transform 1 0 2292 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1680363874
transform 1 0 2252 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1680363874
transform 1 0 2260 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1680363874
transform 1 0 2292 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1680363874
transform 1 0 2244 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1680363874
transform 1 0 2340 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_100
timestamp 1680363874
transform 1 0 2340 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1680363874
transform 1 0 2388 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1680363874
transform 1 0 2428 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1680363874
transform 1 0 2388 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1680363874
transform 1 0 2396 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1680363874
transform 1 0 2428 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1680363874
transform 1 0 2380 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1680363874
transform 1 0 2476 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1680363874
transform 1 0 2428 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1680363874
transform 1 0 2476 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1680363874
transform 1 0 2492 0 1 4645
box -3 -3 3 3
use M2_M1  M2_M1_46
timestamp 1680363874
transform 1 0 2556 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1680363874
transform 1 0 2588 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1680363874
transform 1 0 2508 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1680363874
transform 1 0 2548 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1680363874
transform 1 0 2588 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1680363874
transform 1 0 2508 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1680363874
transform 1 0 2660 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1680363874
transform 1 0 2700 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1680363874
transform 1 0 2660 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1680363874
transform 1 0 2692 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1680363874
transform 1 0 2700 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1680363874
transform 1 0 2612 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1680363874
transform 1 0 2700 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_83
timestamp 1680363874
transform 1 0 2612 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1680363874
transform 1 0 2660 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_51
timestamp 1680363874
transform 1 0 2716 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_26
timestamp 1680363874
transform 1 0 2804 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1680363874
transform 1 0 2844 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1680363874
transform 1 0 2804 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1680363874
transform 1 0 2844 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1680363874
transform 1 0 2828 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1680363874
transform 1 0 2844 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_85
timestamp 1680363874
transform 1 0 2828 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_54
timestamp 1680363874
transform 1 0 2892 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1680363874
transform 1 0 2948 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1680363874
transform 1 0 2972 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_86
timestamp 1680363874
transform 1 0 2972 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1680363874
transform 1 0 3044 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_56
timestamp 1680363874
transform 1 0 3100 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1680363874
transform 1 0 3156 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1680363874
transform 1 0 3180 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_88
timestamp 1680363874
transform 1 0 3180 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_58
timestamp 1680363874
transform 1 0 3276 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1680363874
transform 1 0 3332 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1680363874
transform 1 0 3252 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_101
timestamp 1680363874
transform 1 0 3252 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1680363874
transform 1 0 3396 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1680363874
transform 1 0 3452 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1680363874
transform 1 0 3372 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1680363874
transform 1 0 3372 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_62
timestamp 1680363874
transform 1 0 3476 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1680363874
transform 1 0 3532 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1680363874
transform 1 0 3556 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1680363874
transform 1 0 3556 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_64
timestamp 1680363874
transform 1 0 3572 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1680363874
transform 1 0 3580 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1680363874
transform 1 0 3652 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1680363874
transform 1 0 3684 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1680363874
transform 1 0 3652 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1680363874
transform 1 0 3676 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1680363874
transform 1 0 3676 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1680363874
transform 1 0 3692 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1680363874
transform 1 0 3692 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1680363874
transform 1 0 3764 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1680363874
transform 1 0 3788 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_67
timestamp 1680363874
transform 1 0 3764 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1680363874
transform 1 0 3788 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1680363874
transform 1 0 3708 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1680363874
transform 1 0 3788 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1680363874
transform 1 0 3932 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1680363874
transform 1 0 3956 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_68
timestamp 1680363874
transform 1 0 3828 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1680363874
transform 1 0 3884 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1680363874
transform 1 0 3924 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1680363874
transform 1 0 3956 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1680363874
transform 1 0 3908 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_90
timestamp 1680363874
transform 1 0 3828 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_129
timestamp 1680363874
transform 1 0 4004 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1680363874
transform 1 0 3932 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1680363874
transform 1 0 4052 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1680363874
transform 1 0 4108 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1680363874
transform 1 0 4028 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_9
timestamp 1680363874
transform 1 0 4196 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1680363874
transform 1 0 4196 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1680363874
transform 1 0 4236 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_74
timestamp 1680363874
transform 1 0 4196 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1680363874
transform 1 0 4228 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1680363874
transform 1 0 4236 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1680363874
transform 1 0 4148 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1680363874
transform 1 0 4212 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_132
timestamp 1680363874
transform 1 0 4252 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_10
timestamp 1680363874
transform 1 0 4308 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1680363874
transform 1 0 4308 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1680363874
transform 1 0 4364 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1680363874
transform 1 0 4284 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1680363874
transform 1 0 4364 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_79
timestamp 1680363874
transform 1 0 4388 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1680363874
transform 1 0 4444 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1680363874
transform 1 0 4468 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1680363874
transform 1 0 4492 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_34
timestamp 1680363874
transform 1 0 4564 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_82
timestamp 1680363874
transform 1 0 4564 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1680363874
transform 1 0 4588 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1680363874
transform 1 0 4612 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_35
timestamp 1680363874
transform 1 0 4644 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1680363874
transform 1 0 4756 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_84
timestamp 1680363874
transform 1 0 4756 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1680363874
transform 1 0 4780 0 1 4605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_1
timestamp 1680363874
transform 1 0 4851 0 1 4670
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_2
timestamp 1680363874
transform 1 0 48 0 1 4570
box -10 -3 10 3
use M3_M2  M3_M2_106
timestamp 1680363874
transform 1 0 68 0 1 4575
box -3 -3 3 3
use FILL  FILL_0
timestamp 1680363874
transform 1 0 72 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1680363874
transform -1 0 176 0 1 4570
box -8 -3 104 105
use FILL  FILL_1
timestamp 1680363874
transform 1 0 176 0 1 4570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1680363874
transform 1 0 184 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1680363874
transform 1 0 192 0 1 4570
box -8 -3 104 105
use FILL  FILL_10
timestamp 1680363874
transform 1 0 288 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1680363874
transform 1 0 296 0 1 4570
box -9 -3 26 105
use FILL  FILL_11
timestamp 1680363874
transform 1 0 312 0 1 4570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1680363874
transform 1 0 320 0 1 4570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1680363874
transform 1 0 328 0 1 4570
box -8 -3 16 105
use FILL  FILL_24
timestamp 1680363874
transform 1 0 336 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1680363874
transform 1 0 344 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_3
timestamp 1680363874
transform 1 0 440 0 1 4570
box -9 -3 26 105
use FILL  FILL_25
timestamp 1680363874
transform 1 0 456 0 1 4570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1680363874
transform 1 0 464 0 1 4570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1680363874
transform 1 0 472 0 1 4570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1680363874
transform 1 0 480 0 1 4570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1680363874
transform 1 0 488 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_107
timestamp 1680363874
transform 1 0 508 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_3
timestamp 1680363874
transform 1 0 496 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_4
timestamp 1680363874
transform 1 0 592 0 1 4570
box -9 -3 26 105
use FILL  FILL_38
timestamp 1680363874
transform 1 0 608 0 1 4570
box -8 -3 16 105
use FILL  FILL_39
timestamp 1680363874
transform 1 0 616 0 1 4570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1680363874
transform 1 0 624 0 1 4570
box -8 -3 16 105
use FILL  FILL_47
timestamp 1680363874
transform 1 0 632 0 1 4570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1680363874
transform 1 0 640 0 1 4570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1680363874
transform 1 0 648 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_108
timestamp 1680363874
transform 1 0 676 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_4
timestamp 1680363874
transform 1 0 656 0 1 4570
box -8 -3 104 105
use FILL  FILL_50
timestamp 1680363874
transform 1 0 752 0 1 4570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1680363874
transform 1 0 760 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_109
timestamp 1680363874
transform 1 0 780 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_5
timestamp 1680363874
transform 1 0 768 0 1 4570
box -8 -3 104 105
use FILL  FILL_52
timestamp 1680363874
transform 1 0 864 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_5
timestamp 1680363874
transform 1 0 872 0 1 4570
box -9 -3 26 105
use FILL  FILL_53
timestamp 1680363874
transform 1 0 888 0 1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_7
timestamp 1680363874
transform 1 0 896 0 1 4570
box -8 -3 46 105
use FILL  FILL_54
timestamp 1680363874
transform 1 0 936 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_110
timestamp 1680363874
transform 1 0 956 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_6
timestamp 1680363874
transform 1 0 944 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_7
timestamp 1680363874
transform 1 0 1040 0 1 4570
box -9 -3 26 105
use FILL  FILL_70
timestamp 1680363874
transform 1 0 1056 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_111
timestamp 1680363874
transform 1 0 1076 0 1 4575
box -3 -3 3 3
use FILL  FILL_71
timestamp 1680363874
transform 1 0 1064 0 1 4570
box -8 -3 16 105
use FILL  FILL_72
timestamp 1680363874
transform 1 0 1072 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_112
timestamp 1680363874
transform 1 0 1148 0 1 4575
box -3 -3 3 3
use OAI22X1  OAI22X1_10
timestamp 1680363874
transform 1 0 1080 0 1 4570
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1680363874
transform 1 0 1120 0 1 4570
box -8 -3 46 105
use FILL  FILL_85
timestamp 1680363874
transform 1 0 1160 0 1 4570
box -8 -3 16 105
use FILL  FILL_87
timestamp 1680363874
transform 1 0 1168 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1680363874
transform 1 0 1176 0 1 4570
box -8 -3 104 105
use FILL  FILL_89
timestamp 1680363874
transform 1 0 1272 0 1 4570
box -8 -3 16 105
use FILL  FILL_90
timestamp 1680363874
transform 1 0 1280 0 1 4570
box -8 -3 16 105
use FILL  FILL_91
timestamp 1680363874
transform 1 0 1288 0 1 4570
box -8 -3 16 105
use FILL  FILL_92
timestamp 1680363874
transform 1 0 1296 0 1 4570
box -8 -3 16 105
use FILL  FILL_93
timestamp 1680363874
transform 1 0 1304 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_8
timestamp 1680363874
transform -1 0 1328 0 1 4570
box -9 -3 26 105
use FILL  FILL_94
timestamp 1680363874
transform 1 0 1328 0 1 4570
box -8 -3 16 105
use FILL  FILL_95
timestamp 1680363874
transform 1 0 1336 0 1 4570
box -8 -3 16 105
use FILL  FILL_96
timestamp 1680363874
transform 1 0 1344 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1680363874
transform -1 0 1448 0 1 4570
box -8 -3 104 105
use FILL  FILL_97
timestamp 1680363874
transform 1 0 1448 0 1 4570
box -8 -3 16 105
use FILL  FILL_98
timestamp 1680363874
transform 1 0 1456 0 1 4570
box -8 -3 16 105
use FILL  FILL_99
timestamp 1680363874
transform 1 0 1464 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1680363874
transform 1 0 1472 0 1 4570
box -8 -3 104 105
use FILL  FILL_100
timestamp 1680363874
transform 1 0 1568 0 1 4570
box -8 -3 16 105
use FILL  FILL_101
timestamp 1680363874
transform 1 0 1576 0 1 4570
box -8 -3 16 105
use FILL  FILL_102
timestamp 1680363874
transform 1 0 1584 0 1 4570
box -8 -3 16 105
use FILL  FILL_103
timestamp 1680363874
transform 1 0 1592 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1680363874
transform -1 0 1616 0 1 4570
box -9 -3 26 105
use FILL  FILL_104
timestamp 1680363874
transform 1 0 1616 0 1 4570
box -8 -3 16 105
use FILL  FILL_105
timestamp 1680363874
transform 1 0 1624 0 1 4570
box -8 -3 16 105
use FILL  FILL_106
timestamp 1680363874
transform 1 0 1632 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1680363874
transform 1 0 1640 0 1 4570
box -8 -3 104 105
use FILL  FILL_107
timestamp 1680363874
transform 1 0 1736 0 1 4570
box -8 -3 16 105
use FILL  FILL_122
timestamp 1680363874
transform 1 0 1744 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1680363874
transform 1 0 1752 0 1 4570
box -9 -3 26 105
use FILL  FILL_123
timestamp 1680363874
transform 1 0 1768 0 1 4570
box -8 -3 16 105
use FILL  FILL_124
timestamp 1680363874
transform 1 0 1776 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1680363874
transform -1 0 1880 0 1 4570
box -8 -3 104 105
use FILL  FILL_125
timestamp 1680363874
transform 1 0 1880 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_113
timestamp 1680363874
transform 1 0 1972 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_14
timestamp 1680363874
transform -1 0 1984 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_15
timestamp 1680363874
transform 1 0 1984 0 1 4570
box -9 -3 26 105
use FILL  FILL_126
timestamp 1680363874
transform 1 0 2000 0 1 4570
box -8 -3 16 105
use FILL  FILL_127
timestamp 1680363874
transform 1 0 2008 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_114
timestamp 1680363874
transform 1 0 2100 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_15
timestamp 1680363874
transform -1 0 2112 0 1 4570
box -8 -3 104 105
use FILL  FILL_128
timestamp 1680363874
transform 1 0 2112 0 1 4570
box -8 -3 16 105
use FILL  FILL_129
timestamp 1680363874
transform 1 0 2120 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1680363874
transform 1 0 2128 0 1 4570
box -8 -3 104 105
use FILL  FILL_130
timestamp 1680363874
transform 1 0 2224 0 1 4570
box -8 -3 16 105
use FILL  FILL_131
timestamp 1680363874
transform 1 0 2232 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_16
timestamp 1680363874
transform 1 0 2240 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1680363874
transform -1 0 2352 0 1 4570
box -8 -3 104 105
use FILL  FILL_132
timestamp 1680363874
transform 1 0 2352 0 1 4570
box -8 -3 16 105
use FILL  FILL_162
timestamp 1680363874
transform 1 0 2360 0 1 4570
box -8 -3 16 105
use FILL  FILL_164
timestamp 1680363874
transform 1 0 2368 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1680363874
transform 1 0 2376 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1680363874
transform -1 0 2488 0 1 4570
box -8 -3 104 105
use FILL  FILL_166
timestamp 1680363874
transform 1 0 2488 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1680363874
transform 1 0 2496 0 1 4570
box -8 -3 104 105
use FILL  FILL_177
timestamp 1680363874
transform 1 0 2592 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1680363874
transform 1 0 2600 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_21
timestamp 1680363874
transform 1 0 2696 0 1 4570
box -9 -3 26 105
use FILL  FILL_178
timestamp 1680363874
transform 1 0 2712 0 1 4570
box -8 -3 16 105
use FILL  FILL_185
timestamp 1680363874
transform 1 0 2720 0 1 4570
box -8 -3 16 105
use FILL  FILL_187
timestamp 1680363874
transform 1 0 2728 0 1 4570
box -8 -3 16 105
use FILL  FILL_189
timestamp 1680363874
transform 1 0 2736 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1680363874
transform -1 0 2840 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_23
timestamp 1680363874
transform 1 0 2840 0 1 4570
box -9 -3 26 105
use FILL  FILL_190
timestamp 1680363874
transform 1 0 2856 0 1 4570
box -8 -3 16 105
use FILL  FILL_191
timestamp 1680363874
transform 1 0 2864 0 1 4570
box -8 -3 16 105
use FILL  FILL_202
timestamp 1680363874
transform 1 0 2872 0 1 4570
box -8 -3 16 105
use FILL  FILL_204
timestamp 1680363874
transform 1 0 2880 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1680363874
transform -1 0 2984 0 1 4570
box -8 -3 104 105
use FILL  FILL_205
timestamp 1680363874
transform 1 0 2984 0 1 4570
box -8 -3 16 105
use FILL  FILL_206
timestamp 1680363874
transform 1 0 2992 0 1 4570
box -8 -3 16 105
use FILL  FILL_207
timestamp 1680363874
transform 1 0 3000 0 1 4570
box -8 -3 16 105
use FILL  FILL_208
timestamp 1680363874
transform 1 0 3008 0 1 4570
box -8 -3 16 105
use FILL  FILL_209
timestamp 1680363874
transform 1 0 3016 0 1 4570
box -8 -3 16 105
use FILL  FILL_210
timestamp 1680363874
transform 1 0 3024 0 1 4570
box -8 -3 16 105
use FILL  FILL_211
timestamp 1680363874
transform 1 0 3032 0 1 4570
box -8 -3 16 105
use FILL  FILL_212
timestamp 1680363874
transform 1 0 3040 0 1 4570
box -8 -3 16 105
use FILL  FILL_213
timestamp 1680363874
transform 1 0 3048 0 1 4570
box -8 -3 16 105
use FILL  FILL_214
timestamp 1680363874
transform 1 0 3056 0 1 4570
box -8 -3 16 105
use FILL  FILL_215
timestamp 1680363874
transform 1 0 3064 0 1 4570
box -8 -3 16 105
use FILL  FILL_216
timestamp 1680363874
transform 1 0 3072 0 1 4570
box -8 -3 16 105
use FILL  FILL_217
timestamp 1680363874
transform 1 0 3080 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_115
timestamp 1680363874
transform 1 0 3100 0 1 4575
box -3 -3 3 3
use FILL  FILL_218
timestamp 1680363874
transform 1 0 3088 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_116
timestamp 1680363874
transform 1 0 3188 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_24
timestamp 1680363874
transform -1 0 3192 0 1 4570
box -8 -3 104 105
use FILL  FILL_219
timestamp 1680363874
transform 1 0 3192 0 1 4570
box -8 -3 16 105
use FILL  FILL_220
timestamp 1680363874
transform 1 0 3200 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_117
timestamp 1680363874
transform 1 0 3220 0 1 4575
box -3 -3 3 3
use FILL  FILL_221
timestamp 1680363874
transform 1 0 3208 0 1 4570
box -8 -3 16 105
use FILL  FILL_222
timestamp 1680363874
transform 1 0 3216 0 1 4570
box -8 -3 16 105
use FILL  FILL_223
timestamp 1680363874
transform 1 0 3224 0 1 4570
box -8 -3 16 105
use FILL  FILL_224
timestamp 1680363874
transform 1 0 3232 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1680363874
transform 1 0 3240 0 1 4570
box -8 -3 104 105
use FILL  FILL_237
timestamp 1680363874
transform 1 0 3336 0 1 4570
box -8 -3 16 105
use FILL  FILL_238
timestamp 1680363874
transform 1 0 3344 0 1 4570
box -8 -3 16 105
use FILL  FILL_246
timestamp 1680363874
transform 1 0 3352 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1680363874
transform 1 0 3360 0 1 4570
box -8 -3 104 105
use FILL  FILL_248
timestamp 1680363874
transform 1 0 3456 0 1 4570
box -8 -3 16 105
use FILL  FILL_249
timestamp 1680363874
transform 1 0 3464 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1680363874
transform -1 0 3568 0 1 4570
box -8 -3 104 105
use FILL  FILL_250
timestamp 1680363874
transform 1 0 3568 0 1 4570
box -8 -3 16 105
use FILL  FILL_259
timestamp 1680363874
transform 1 0 3576 0 1 4570
box -8 -3 16 105
use FILL  FILL_260
timestamp 1680363874
transform 1 0 3584 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1680363874
transform -1 0 3688 0 1 4570
box -8 -3 104 105
use FILL  FILL_261
timestamp 1680363874
transform 1 0 3688 0 1 4570
box -8 -3 16 105
use FILL  FILL_262
timestamp 1680363874
transform 1 0 3696 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1680363874
transform -1 0 3800 0 1 4570
box -8 -3 104 105
use FILL  FILL_263
timestamp 1680363874
transform 1 0 3800 0 1 4570
box -8 -3 16 105
use FILL  FILL_264
timestamp 1680363874
transform 1 0 3808 0 1 4570
box -8 -3 16 105
use FILL  FILL_265
timestamp 1680363874
transform 1 0 3816 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_118
timestamp 1680363874
transform 1 0 3852 0 1 4575
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1680363874
transform 1 0 3908 0 1 4575
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1680363874
transform 1 0 4004 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_31
timestamp 1680363874
transform -1 0 3920 0 1 4570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1680363874
transform -1 0 4016 0 1 4570
box -8 -3 104 105
use M3_M2  M3_M2_121
timestamp 1680363874
transform 1 0 4028 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_33
timestamp 1680363874
transform 1 0 4016 0 1 4570
box -8 -3 104 105
use FILL  FILL_266
timestamp 1680363874
transform 1 0 4112 0 1 4570
box -8 -3 16 105
use FILL  FILL_267
timestamp 1680363874
transform 1 0 4120 0 1 4570
box -8 -3 16 105
use FILL  FILL_268
timestamp 1680363874
transform 1 0 4128 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1680363874
transform 1 0 4136 0 1 4570
box -8 -3 104 105
use FILL  FILL_269
timestamp 1680363874
transform 1 0 4232 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1680363874
transform -1 0 4256 0 1 4570
box -9 -3 26 105
use FILL  FILL_270
timestamp 1680363874
transform 1 0 4256 0 1 4570
box -8 -3 16 105
use FILL  FILL_271
timestamp 1680363874
transform 1 0 4264 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_122
timestamp 1680363874
transform 1 0 4284 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_35
timestamp 1680363874
transform 1 0 4272 0 1 4570
box -8 -3 104 105
use FILL  FILL_272
timestamp 1680363874
transform 1 0 4368 0 1 4570
box -8 -3 16 105
use FILL  FILL_273
timestamp 1680363874
transform 1 0 4376 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1680363874
transform -1 0 4480 0 1 4570
box -8 -3 104 105
use FILL  FILL_274
timestamp 1680363874
transform 1 0 4480 0 1 4570
box -8 -3 16 105
use FILL  FILL_304
timestamp 1680363874
transform 1 0 4488 0 1 4570
box -8 -3 16 105
use FILL  FILL_306
timestamp 1680363874
transform 1 0 4496 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_123
timestamp 1680363874
transform 1 0 4588 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_42
timestamp 1680363874
transform -1 0 4600 0 1 4570
box -8 -3 104 105
use FILL  FILL_308
timestamp 1680363874
transform 1 0 4600 0 1 4570
box -8 -3 16 105
use FILL  FILL_309
timestamp 1680363874
transform 1 0 4608 0 1 4570
box -8 -3 16 105
use FILL  FILL_310
timestamp 1680363874
transform 1 0 4616 0 1 4570
box -8 -3 16 105
use FILL  FILL_311
timestamp 1680363874
transform 1 0 4624 0 1 4570
box -8 -3 16 105
use FILL  FILL_312
timestamp 1680363874
transform 1 0 4632 0 1 4570
box -8 -3 16 105
use FILL  FILL_313
timestamp 1680363874
transform 1 0 4640 0 1 4570
box -8 -3 16 105
use FILL  FILL_314
timestamp 1680363874
transform 1 0 4648 0 1 4570
box -8 -3 16 105
use FILL  FILL_315
timestamp 1680363874
transform 1 0 4656 0 1 4570
box -8 -3 16 105
use FILL  FILL_316
timestamp 1680363874
transform 1 0 4664 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_124
timestamp 1680363874
transform 1 0 4684 0 1 4575
box -3 -3 3 3
use FILL  FILL_317
timestamp 1680363874
transform 1 0 4672 0 1 4570
box -8 -3 16 105
use FILL  FILL_318
timestamp 1680363874
transform 1 0 4680 0 1 4570
box -8 -3 16 105
use FILL  FILL_319
timestamp 1680363874
transform 1 0 4688 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_125
timestamp 1680363874
transform 1 0 4780 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_43
timestamp 1680363874
transform -1 0 4792 0 1 4570
box -8 -3 104 105
use FILL  FILL_320
timestamp 1680363874
transform 1 0 4792 0 1 4570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_3
timestamp 1680363874
transform 1 0 4827 0 1 4570
box -10 -3 10 3
use M2_M1  M2_M1_137
timestamp 1680363874
transform 1 0 68 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1680363874
transform 1 0 116 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_176
timestamp 1680363874
transform 1 0 132 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1680363874
transform 1 0 132 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1680363874
transform 1 0 148 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1680363874
transform 1 0 156 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_304
timestamp 1680363874
transform 1 0 156 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1680363874
transform 1 0 188 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1680363874
transform 1 0 188 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_140
timestamp 1680363874
transform 1 0 188 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1680363874
transform 1 0 212 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_127
timestamp 1680363874
transform 1 0 228 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1680363874
transform 1 0 308 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1680363874
transform 1 0 300 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1680363874
transform 1 0 276 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_141
timestamp 1680363874
transform 1 0 276 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1680363874
transform 1 0 292 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1680363874
transform 1 0 308 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1680363874
transform 1 0 284 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1680363874
transform 1 0 300 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1680363874
transform 1 0 308 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_256
timestamp 1680363874
transform 1 0 308 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1680363874
transform 1 0 284 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1680363874
transform 1 0 324 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1680363874
transform 1 0 340 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_214
timestamp 1680363874
transform 1 0 348 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1680363874
transform 1 0 324 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_284
timestamp 1680363874
transform 1 0 348 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1680363874
transform 1 0 380 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1680363874
transform 1 0 396 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_129
timestamp 1680363874
transform 1 0 460 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1680363874
transform 1 0 436 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1680363874
transform 1 0 452 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1680363874
transform 1 0 428 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1680363874
transform 1 0 452 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1680363874
transform 1 0 468 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_286
timestamp 1680363874
transform 1 0 460 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1680363874
transform 1 0 468 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1680363874
transform 1 0 484 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1680363874
transform 1 0 492 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1680363874
transform 1 0 508 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1680363874
transform 1 0 484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1680363874
transform 1 0 476 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1680363874
transform 1 0 532 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1680363874
transform 1 0 524 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_147
timestamp 1680363874
transform 1 0 564 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1680363874
transform 1 0 548 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1680363874
transform 1 0 564 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1680363874
transform 1 0 572 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1680363874
transform 1 0 532 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1680363874
transform 1 0 540 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1680363874
transform 1 0 556 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_306
timestamp 1680363874
transform 1 0 548 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1680363874
transform 1 0 556 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1680363874
transform 1 0 540 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_291
timestamp 1680363874
transform 1 0 580 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_257
timestamp 1680363874
transform 1 0 572 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1680363874
transform 1 0 580 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1680363874
transform 1 0 604 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1680363874
transform 1 0 620 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1680363874
transform 1 0 604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1680363874
transform 1 0 620 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1680363874
transform 1 0 612 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_332
timestamp 1680363874
transform 1 0 612 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1680363874
transform 1 0 620 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1680363874
transform 1 0 644 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1680363874
transform 1 0 684 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1680363874
transform 1 0 636 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1680363874
transform 1 0 644 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1680363874
transform 1 0 660 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1680363874
transform 1 0 676 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1680363874
transform 1 0 684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1680363874
transform 1 0 652 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1680363874
transform 1 0 716 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_183
timestamp 1680363874
transform 1 0 740 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_164
timestamp 1680363874
transform 1 0 740 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1680363874
transform 1 0 756 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1680363874
transform 1 0 724 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1680363874
transform 1 0 732 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1680363874
transform 1 0 748 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1680363874
transform 1 0 764 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1680363874
transform 1 0 724 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1680363874
transform 1 0 780 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1680363874
transform 1 0 772 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1680363874
transform 1 0 780 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1680363874
transform 1 0 764 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1680363874
transform 1 0 748 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1680363874
transform 1 0 732 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1680363874
transform 1 0 836 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1680363874
transform 1 0 828 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1680363874
transform 1 0 812 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1680363874
transform 1 0 820 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1680363874
transform 1 0 836 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1680363874
transform 1 0 852 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_427
timestamp 1680363874
transform 1 0 860 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1680363874
transform 1 0 884 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1680363874
transform 1 0 900 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1680363874
transform 1 0 908 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1680363874
transform 1 0 916 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1680363874
transform 1 0 892 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1680363874
transform 1 0 876 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_260
timestamp 1680363874
transform 1 0 884 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1680363874
transform 1 0 900 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1680363874
transform 1 0 908 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_219
timestamp 1680363874
transform 1 0 924 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1680363874
transform 1 0 940 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_172
timestamp 1680363874
transform 1 0 932 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1680363874
transform 1 0 892 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1680363874
transform 1 0 916 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1680363874
transform 1 0 924 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_429
timestamp 1680363874
transform 1 0 932 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_307
timestamp 1680363874
transform 1 0 908 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_173
timestamp 1680363874
transform 1 0 940 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1680363874
transform 1 0 972 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1680363874
transform 1 0 988 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1680363874
transform 1 0 980 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_230
timestamp 1680363874
transform 1 0 988 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_176
timestamp 1680363874
transform 1 0 1012 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1680363874
transform 1 0 1004 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_262
timestamp 1680363874
transform 1 0 980 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1680363874
transform 1 0 1020 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1680363874
transform 1 0 1060 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1680363874
transform 1 0 1060 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1680363874
transform 1 0 1068 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1680363874
transform 1 0 1092 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1680363874
transform 1 0 1092 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1680363874
transform 1 0 1052 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1680363874
transform 1 0 1068 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1680363874
transform 1 0 1084 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1680363874
transform 1 0 1060 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1680363874
transform 1 0 1076 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1680363874
transform 1 0 1076 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1680363874
transform 1 0 1052 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_305
timestamp 1680363874
transform 1 0 1092 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_264
timestamp 1680363874
transform 1 0 1100 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1680363874
transform 1 0 1124 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1680363874
transform 1 0 1132 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_180
timestamp 1680363874
transform 1 0 1124 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1680363874
transform 1 0 1140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1680363874
transform 1 0 1156 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1680363874
transform 1 0 1148 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1680363874
transform 1 0 1180 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1680363874
transform 1 0 1180 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1680363874
transform 1 0 1204 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1680363874
transform 1 0 1220 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1680363874
transform 1 0 1196 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1680363874
transform 1 0 1212 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1680363874
transform 1 0 1228 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_265
timestamp 1680363874
transform 1 0 1196 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1680363874
transform 1 0 1228 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1680363874
transform 1 0 1212 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1680363874
transform 1 0 1292 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1680363874
transform 1 0 1276 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_186
timestamp 1680363874
transform 1 0 1252 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1680363874
transform 1 0 1260 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1680363874
transform 1 0 1276 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_221
timestamp 1680363874
transform 1 0 1284 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1680363874
transform 1 0 1332 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1680363874
transform 1 0 1348 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1680363874
transform 1 0 1436 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1680363874
transform 1 0 1372 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1680363874
transform 1 0 1396 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1680363874
transform 1 0 1436 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1680363874
transform 1 0 1292 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1680363874
transform 1 0 1300 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1680363874
transform 1 0 1316 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1680363874
transform 1 0 1332 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1680363874
transform 1 0 1348 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1680363874
transform 1 0 1260 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_310
timestamp 1680363874
transform 1 0 1268 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1680363874
transform 1 0 1284 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1680363874
transform 1 0 1300 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_312
timestamp 1680363874
transform 1 0 1308 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1680363874
transform 1 0 1324 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_309
timestamp 1680363874
transform 1 0 1324 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1680363874
transform 1 0 1388 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_194
timestamp 1680363874
transform 1 0 1436 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1680363874
transform 1 0 1452 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1680363874
transform 1 0 1372 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1680363874
transform 1 0 1428 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1680363874
transform 1 0 1444 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1680363874
transform 1 0 1452 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1680363874
transform 1 0 1348 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1680363874
transform 1 0 1372 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1680363874
transform 1 0 1396 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1680363874
transform 1 0 1420 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1680363874
transform 1 0 1436 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1680363874
transform 1 0 1484 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1680363874
transform 1 0 1516 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1680363874
transform 1 0 1476 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1680363874
transform 1 0 1492 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1680363874
transform 1 0 1500 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1680363874
transform 1 0 1516 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1680363874
transform 1 0 1532 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1680363874
transform 1 0 1468 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1680363874
transform 1 0 1484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1680363874
transform 1 0 1500 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_319
timestamp 1680363874
transform 1 0 1508 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1680363874
transform 1 0 1524 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1680363874
transform 1 0 1508 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1680363874
transform 1 0 1524 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1680363874
transform 1 0 1492 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1680363874
transform 1 0 1468 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1680363874
transform 1 0 1532 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1680363874
transform 1 0 1620 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1680363874
transform 1 0 1588 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_201
timestamp 1680363874
transform 1 0 1564 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1680363874
transform 1 0 1588 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1680363874
transform 1 0 1644 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1680363874
transform 1 0 1652 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_274
timestamp 1680363874
transform 1 0 1652 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1680363874
transform 1 0 1660 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1680363874
transform 1 0 1668 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_275
timestamp 1680363874
transform 1 0 1668 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1680363874
transform 1 0 1676 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1680363874
transform 1 0 1716 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_158
timestamp 1680363874
transform 1 0 1756 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1680363874
transform 1 0 1756 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1680363874
transform 1 0 1820 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1680363874
transform 1 0 1796 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1680363874
transform 1 0 1788 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1680363874
transform 1 0 1796 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1680363874
transform 1 0 1820 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1680363874
transform 1 0 1748 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1680363874
transform 1 0 1764 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1680363874
transform 1 0 1780 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1680363874
transform 1 0 1748 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_329
timestamp 1680363874
transform 1 0 1812 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1680363874
transform 1 0 1820 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1680363874
transform 1 0 1836 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_330
timestamp 1680363874
transform 1 0 1828 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_276
timestamp 1680363874
transform 1 0 1812 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1680363874
transform 1 0 1828 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1680363874
transform 1 0 1924 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1680363874
transform 1 0 1924 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1680363874
transform 1 0 1844 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1680363874
transform 1 0 1884 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1680363874
transform 1 0 1948 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1680363874
transform 1 0 1980 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1680363874
transform 1 0 1972 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_209
timestamp 1680363874
transform 1 0 1948 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1680363874
transform 1 0 1964 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1680363874
transform 1 0 1900 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1680363874
transform 1 0 1940 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1680363874
transform 1 0 1956 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_237
timestamp 1680363874
transform 1 0 1964 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1680363874
transform 1 0 1980 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1680363874
transform 1 0 1972 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1680363874
transform 1 0 1980 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_313
timestamp 1680363874
transform 1 0 1940 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1680363874
transform 1 0 1980 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1680363874
transform 1 0 1972 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_212
timestamp 1680363874
transform 1 0 2020 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1680363874
transform 1 0 2036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1680363874
transform 1 0 1996 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1680363874
transform 1 0 2012 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1680363874
transform 1 0 2028 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_279
timestamp 1680363874
transform 1 0 2012 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1680363874
transform 1 0 2036 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1680363874
transform 1 0 2028 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1680363874
transform 1 0 2036 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_340
timestamp 1680363874
transform 1 0 2060 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1680363874
transform 1 0 2068 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1680363874
transform 1 0 2068 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1680363874
transform 1 0 2084 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1680363874
transform 1 0 2108 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_214
timestamp 1680363874
transform 1 0 2100 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1680363874
transform 1 0 2108 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1680363874
transform 1 0 2132 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1680363874
transform 1 0 2140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1680363874
transform 1 0 2108 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1680363874
transform 1 0 2124 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1680363874
transform 1 0 2132 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_344
timestamp 1680363874
transform 1 0 2148 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1680363874
transform 1 0 2148 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_345
timestamp 1680363874
transform 1 0 2164 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1680363874
transform 1 0 2172 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_282
timestamp 1680363874
transform 1 0 2172 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1680363874
transform 1 0 2212 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1680363874
transform 1 0 2220 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1680363874
transform 1 0 2236 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1680363874
transform 1 0 2244 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1680363874
transform 1 0 2260 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1680363874
transform 1 0 2244 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_139
timestamp 1680363874
transform 1 0 2276 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1680363874
transform 1 0 2276 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1680363874
transform 1 0 2236 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1680363874
transform 1 0 2252 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1680363874
transform 1 0 2268 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1680363874
transform 1 0 2372 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_163
timestamp 1680363874
transform 1 0 2412 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1680363874
transform 1 0 2404 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1680363874
transform 1 0 2412 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1680363874
transform 1 0 2396 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_223
timestamp 1680363874
transform 1 0 2428 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_352
timestamp 1680363874
transform 1 0 2444 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1680363874
transform 1 0 2452 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_283
timestamp 1680363874
transform 1 0 2444 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_222
timestamp 1680363874
transform 1 0 2508 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1680363874
transform 1 0 2532 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1680363874
transform 1 0 2548 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1680363874
transform 1 0 2524 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1680363874
transform 1 0 2540 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_240
timestamp 1680363874
transform 1 0 2548 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_356
timestamp 1680363874
transform 1 0 2556 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_317
timestamp 1680363874
transform 1 0 2540 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1680363874
transform 1 0 2524 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1680363874
transform 1 0 2612 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_225
timestamp 1680363874
transform 1 0 2580 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1680363874
transform 1 0 2588 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1680363874
transform 1 0 2580 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1680363874
transform 1 0 2588 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_227
timestamp 1680363874
transform 1 0 2620 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1680363874
transform 1 0 2596 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1680363874
transform 1 0 2612 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_284
timestamp 1680363874
transform 1 0 2580 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1680363874
transform 1 0 2620 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1680363874
transform 1 0 2636 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_228
timestamp 1680363874
transform 1 0 2636 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1680363874
transform 1 0 2652 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1680363874
transform 1 0 2628 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1680363874
transform 1 0 2628 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1680363874
transform 1 0 2716 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1680363874
transform 1 0 2684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1680363874
transform 1 0 2700 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1680363874
transform 1 0 2708 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1680363874
transform 1 0 2660 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1680363874
transform 1 0 2676 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1680363874
transform 1 0 2692 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1680363874
transform 1 0 2700 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1680363874
transform 1 0 2676 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1680363874
transform 1 0 2660 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1680363874
transform 1 0 2716 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1680363874
transform 1 0 2732 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_364
timestamp 1680363874
transform 1 0 2732 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1680363874
transform 1 0 2764 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1680363874
transform 1 0 2764 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1680363874
transform 1 0 2796 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1680363874
transform 1 0 2828 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1680363874
transform 1 0 2860 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1680363874
transform 1 0 2860 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_234
timestamp 1680363874
transform 1 0 2852 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1680363874
transform 1 0 2860 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1680363874
transform 1 0 2868 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1680363874
transform 1 0 2828 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1680363874
transform 1 0 2844 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1680363874
transform 1 0 2852 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1680363874
transform 1 0 2828 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_368
timestamp 1680363874
transform 1 0 2876 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1680363874
transform 1 0 2876 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1680363874
transform 1 0 2892 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1680363874
transform 1 0 2908 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1680363874
transform 1 0 2948 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1680363874
transform 1 0 2972 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1680363874
transform 1 0 2956 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1680363874
transform 1 0 2964 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1680363874
transform 1 0 2932 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1680363874
transform 1 0 2948 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1680363874
transform 1 0 2956 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1680363874
transform 1 0 2964 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1680363874
transform 1 0 2972 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1680363874
transform 1 0 2964 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_240
timestamp 1680363874
transform 1 0 3084 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1680363874
transform 1 0 3116 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1680363874
transform 1 0 3124 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1680363874
transform 1 0 3140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1680363874
transform 1 0 3004 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1680363874
transform 1 0 3060 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1680363874
transform 1 0 3100 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1680363874
transform 1 0 3108 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_288
timestamp 1680363874
transform 1 0 3060 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1680363874
transform 1 0 3100 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1680363874
transform 1 0 3004 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1680363874
transform 1 0 3124 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1680363874
transform 1 0 3132 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1680363874
transform 1 0 3148 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1680363874
transform 1 0 3156 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_205
timestamp 1680363874
transform 1 0 3164 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_380
timestamp 1680363874
transform 1 0 3164 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1680363874
transform 1 0 3140 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1680363874
transform 1 0 3156 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1680363874
transform 1 0 3108 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1680363874
transform 1 0 3084 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1680363874
transform 1 0 3140 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_244
timestamp 1680363874
transform 1 0 3196 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1680363874
transform 1 0 3204 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1680363874
transform 1 0 3220 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1680363874
transform 1 0 3212 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1680363874
transform 1 0 3204 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_382
timestamp 1680363874
transform 1 0 3244 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1680363874
transform 1 0 3252 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1680363874
transform 1 0 3268 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_206
timestamp 1680363874
transform 1 0 3292 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_248
timestamp 1680363874
transform 1 0 3284 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1680363874
transform 1 0 3276 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1680363874
transform 1 0 3268 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1680363874
transform 1 0 3268 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1680363874
transform 1 0 3284 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1680363874
transform 1 0 3276 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1680363874
transform 1 0 3292 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1680363874
transform 1 0 3316 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1680363874
transform 1 0 3332 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_250
timestamp 1680363874
transform 1 0 3316 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_385
timestamp 1680363874
transform 1 0 3324 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1680363874
transform 1 0 3340 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1680363874
transform 1 0 3348 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_291
timestamp 1680363874
transform 1 0 3324 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1680363874
transform 1 0 3340 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1680363874
transform 1 0 3404 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1680363874
transform 1 0 3404 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_388
timestamp 1680363874
transform 1 0 3388 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1680363874
transform 1 0 3396 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1680363874
transform 1 0 3412 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1680363874
transform 1 0 3420 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1680363874
transform 1 0 3404 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1680363874
transform 1 0 3420 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1680363874
transform 1 0 3452 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1680363874
transform 1 0 3428 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1680363874
transform 1 0 3444 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1680363874
transform 1 0 3444 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_254
timestamp 1680363874
transform 1 0 3476 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1680363874
transform 1 0 3492 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1680363874
transform 1 0 3468 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1680363874
transform 1 0 3484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_168
timestamp 1680363874
transform 1 0 3508 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1680363874
transform 1 0 3500 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1680363874
transform 1 0 3524 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_395
timestamp 1680363874
transform 1 0 3516 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1680363874
transform 1 0 3532 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1680363874
transform 1 0 3572 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1680363874
transform 1 0 3564 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1680363874
transform 1 0 3580 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_256
timestamp 1680363874
transform 1 0 3556 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1680363874
transform 1 0 3564 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1680363874
transform 1 0 3548 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1680363874
transform 1 0 3548 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1680363874
transform 1 0 3572 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_397
timestamp 1680363874
transform 1 0 3572 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1680363874
transform 1 0 3596 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1680363874
transform 1 0 3604 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_295
timestamp 1680363874
transform 1 0 3596 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1680363874
transform 1 0 3604 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_259
timestamp 1680363874
transform 1 0 3708 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1680363874
transform 1 0 3684 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1680363874
transform 1 0 3724 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_170
timestamp 1680363874
transform 1 0 3836 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1680363874
transform 1 0 3852 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1680363874
transform 1 0 3820 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1680363874
transform 1 0 3892 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1680363874
transform 1 0 3924 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1680363874
transform 1 0 3964 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1680363874
transform 1 0 3932 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1680363874
transform 1 0 3932 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1680363874
transform 1 0 3980 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1680363874
transform 1 0 4020 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_403
timestamp 1680363874
transform 1 0 4020 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1680363874
transform 1 0 4108 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_262
timestamp 1680363874
transform 1 0 4124 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1680363874
transform 1 0 4044 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1680363874
transform 1 0 4100 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_296
timestamp 1680363874
transform 1 0 4100 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1680363874
transform 1 0 4100 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1680363874
transform 1 0 4148 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1680363874
transform 1 0 4140 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_297
timestamp 1680363874
transform 1 0 4140 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1680363874
transform 1 0 4148 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1680363874
transform 1 0 4164 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1680363874
transform 1 0 4164 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1680363874
transform 1 0 4196 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1680363874
transform 1 0 4196 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1680363874
transform 1 0 4204 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1680363874
transform 1 0 4164 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1680363874
transform 1 0 4180 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1680363874
transform 1 0 4196 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1680363874
transform 1 0 4164 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1680363874
transform 1 0 4204 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1680363874
transform 1 0 4172 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1680363874
transform 1 0 4196 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_267
timestamp 1680363874
transform 1 0 4228 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1680363874
transform 1 0 4284 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1680363874
transform 1 0 4300 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1680363874
transform 1 0 4268 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_268
timestamp 1680363874
transform 1 0 4244 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1680363874
transform 1 0 4260 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1680363874
transform 1 0 4268 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1680363874
transform 1 0 4300 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1680363874
transform 1 0 4228 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1680363874
transform 1 0 4236 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1680363874
transform 1 0 4252 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1680363874
transform 1 0 4268 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1680363874
transform 1 0 4276 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1680363874
transform 1 0 4300 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1680363874
transform 1 0 4388 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1680363874
transform 1 0 4348 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1680363874
transform 1 0 4380 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_300
timestamp 1680363874
transform 1 0 4268 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1680363874
transform 1 0 4276 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1680363874
transform 1 0 4388 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_417
timestamp 1680363874
transform 1 0 4396 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1680363874
transform 1 0 4396 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_273
timestamp 1680363874
transform 1 0 4436 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1680363874
transform 1 0 4444 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1680363874
transform 1 0 4428 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1680363874
transform 1 0 4444 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1680363874
transform 1 0 4452 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1680363874
transform 1 0 4444 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1680363874
transform 1 0 4468 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_421
timestamp 1680363874
transform 1 0 4484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_302
timestamp 1680363874
transform 1 0 4492 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1680363874
transform 1 0 4588 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1680363874
transform 1 0 4684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1680363874
transform 1 0 4556 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1680363874
transform 1 0 4604 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1680363874
transform 1 0 4612 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_424
timestamp 1680363874
transform 1 0 4660 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_345
timestamp 1680363874
transform 1 0 4652 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1680363874
transform 1 0 4700 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_346
timestamp 1680363874
transform 1 0 4700 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1680363874
transform 1 0 4788 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1680363874
transform 1 0 4756 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1680363874
transform 1 0 4756 0 1 4515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_4
timestamp 1680363874
transform 1 0 24 0 1 4470
box -10 -3 10 3
use FILL  FILL_2
timestamp 1680363874
transform 1 0 72 0 -1 4570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1680363874
transform 1 0 80 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1680363874
transform 1 0 88 0 -1 4570
box -9 -3 26 105
use FILL  FILL_4
timestamp 1680363874
transform 1 0 104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1680363874
transform 1 0 112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1680363874
transform 1 0 120 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_0
timestamp 1680363874
transform 1 0 128 0 -1 4570
box -8 -3 46 105
use FILL  FILL_7
timestamp 1680363874
transform 1 0 168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1680363874
transform 1 0 176 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1680363874
transform 1 0 184 0 -1 4570
box -9 -3 26 105
use FILL  FILL_12
timestamp 1680363874
transform 1 0 200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_13
timestamp 1680363874
transform 1 0 208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_14
timestamp 1680363874
transform 1 0 216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_15
timestamp 1680363874
transform 1 0 224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_16
timestamp 1680363874
transform 1 0 232 0 -1 4570
box -8 -3 16 105
use FILL  FILL_17
timestamp 1680363874
transform 1 0 240 0 -1 4570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1680363874
transform 1 0 248 0 -1 4570
box -8 -3 16 105
use FILL  FILL_19
timestamp 1680363874
transform 1 0 256 0 -1 4570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1680363874
transform 1 0 264 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_1
timestamp 1680363874
transform -1 0 312 0 -1 4570
box -8 -3 46 105
use FILL  FILL_21
timestamp 1680363874
transform 1 0 312 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_2
timestamp 1680363874
transform 1 0 320 0 -1 4570
box -8 -3 46 105
use FILL  FILL_26
timestamp 1680363874
transform 1 0 360 0 -1 4570
box -8 -3 16 105
use FILL  FILL_27
timestamp 1680363874
transform 1 0 368 0 -1 4570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1680363874
transform 1 0 376 0 -1 4570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1680363874
transform 1 0 384 0 -1 4570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1680363874
transform 1 0 392 0 -1 4570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1680363874
transform 1 0 400 0 -1 4570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1680363874
transform 1 0 408 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_354
timestamp 1680363874
transform 1 0 428 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_3
timestamp 1680363874
transform -1 0 456 0 -1 4570
box -8 -3 46 105
use FILL  FILL_33
timestamp 1680363874
transform 1 0 456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1680363874
transform 1 0 464 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_4
timestamp 1680363874
transform -1 0 512 0 -1 4570
box -8 -3 46 105
use FILL  FILL_42
timestamp 1680363874
transform 1 0 512 0 -1 4570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1680363874
transform 1 0 520 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1680363874
transform 1 0 528 0 -1 4570
box -8 -3 46 105
use FILL  FILL_44
timestamp 1680363874
transform 1 0 568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_45
timestamp 1680363874
transform 1 0 576 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_6
timestamp 1680363874
transform 1 0 584 0 -1 4570
box -8 -3 46 105
use FILL  FILL_46
timestamp 1680363874
transform 1 0 624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1680363874
transform 1 0 632 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_355
timestamp 1680363874
transform 1 0 652 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_8
timestamp 1680363874
transform -1 0 680 0 -1 4570
box -8 -3 46 105
use FILL  FILL_56
timestamp 1680363874
transform 1 0 680 0 -1 4570
box -8 -3 16 105
use FILL  FILL_57
timestamp 1680363874
transform 1 0 688 0 -1 4570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1680363874
transform 1 0 696 0 -1 4570
box -8 -3 16 105
use FILL  FILL_59
timestamp 1680363874
transform 1 0 704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1680363874
transform 1 0 712 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1680363874
transform 1 0 720 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_6
timestamp 1680363874
transform -1 0 776 0 -1 4570
box -9 -3 26 105
use FILL  FILL_61
timestamp 1680363874
transform 1 0 776 0 -1 4570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1680363874
transform 1 0 784 0 -1 4570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1680363874
transform 1 0 792 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1680363874
transform 1 0 800 0 -1 4570
box -8 -3 34 105
use FILL  FILL_64
timestamp 1680363874
transform 1 0 832 0 -1 4570
box -8 -3 16 105
use FILL  FILL_65
timestamp 1680363874
transform 1 0 840 0 -1 4570
box -8 -3 16 105
use FILL  FILL_66
timestamp 1680363874
transform 1 0 848 0 -1 4570
box -8 -3 16 105
use FILL  FILL_67
timestamp 1680363874
transform 1 0 856 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1680363874
transform 1 0 864 0 -1 4570
box -8 -3 34 105
use FILL  FILL_68
timestamp 1680363874
transform 1 0 896 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1680363874
transform 1 0 904 0 -1 4570
box -8 -3 34 105
use FILL  FILL_69
timestamp 1680363874
transform 1 0 936 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_356
timestamp 1680363874
transform 1 0 956 0 1 4475
box -3 -3 3 3
use FILL  FILL_73
timestamp 1680363874
transform 1 0 944 0 -1 4570
box -8 -3 16 105
use FILL  FILL_74
timestamp 1680363874
transform 1 0 952 0 -1 4570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1680363874
transform 1 0 960 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_12
timestamp 1680363874
transform -1 0 1008 0 -1 4570
box -8 -3 46 105
use FILL  FILL_76
timestamp 1680363874
transform 1 0 1008 0 -1 4570
box -8 -3 16 105
use FILL  FILL_77
timestamp 1680363874
transform 1 0 1016 0 -1 4570
box -8 -3 16 105
use FILL  FILL_78
timestamp 1680363874
transform 1 0 1024 0 -1 4570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1680363874
transform 1 0 1032 0 -1 4570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1680363874
transform 1 0 1040 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_13
timestamp 1680363874
transform 1 0 1048 0 -1 4570
box -8 -3 46 105
use FILL  FILL_81
timestamp 1680363874
transform 1 0 1088 0 -1 4570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1680363874
transform 1 0 1096 0 -1 4570
box -8 -3 16 105
use FILL  FILL_83
timestamp 1680363874
transform 1 0 1104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_84
timestamp 1680363874
transform 1 0 1112 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_357
timestamp 1680363874
transform 1 0 1140 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_14
timestamp 1680363874
transform 1 0 1120 0 -1 4570
box -8 -3 46 105
use FILL  FILL_86
timestamp 1680363874
transform 1 0 1160 0 -1 4570
box -8 -3 16 105
use FILL  FILL_88
timestamp 1680363874
transform 1 0 1168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_108
timestamp 1680363874
transform 1 0 1176 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_15
timestamp 1680363874
transform 1 0 1184 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_10
timestamp 1680363874
transform -1 0 1240 0 -1 4570
box -9 -3 26 105
use FILL  FILL_109
timestamp 1680363874
transform 1 0 1240 0 -1 4570
box -8 -3 16 105
use FILL  FILL_110
timestamp 1680363874
transform 1 0 1248 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_16
timestamp 1680363874
transform -1 0 1296 0 -1 4570
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1680363874
transform -1 0 1336 0 -1 4570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1680363874
transform 1 0 1336 0 -1 4570
box -8 -3 104 105
use INVX2  INVX2_11
timestamp 1680363874
transform 1 0 1432 0 -1 4570
box -9 -3 26 105
use FILL  FILL_111
timestamp 1680363874
transform 1 0 1448 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_18
timestamp 1680363874
transform -1 0 1496 0 -1 4570
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1680363874
transform -1 0 1536 0 -1 4570
box -8 -3 46 105
use FILL  FILL_112
timestamp 1680363874
transform 1 0 1536 0 -1 4570
box -8 -3 16 105
use FILL  FILL_113
timestamp 1680363874
transform 1 0 1544 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1680363874
transform 1 0 1552 0 -1 4570
box -8 -3 104 105
use INVX2  INVX2_12
timestamp 1680363874
transform -1 0 1664 0 -1 4570
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1680363874
transform 1 0 1664 0 -1 4570
box -9 -3 26 105
use FILL  FILL_114
timestamp 1680363874
transform 1 0 1680 0 -1 4570
box -8 -3 16 105
use FILL  FILL_115
timestamp 1680363874
transform 1 0 1688 0 -1 4570
box -8 -3 16 105
use FILL  FILL_116
timestamp 1680363874
transform 1 0 1696 0 -1 4570
box -8 -3 16 105
use FILL  FILL_117
timestamp 1680363874
transform 1 0 1704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_118
timestamp 1680363874
transform 1 0 1712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_119
timestamp 1680363874
transform 1 0 1720 0 -1 4570
box -8 -3 16 105
use FILL  FILL_120
timestamp 1680363874
transform 1 0 1728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_121
timestamp 1680363874
transform 1 0 1736 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1680363874
transform 1 0 1744 0 -1 4570
box -8 -3 46 105
use FILL  FILL_133
timestamp 1680363874
transform 1 0 1784 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1680363874
transform -1 0 1832 0 -1 4570
box -8 -3 46 105
use FILL  FILL_134
timestamp 1680363874
transform 1 0 1832 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1680363874
transform -1 0 1936 0 -1 4570
box -8 -3 104 105
use AOI22X1  AOI22X1_2
timestamp 1680363874
transform 1 0 1936 0 -1 4570
box -8 -3 46 105
use FILL  FILL_135
timestamp 1680363874
transform 1 0 1976 0 -1 4570
box -8 -3 16 105
use FILL  FILL_136
timestamp 1680363874
transform 1 0 1984 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1680363874
transform 1 0 1992 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_17
timestamp 1680363874
transform 1 0 2032 0 -1 4570
box -9 -3 26 105
use FILL  FILL_137
timestamp 1680363874
transform 1 0 2048 0 -1 4570
box -8 -3 16 105
use FILL  FILL_138
timestamp 1680363874
transform 1 0 2056 0 -1 4570
box -8 -3 16 105
use FILL  FILL_139
timestamp 1680363874
transform 1 0 2064 0 -1 4570
box -8 -3 16 105
use FILL  FILL_140
timestamp 1680363874
transform 1 0 2072 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_18
timestamp 1680363874
transform -1 0 2096 0 -1 4570
box -9 -3 26 105
use FILL  FILL_141
timestamp 1680363874
transform 1 0 2096 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1680363874
transform 1 0 2104 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_19
timestamp 1680363874
transform 1 0 2144 0 -1 4570
box -9 -3 26 105
use FILL  FILL_142
timestamp 1680363874
transform 1 0 2160 0 -1 4570
box -8 -3 16 105
use FILL  FILL_143
timestamp 1680363874
transform 1 0 2168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_144
timestamp 1680363874
transform 1 0 2176 0 -1 4570
box -8 -3 16 105
use FILL  FILL_145
timestamp 1680363874
transform 1 0 2184 0 -1 4570
box -8 -3 16 105
use FILL  FILL_146
timestamp 1680363874
transform 1 0 2192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_147
timestamp 1680363874
transform 1 0 2200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_148
timestamp 1680363874
transform 1 0 2208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_149
timestamp 1680363874
transform 1 0 2216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_150
timestamp 1680363874
transform 1 0 2224 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1680363874
transform -1 0 2272 0 -1 4570
box -8 -3 46 105
use FILL  FILL_151
timestamp 1680363874
transform 1 0 2272 0 -1 4570
box -8 -3 16 105
use FILL  FILL_152
timestamp 1680363874
transform 1 0 2280 0 -1 4570
box -8 -3 16 105
use FILL  FILL_153
timestamp 1680363874
transform 1 0 2288 0 -1 4570
box -8 -3 16 105
use FILL  FILL_154
timestamp 1680363874
transform 1 0 2296 0 -1 4570
box -8 -3 16 105
use FILL  FILL_155
timestamp 1680363874
transform 1 0 2304 0 -1 4570
box -8 -3 16 105
use FILL  FILL_156
timestamp 1680363874
transform 1 0 2312 0 -1 4570
box -8 -3 16 105
use FILL  FILL_157
timestamp 1680363874
transform 1 0 2320 0 -1 4570
box -8 -3 16 105
use FILL  FILL_158
timestamp 1680363874
transform 1 0 2328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_159
timestamp 1680363874
transform 1 0 2336 0 -1 4570
box -8 -3 16 105
use FILL  FILL_160
timestamp 1680363874
transform 1 0 2344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_161
timestamp 1680363874
transform 1 0 2352 0 -1 4570
box -8 -3 16 105
use FILL  FILL_163
timestamp 1680363874
transform 1 0 2360 0 -1 4570
box -8 -3 16 105
use FILL  FILL_165
timestamp 1680363874
transform 1 0 2368 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1680363874
transform 1 0 2376 0 -1 4570
box -8 -3 46 105
use FILL  FILL_167
timestamp 1680363874
transform 1 0 2416 0 -1 4570
box -8 -3 16 105
use FILL  FILL_168
timestamp 1680363874
transform 1 0 2424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_169
timestamp 1680363874
transform 1 0 2432 0 -1 4570
box -8 -3 16 105
use FILL  FILL_170
timestamp 1680363874
transform 1 0 2440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_171
timestamp 1680363874
transform 1 0 2448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_172
timestamp 1680363874
transform 1 0 2456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_173
timestamp 1680363874
transform 1 0 2464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_174
timestamp 1680363874
transform 1 0 2472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_175
timestamp 1680363874
transform 1 0 2480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_176
timestamp 1680363874
transform 1 0 2488 0 -1 4570
box -8 -3 16 105
use FILL  FILL_179
timestamp 1680363874
transform 1 0 2496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_180
timestamp 1680363874
transform 1 0 2504 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_20
timestamp 1680363874
transform 1 0 2512 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_22
timestamp 1680363874
transform -1 0 2568 0 -1 4570
box -9 -3 26 105
use FILL  FILL_181
timestamp 1680363874
transform 1 0 2568 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_7
timestamp 1680363874
transform -1 0 2616 0 -1 4570
box -8 -3 46 105
use FILL  FILL_182
timestamp 1680363874
transform 1 0 2616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_183
timestamp 1680363874
transform 1 0 2624 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_358
timestamp 1680363874
transform 1 0 2660 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_21
timestamp 1680363874
transform 1 0 2632 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1680363874
transform -1 0 2712 0 -1 4570
box -8 -3 46 105
use FILL  FILL_184
timestamp 1680363874
transform 1 0 2712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_186
timestamp 1680363874
transform 1 0 2720 0 -1 4570
box -8 -3 16 105
use FILL  FILL_188
timestamp 1680363874
transform 1 0 2728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_192
timestamp 1680363874
transform 1 0 2736 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_24
timestamp 1680363874
transform 1 0 2744 0 -1 4570
box -9 -3 26 105
use FILL  FILL_193
timestamp 1680363874
transform 1 0 2760 0 -1 4570
box -8 -3 16 105
use FILL  FILL_194
timestamp 1680363874
transform 1 0 2768 0 -1 4570
box -8 -3 16 105
use FILL  FILL_195
timestamp 1680363874
transform 1 0 2776 0 -1 4570
box -8 -3 16 105
use FILL  FILL_196
timestamp 1680363874
transform 1 0 2784 0 -1 4570
box -8 -3 16 105
use FILL  FILL_197
timestamp 1680363874
transform 1 0 2792 0 -1 4570
box -8 -3 16 105
use FILL  FILL_198
timestamp 1680363874
transform 1 0 2800 0 -1 4570
box -8 -3 16 105
use FILL  FILL_199
timestamp 1680363874
transform 1 0 2808 0 -1 4570
box -8 -3 16 105
use FILL  FILL_200
timestamp 1680363874
transform 1 0 2816 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_9
timestamp 1680363874
transform -1 0 2864 0 -1 4570
box -8 -3 46 105
use FILL  FILL_201
timestamp 1680363874
transform 1 0 2864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_203
timestamp 1680363874
transform 1 0 2872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_225
timestamp 1680363874
transform 1 0 2880 0 -1 4570
box -8 -3 16 105
use FILL  FILL_226
timestamp 1680363874
transform 1 0 2888 0 -1 4570
box -8 -3 16 105
use FILL  FILL_227
timestamp 1680363874
transform 1 0 2896 0 -1 4570
box -8 -3 16 105
use FILL  FILL_228
timestamp 1680363874
transform 1 0 2904 0 -1 4570
box -8 -3 16 105
use FILL  FILL_229
timestamp 1680363874
transform 1 0 2912 0 -1 4570
box -8 -3 16 105
use FILL  FILL_230
timestamp 1680363874
transform 1 0 2920 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1680363874
transform -1 0 2968 0 -1 4570
box -8 -3 46 105
use FILL  FILL_231
timestamp 1680363874
transform 1 0 2968 0 -1 4570
box -8 -3 16 105
use FILL  FILL_232
timestamp 1680363874
transform 1 0 2976 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_25
timestamp 1680363874
transform 1 0 2984 0 -1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1680363874
transform -1 0 3096 0 -1 4570
box -8 -3 104 105
use INVX2  INVX2_26
timestamp 1680363874
transform -1 0 3112 0 -1 4570
box -9 -3 26 105
use AOI22X1  AOI22X1_11
timestamp 1680363874
transform 1 0 3112 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_27
timestamp 1680363874
transform -1 0 3168 0 -1 4570
box -9 -3 26 105
use FILL  FILL_233
timestamp 1680363874
transform 1 0 3168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_234
timestamp 1680363874
transform 1 0 3176 0 -1 4570
box -8 -3 16 105
use FILL  FILL_235
timestamp 1680363874
transform 1 0 3184 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_359
timestamp 1680363874
transform 1 0 3220 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_12
timestamp 1680363874
transform 1 0 3192 0 -1 4570
box -8 -3 46 105
use FILL  FILL_236
timestamp 1680363874
transform 1 0 3232 0 -1 4570
box -8 -3 16 105
use FILL  FILL_239
timestamp 1680363874
transform 1 0 3240 0 -1 4570
box -8 -3 16 105
use FILL  FILL_240
timestamp 1680363874
transform 1 0 3248 0 -1 4570
box -8 -3 16 105
use FILL  FILL_241
timestamp 1680363874
transform 1 0 3256 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_28
timestamp 1680363874
transform 1 0 3264 0 -1 4570
box -9 -3 26 105
use FILL  FILL_242
timestamp 1680363874
transform 1 0 3280 0 -1 4570
box -8 -3 16 105
use FILL  FILL_243
timestamp 1680363874
transform 1 0 3288 0 -1 4570
box -8 -3 16 105
use FILL  FILL_244
timestamp 1680363874
transform 1 0 3296 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_13
timestamp 1680363874
transform 1 0 3304 0 -1 4570
box -8 -3 46 105
use FILL  FILL_245
timestamp 1680363874
transform 1 0 3344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_247
timestamp 1680363874
transform 1 0 3352 0 -1 4570
box -8 -3 16 105
use FILL  FILL_251
timestamp 1680363874
transform 1 0 3360 0 -1 4570
box -8 -3 16 105
use FILL  FILL_252
timestamp 1680363874
transform 1 0 3368 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_29
timestamp 1680363874
transform 1 0 3376 0 -1 4570
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1680363874
transform -1 0 3408 0 -1 4570
box -9 -3 26 105
use AOI22X1  AOI22X1_14
timestamp 1680363874
transform 1 0 3408 0 -1 4570
box -8 -3 46 105
use FILL  FILL_253
timestamp 1680363874
transform 1 0 3448 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_360
timestamp 1680363874
transform 1 0 3468 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_22
timestamp 1680363874
transform -1 0 3496 0 -1 4570
box -8 -3 46 105
use FILL  FILL_254
timestamp 1680363874
transform 1 0 3496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_255
timestamp 1680363874
transform 1 0 3504 0 -1 4570
box -8 -3 16 105
use FILL  FILL_256
timestamp 1680363874
transform 1 0 3512 0 -1 4570
box -8 -3 16 105
use FILL  FILL_257
timestamp 1680363874
transform 1 0 3520 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_15
timestamp 1680363874
transform -1 0 3568 0 -1 4570
box -8 -3 46 105
use FILL  FILL_258
timestamp 1680363874
transform 1 0 3568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_275
timestamp 1680363874
transform 1 0 3576 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_32
timestamp 1680363874
transform -1 0 3600 0 -1 4570
box -9 -3 26 105
use FILL  FILL_276
timestamp 1680363874
transform 1 0 3600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_277
timestamp 1680363874
transform 1 0 3608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_278
timestamp 1680363874
transform 1 0 3616 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1680363874
transform -1 0 3720 0 -1 4570
box -8 -3 104 105
use FILL  FILL_279
timestamp 1680363874
transform 1 0 3720 0 -1 4570
box -8 -3 16 105
use FILL  FILL_280
timestamp 1680363874
transform 1 0 3728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_281
timestamp 1680363874
transform 1 0 3736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_282
timestamp 1680363874
transform 1 0 3744 0 -1 4570
box -8 -3 16 105
use FILL  FILL_283
timestamp 1680363874
transform 1 0 3752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_284
timestamp 1680363874
transform 1 0 3760 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_361
timestamp 1680363874
transform 1 0 3788 0 1 4475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_38
timestamp 1680363874
transform -1 0 3864 0 -1 4570
box -8 -3 104 105
use FILL  FILL_285
timestamp 1680363874
transform 1 0 3864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_286
timestamp 1680363874
transform 1 0 3872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_287
timestamp 1680363874
transform 1 0 3880 0 -1 4570
box -8 -3 16 105
use FILL  FILL_288
timestamp 1680363874
transform 1 0 3888 0 -1 4570
box -8 -3 16 105
use FILL  FILL_289
timestamp 1680363874
transform 1 0 3896 0 -1 4570
box -8 -3 16 105
use FILL  FILL_290
timestamp 1680363874
transform 1 0 3904 0 -1 4570
box -8 -3 16 105
use FILL  FILL_291
timestamp 1680363874
transform 1 0 3912 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1680363874
transform 1 0 3920 0 -1 4570
box -8 -3 104 105
use FILL  FILL_292
timestamp 1680363874
transform 1 0 4016 0 -1 4570
box -8 -3 16 105
use FILL  FILL_293
timestamp 1680363874
transform 1 0 4024 0 -1 4570
box -8 -3 16 105
use FILL  FILL_294
timestamp 1680363874
transform 1 0 4032 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1680363874
transform -1 0 4136 0 -1 4570
box -8 -3 104 105
use FILL  FILL_295
timestamp 1680363874
transform 1 0 4136 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_33
timestamp 1680363874
transform 1 0 4144 0 -1 4570
box -9 -3 26 105
use AOI22X1  AOI22X1_16
timestamp 1680363874
transform -1 0 4200 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_34
timestamp 1680363874
transform 1 0 4200 0 -1 4570
box -9 -3 26 105
use FILL  FILL_296
timestamp 1680363874
transform 1 0 4216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_297
timestamp 1680363874
transform 1 0 4224 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_17
timestamp 1680363874
transform -1 0 4272 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_35
timestamp 1680363874
transform 1 0 4272 0 -1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1680363874
transform 1 0 4288 0 -1 4570
box -8 -3 104 105
use FILL  FILL_298
timestamp 1680363874
transform 1 0 4384 0 -1 4570
box -8 -3 16 105
use FILL  FILL_299
timestamp 1680363874
transform 1 0 4392 0 -1 4570
box -8 -3 16 105
use FILL  FILL_300
timestamp 1680363874
transform 1 0 4400 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_18
timestamp 1680363874
transform -1 0 4448 0 -1 4570
box -8 -3 46 105
use FILL  FILL_301
timestamp 1680363874
transform 1 0 4448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_302
timestamp 1680363874
transform 1 0 4456 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_36
timestamp 1680363874
transform 1 0 4464 0 -1 4570
box -9 -3 26 105
use FILL  FILL_303
timestamp 1680363874
transform 1 0 4480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_305
timestamp 1680363874
transform 1 0 4488 0 -1 4570
box -8 -3 16 105
use FILL  FILL_307
timestamp 1680363874
transform 1 0 4496 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1680363874
transform -1 0 4600 0 -1 4570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1680363874
transform -1 0 4696 0 -1 4570
box -8 -3 104 105
use FILL  FILL_321
timestamp 1680363874
transform 1 0 4696 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1680363874
transform -1 0 4800 0 -1 4570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_5
timestamp 1680363874
transform 1 0 4851 0 1 4470
box -10 -3 10 3
use M2_M1  M2_M1_433
timestamp 1680363874
transform 1 0 76 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1680363874
transform 1 0 132 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_434
timestamp 1680363874
transform 1 0 244 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1680363874
transform 1 0 180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1680363874
transform 1 0 244 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1680363874
transform 1 0 156 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1680363874
transform 1 0 172 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1680363874
transform 1 0 196 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_515
timestamp 1680363874
transform 1 0 196 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1680363874
transform 1 0 236 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_437
timestamp 1680363874
transform 1 0 300 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_435
timestamp 1680363874
transform 1 0 340 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_438
timestamp 1680363874
transform 1 0 364 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1680363874
transform 1 0 316 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1680363874
transform 1 0 316 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1680363874
transform 1 0 364 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1680363874
transform 1 0 396 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1680363874
transform 1 0 484 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1680363874
transform 1 0 460 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_476
timestamp 1680363874
transform 1 0 468 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1680363874
transform 1 0 476 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1680363874
transform 1 0 452 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1680363874
transform 1 0 468 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1680363874
transform 1 0 484 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_519
timestamp 1680363874
transform 1 0 468 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1680363874
transform 1 0 484 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_441
timestamp 1680363874
transform 1 0 500 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1680363874
transform 1 0 508 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_520
timestamp 1680363874
transform 1 0 500 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1680363874
transform 1 0 524 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1680363874
transform 1 0 524 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_376
timestamp 1680363874
transform 1 0 556 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1680363874
transform 1 0 548 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1680363874
transform 1 0 564 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_442
timestamp 1680363874
transform 1 0 548 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1680363874
transform 1 0 564 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1680363874
transform 1 0 556 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1680363874
transform 1 0 564 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1680363874
transform 1 0 572 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1680363874
transform 1 0 580 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1680363874
transform 1 0 556 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1680363874
transform 1 0 588 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1680363874
transform 1 0 588 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_444
timestamp 1680363874
transform 1 0 588 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_377
timestamp 1680363874
transform 1 0 636 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1680363874
transform 1 0 628 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_445
timestamp 1680363874
transform 1 0 636 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_438
timestamp 1680363874
transform 1 0 652 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_446
timestamp 1680363874
transform 1 0 652 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1680363874
transform 1 0 628 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1680363874
transform 1 0 644 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1680363874
transform 1 0 652 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_521
timestamp 1680363874
transform 1 0 652 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1680363874
transform 1 0 668 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1680363874
transform 1 0 700 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_447
timestamp 1680363874
transform 1 0 676 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1680363874
transform 1 0 692 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_448
timestamp 1680363874
transform 1 0 700 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_380
timestamp 1680363874
transform 1 0 748 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1680363874
transform 1 0 724 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_449
timestamp 1680363874
transform 1 0 724 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1680363874
transform 1 0 748 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1680363874
transform 1 0 692 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1680363874
transform 1 0 708 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1680363874
transform 1 0 716 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_440
timestamp 1680363874
transform 1 0 772 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_451
timestamp 1680363874
transform 1 0 772 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1680363874
transform 1 0 740 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1680363874
transform 1 0 756 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1680363874
transform 1 0 764 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1680363874
transform 1 0 788 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_522
timestamp 1680363874
transform 1 0 716 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1680363874
transform 1 0 740 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1680363874
transform 1 0 764 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_582
timestamp 1680363874
transform 1 0 796 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1680363874
transform 1 0 796 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1680363874
transform 1 0 820 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_430
timestamp 1680363874
transform 1 0 820 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_368
timestamp 1680363874
transform 1 0 852 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1680363874
transform 1 0 852 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1680363874
transform 1 0 852 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1680363874
transform 1 0 836 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1680363874
transform 1 0 836 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_583
timestamp 1680363874
transform 1 0 876 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_369
timestamp 1680363874
transform 1 0 892 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_584
timestamp 1680363874
transform 1 0 884 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1680363874
transform 1 0 908 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_585
timestamp 1680363874
transform 1 0 908 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_404
timestamp 1680363874
transform 1 0 924 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_586
timestamp 1680363874
transform 1 0 924 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1680363874
transform 1 0 940 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_501
timestamp 1680363874
transform 1 0 940 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1680363874
transform 1 0 972 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1680363874
transform 1 0 988 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_432
timestamp 1680363874
transform 1 0 972 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1680363874
transform 1 0 956 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_441
timestamp 1680363874
transform 1 0 996 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_455
timestamp 1680363874
transform 1 0 988 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1680363874
transform 1 0 972 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1680363874
transform 1 0 980 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1680363874
transform 1 0 996 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1680363874
transform 1 0 1012 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1680363874
transform 1 0 1028 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_406
timestamp 1680363874
transform 1 0 1044 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1680363874
transform 1 0 1076 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1680363874
transform 1 0 1060 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_457
timestamp 1680363874
transform 1 0 1060 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1680363874
transform 1 0 1076 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_443
timestamp 1680363874
transform 1 0 1092 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1680363874
transform 1 0 1092 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1680363874
transform 1 0 1052 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1680363874
transform 1 0 1068 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1680363874
transform 1 0 1084 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1680363874
transform 1 0 1092 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1680363874
transform 1 0 1068 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1680363874
transform 1 0 1092 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1680363874
transform 1 0 1148 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_460
timestamp 1680363874
transform 1 0 1148 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_502
timestamp 1680363874
transform 1 0 1132 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_461
timestamp 1680363874
transform 1 0 1164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1680363874
transform 1 0 1140 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1680363874
transform 1 0 1156 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_528
timestamp 1680363874
transform 1 0 1164 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1680363874
transform 1 0 1212 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1680363874
transform 1 0 1244 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1680363874
transform 1 0 1228 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_462
timestamp 1680363874
transform 1 0 1252 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1680363874
transform 1 0 1268 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1680363874
transform 1 0 1220 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1680363874
transform 1 0 1228 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1680363874
transform 1 0 1244 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1680363874
transform 1 0 1260 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_529
timestamp 1680363874
transform 1 0 1220 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1680363874
transform 1 0 1268 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1680363874
transform 1 0 1324 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1680363874
transform 1 0 1292 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_464
timestamp 1680363874
transform 1 0 1324 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1680363874
transform 1 0 1388 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1680363874
transform 1 0 1396 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1680363874
transform 1 0 1372 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_446
timestamp 1680363874
transform 1 0 1428 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_467
timestamp 1680363874
transform 1 0 1428 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1680363874
transform 1 0 1444 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1680363874
transform 1 0 1460 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1680363874
transform 1 0 1412 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1680363874
transform 1 0 1420 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1680363874
transform 1 0 1436 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1680363874
transform 1 0 1452 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_531
timestamp 1680363874
transform 1 0 1436 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1680363874
transform 1 0 1468 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1680363874
transform 1 0 1484 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1680363874
transform 1 0 1508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1680363874
transform 1 0 1468 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1680363874
transform 1 0 1484 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1680363874
transform 1 0 1508 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1680363874
transform 1 0 1588 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_471
timestamp 1680363874
transform 1 0 1580 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1680363874
transform 1 0 1588 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1680363874
transform 1 0 1692 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1680363874
transform 1 0 1660 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1680363874
transform 1 0 1700 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_473
timestamp 1680363874
transform 1 0 1660 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1680363874
transform 1 0 1692 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1680363874
transform 1 0 1700 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1680363874
transform 1 0 1596 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1680363874
transform 1 0 1612 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1680363874
transform 1 0 1612 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1680363874
transform 1 0 1636 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1680363874
transform 1 0 1652 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1680363874
transform 1 0 1724 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1680363874
transform 1 0 1748 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1680363874
transform 1 0 1732 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_476
timestamp 1680363874
transform 1 0 1724 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1680363874
transform 1 0 1740 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_450
timestamp 1680363874
transform 1 0 1764 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1680363874
transform 1 0 1764 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1680363874
transform 1 0 1724 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1680363874
transform 1 0 1732 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1680363874
transform 1 0 1756 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1680363874
transform 1 0 1780 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1680363874
transform 1 0 1780 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_613
timestamp 1680363874
transform 1 0 1772 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_451
timestamp 1680363874
transform 1 0 1828 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_479
timestamp 1680363874
transform 1 0 1796 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1680363874
transform 1 0 1812 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1680363874
transform 1 0 1788 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1680363874
transform 1 0 1804 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1680363874
transform 1 0 1812 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_616
timestamp 1680363874
transform 1 0 1820 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_536
timestamp 1680363874
transform 1 0 1796 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1680363874
transform 1 0 1860 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1680363874
transform 1 0 1844 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_481
timestamp 1680363874
transform 1 0 1844 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1680363874
transform 1 0 1860 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1680363874
transform 1 0 1836 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1680363874
transform 1 0 1852 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1680363874
transform 1 0 1860 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1680363874
transform 1 0 1844 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1680363874
transform 1 0 1892 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1680363874
transform 1 0 1908 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1680363874
transform 1 0 1900 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1680363874
transform 1 0 1908 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1680363874
transform 1 0 1892 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_413
timestamp 1680363874
transform 1 0 1948 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1680363874
transform 1 0 1964 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_485
timestamp 1680363874
transform 1 0 1956 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1680363874
transform 1 0 2012 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1680363874
transform 1 0 2020 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1680363874
transform 1 0 2036 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1680363874
transform 1 0 1940 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1680363874
transform 1 0 1948 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1680363874
transform 1 0 1964 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1680363874
transform 1 0 1972 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1680363874
transform 1 0 1988 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_538
timestamp 1680363874
transform 1 0 2012 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1680363874
transform 1 0 2084 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1680363874
transform 1 0 2100 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1680363874
transform 1 0 2116 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1680363874
transform 1 0 2092 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1680363874
transform 1 0 2108 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_539
timestamp 1680363874
transform 1 0 2108 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1680363874
transform 1 0 2228 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1680363874
transform 1 0 2196 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1680363874
transform 1 0 2236 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_490
timestamp 1680363874
transform 1 0 2196 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1680363874
transform 1 0 2228 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1680363874
transform 1 0 2236 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1680363874
transform 1 0 2148 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_547
timestamp 1680363874
transform 1 0 2148 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1680363874
transform 1 0 2260 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_628
timestamp 1680363874
transform 1 0 2252 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1680363874
transform 1 0 2308 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1680363874
transform 1 0 2284 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_548
timestamp 1680363874
transform 1 0 2284 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1680363874
transform 1 0 2300 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1680363874
transform 1 0 2372 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1680363874
transform 1 0 2404 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1680363874
transform 1 0 2388 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1680363874
transform 1 0 2388 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1680363874
transform 1 0 2404 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1680363874
transform 1 0 2380 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1680363874
transform 1 0 2396 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1680363874
transform 1 0 2404 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1680363874
transform 1 0 2452 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1680363874
transform 1 0 2476 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1680363874
transform 1 0 2516 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_496
timestamp 1680363874
transform 1 0 2476 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1680363874
transform 1 0 2508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1680363874
transform 1 0 2516 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1680363874
transform 1 0 2412 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1680363874
transform 1 0 2428 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_550
timestamp 1680363874
transform 1 0 2428 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1680363874
transform 1 0 2540 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_634
timestamp 1680363874
transform 1 0 2548 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_387
timestamp 1680363874
transform 1 0 2564 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1680363874
transform 1 0 2628 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1680363874
transform 1 0 2612 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1680363874
transform 1 0 2684 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_499
timestamp 1680363874
transform 1 0 2620 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1680363874
transform 1 0 2676 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1680363874
transform 1 0 2684 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1680363874
transform 1 0 2700 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1680363874
transform 1 0 2596 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_507
timestamp 1680363874
transform 1 0 2644 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1680363874
transform 1 0 2684 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1680363874
transform 1 0 2692 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_551
timestamp 1680363874
transform 1 0 2596 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1680363874
transform 1 0 2724 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1680363874
transform 1 0 2756 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1680363874
transform 1 0 2796 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1680363874
transform 1 0 2852 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1680363874
transform 1 0 2772 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_552
timestamp 1680363874
transform 1 0 2772 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1680363874
transform 1 0 2788 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_506
timestamp 1680363874
transform 1 0 2868 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_508
timestamp 1680363874
transform 1 0 2868 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1680363874
transform 1 0 2924 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_507
timestamp 1680363874
transform 1 0 2916 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1680363874
transform 1 0 2932 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1680363874
transform 1 0 2908 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1680363874
transform 1 0 2924 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1680363874
transform 1 0 2932 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1680363874
transform 1 0 2964 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1680363874
transform 1 0 2964 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1680363874
transform 1 0 2956 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1680363874
transform 1 0 2996 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1680363874
transform 1 0 3076 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1680363874
transform 1 0 3124 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1680363874
transform 1 0 3116 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1680363874
transform 1 0 3148 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_509
timestamp 1680363874
transform 1 0 2956 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1680363874
transform 1 0 2964 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1680363874
transform 1 0 2996 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1680363874
transform 1 0 3060 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1680363874
transform 1 0 3092 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1680363874
transform 1 0 3044 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1680363874
transform 1 0 3140 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_365
timestamp 1680363874
transform 1 0 3164 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_514
timestamp 1680363874
transform 1 0 3164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1680363874
transform 1 0 3188 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1680363874
transform 1 0 3236 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_515
timestamp 1680363874
transform 1 0 3220 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1680363874
transform 1 0 3212 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1680363874
transform 1 0 3244 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1680363874
transform 1 0 3260 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1680363874
transform 1 0 3268 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_518
timestamp 1680363874
transform 1 0 3276 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1680363874
transform 1 0 3284 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1680363874
transform 1 0 3236 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1680363874
transform 1 0 3244 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1680363874
transform 1 0 3268 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1680363874
transform 1 0 3276 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_554
timestamp 1680363874
transform 1 0 3260 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1680363874
transform 1 0 3300 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1680363874
transform 1 0 3308 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1680363874
transform 1 0 3300 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_651
timestamp 1680363874
transform 1 0 3316 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_423
timestamp 1680363874
transform 1 0 3340 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1680363874
transform 1 0 3364 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1680363874
transform 1 0 3332 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1680363874
transform 1 0 3332 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1680363874
transform 1 0 3348 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1680363874
transform 1 0 3364 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1680363874
transform 1 0 3332 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_652
timestamp 1680363874
transform 1 0 3356 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_488
timestamp 1680363874
transform 1 0 3372 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1680363874
transform 1 0 3388 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1680363874
transform 1 0 3484 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1680363874
transform 1 0 3444 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1680363874
transform 1 0 3428 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_524
timestamp 1680363874
transform 1 0 3428 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1680363874
transform 1 0 3476 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_653
timestamp 1680363874
transform 1 0 3476 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_490
timestamp 1680363874
transform 1 0 3500 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_654
timestamp 1680363874
transform 1 0 3500 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1680363874
transform 1 0 3556 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1680363874
transform 1 0 3548 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_525
timestamp 1680363874
transform 1 0 3524 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1680363874
transform 1 0 3540 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1680363874
transform 1 0 3556 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_555
timestamp 1680363874
transform 1 0 3516 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_655
timestamp 1680363874
transform 1 0 3548 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1680363874
transform 1 0 3556 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_556
timestamp 1680363874
transform 1 0 3540 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1680363874
transform 1 0 3596 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1680363874
transform 1 0 3652 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1680363874
transform 1 0 3588 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1680363874
transform 1 0 3628 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1680363874
transform 1 0 3588 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1680363874
transform 1 0 3596 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1680363874
transform 1 0 3628 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1680363874
transform 1 0 3676 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1680363874
transform 1 0 3700 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_367
timestamp 1680363874
transform 1 0 3756 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1680363874
transform 1 0 3732 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1680363874
transform 1 0 3772 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1680363874
transform 1 0 3732 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1680363874
transform 1 0 3740 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1680363874
transform 1 0 3772 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1680363874
transform 1 0 3724 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1680363874
transform 1 0 3772 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_659
timestamp 1680363874
transform 1 0 3820 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_557
timestamp 1680363874
transform 1 0 3796 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1680363874
transform 1 0 3836 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_534
timestamp 1680363874
transform 1 0 3836 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1680363874
transform 1 0 3836 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_558
timestamp 1680363874
transform 1 0 3836 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_535
timestamp 1680363874
transform 1 0 3876 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_491
timestamp 1680363874
transform 1 0 3884 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1680363874
transform 1 0 3900 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1680363874
transform 1 0 3900 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1680363874
transform 1 0 3884 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1680363874
transform 1 0 3892 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1680363874
transform 1 0 3948 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1680363874
transform 1 0 3956 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_663
timestamp 1680363874
transform 1 0 3940 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1680363874
transform 1 0 3956 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1680363874
transform 1 0 3964 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1680363874
transform 1 0 3980 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_397
timestamp 1680363874
transform 1 0 4028 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1680363874
transform 1 0 4036 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_539
timestamp 1680363874
transform 1 0 4028 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1680363874
transform 1 0 4036 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1680363874
transform 1 0 4044 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_540
timestamp 1680363874
transform 1 0 4044 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1680363874
transform 1 0 4060 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_540
timestamp 1680363874
transform 1 0 4084 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1680363874
transform 1 0 4100 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1680363874
transform 1 0 4076 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_493
timestamp 1680363874
transform 1 0 4108 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_669
timestamp 1680363874
transform 1 0 4108 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1680363874
transform 1 0 4116 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1680363874
transform 1 0 4140 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1680363874
transform 1 0 4132 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1680363874
transform 1 0 4132 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1680363874
transform 1 0 4140 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1680363874
transform 1 0 4140 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1680363874
transform 1 0 4180 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1680363874
transform 1 0 4164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1680363874
transform 1 0 4180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1680363874
transform 1 0 4148 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1680363874
transform 1 0 4172 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_373
timestamp 1680363874
transform 1 0 4268 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1680363874
transform 1 0 4260 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1680363874
transform 1 0 4196 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1680363874
transform 1 0 4236 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_546
timestamp 1680363874
transform 1 0 4228 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_494
timestamp 1680363874
transform 1 0 4252 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1680363874
transform 1 0 4276 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_495
timestamp 1680363874
transform 1 0 4340 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_547
timestamp 1680363874
transform 1 0 4348 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_514
timestamp 1680363874
transform 1 0 4332 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1680363874
transform 1 0 4380 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1680363874
transform 1 0 4404 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_548
timestamp 1680363874
transform 1 0 4396 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1680363874
transform 1 0 4420 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1680363874
transform 1 0 4460 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1680363874
transform 1 0 4484 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1680363874
transform 1 0 4428 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1680363874
transform 1 0 4452 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1680363874
transform 1 0 4468 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_498
timestamp 1680363874
transform 1 0 4476 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_552
timestamp 1680363874
transform 1 0 4484 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1680363874
transform 1 0 4412 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1680363874
transform 1 0 4420 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1680363874
transform 1 0 4436 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1680363874
transform 1 0 4444 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1680363874
transform 1 0 4460 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1680363874
transform 1 0 4476 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1680363874
transform 1 0 4484 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1680363874
transform 1 0 4444 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1680363874
transform 1 0 4548 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1680363874
transform 1 0 4548 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_374
timestamp 1680363874
transform 1 0 4564 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1680363874
transform 1 0 4604 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1680363874
transform 1 0 4596 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1680363874
transform 1 0 4588 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_553
timestamp 1680363874
transform 1 0 4556 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1680363874
transform 1 0 4564 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1680363874
transform 1 0 4580 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1680363874
transform 1 0 4596 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1680363874
transform 1 0 4572 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1680363874
transform 1 0 4588 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1680363874
transform 1 0 4596 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1680363874
transform 1 0 4564 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1680363874
transform 1 0 4644 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1680363874
transform 1 0 4636 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1680363874
transform 1 0 4676 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_557
timestamp 1680363874
transform 1 0 4636 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1680363874
transform 1 0 4644 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_499
timestamp 1680363874
transform 1 0 4660 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_559
timestamp 1680363874
transform 1 0 4676 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1680363874
transform 1 0 4724 0 1 4405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_6
timestamp 1680363874
transform 1 0 48 0 1 4370
box -10 -3 10 3
use M3_M2  M3_M2_559
timestamp 1680363874
transform 1 0 76 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1680363874
transform 1 0 172 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1680363874
transform 1 0 188 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_47
timestamp 1680363874
transform -1 0 168 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_37
timestamp 1680363874
transform 1 0 168 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1680363874
transform 1 0 184 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_38
timestamp 1680363874
transform 1 0 280 0 1 4370
box -9 -3 26 105
use FILL  FILL_322
timestamp 1680363874
transform 1 0 296 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1680363874
transform 1 0 304 0 1 4370
box -8 -3 104 105
use FILL  FILL_323
timestamp 1680363874
transform 1 0 400 0 1 4370
box -8 -3 16 105
use FILL  FILL_330
timestamp 1680363874
transform 1 0 408 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_40
timestamp 1680363874
transform 1 0 416 0 1 4370
box -9 -3 26 105
use FILL  FILL_332
timestamp 1680363874
transform 1 0 432 0 1 4370
box -8 -3 16 105
use FILL  FILL_334
timestamp 1680363874
transform 1 0 440 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_25
timestamp 1680363874
transform 1 0 448 0 1 4370
box -8 -3 46 105
use FILL  FILL_336
timestamp 1680363874
transform 1 0 488 0 1 4370
box -8 -3 16 105
use FILL  FILL_337
timestamp 1680363874
transform 1 0 496 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1680363874
transform 1 0 504 0 1 4370
box -9 -3 26 105
use FILL  FILL_338
timestamp 1680363874
transform 1 0 520 0 1 4370
box -8 -3 16 105
use FILL  FILL_339
timestamp 1680363874
transform 1 0 528 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_26
timestamp 1680363874
transform 1 0 536 0 1 4370
box -8 -3 46 105
use FILL  FILL_340
timestamp 1680363874
transform 1 0 576 0 1 4370
box -8 -3 16 105
use FILL  FILL_341
timestamp 1680363874
transform 1 0 584 0 1 4370
box -8 -3 16 105
use FILL  FILL_342
timestamp 1680363874
transform 1 0 592 0 1 4370
box -8 -3 16 105
use FILL  FILL_343
timestamp 1680363874
transform 1 0 600 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_28
timestamp 1680363874
transform 1 0 608 0 1 4370
box -8 -3 46 105
use FILL  FILL_347
timestamp 1680363874
transform 1 0 648 0 1 4370
box -8 -3 16 105
use FILL  FILL_349
timestamp 1680363874
transform 1 0 656 0 1 4370
box -8 -3 16 105
use FILL  FILL_351
timestamp 1680363874
transform 1 0 664 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_562
timestamp 1680363874
transform 1 0 708 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_30
timestamp 1680363874
transform 1 0 672 0 1 4370
box -8 -3 46 105
use FILL  FILL_352
timestamp 1680363874
transform 1 0 712 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_563
timestamp 1680363874
transform 1 0 748 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_32
timestamp 1680363874
transform 1 0 720 0 1 4370
box -8 -3 46 105
use OAI21X1  OAI21X1_3
timestamp 1680363874
transform 1 0 760 0 1 4370
box -8 -3 34 105
use FILL  FILL_360
timestamp 1680363874
transform 1 0 792 0 1 4370
box -8 -3 16 105
use FILL  FILL_362
timestamp 1680363874
transform 1 0 800 0 1 4370
box -8 -3 16 105
use FILL  FILL_364
timestamp 1680363874
transform 1 0 808 0 1 4370
box -8 -3 16 105
use FILL  FILL_366
timestamp 1680363874
transform 1 0 816 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1680363874
transform 1 0 824 0 1 4370
box -8 -3 34 105
use FILL  FILL_368
timestamp 1680363874
transform 1 0 856 0 1 4370
box -8 -3 16 105
use FILL  FILL_370
timestamp 1680363874
transform 1 0 864 0 1 4370
box -8 -3 16 105
use FILL  FILL_372
timestamp 1680363874
transform 1 0 872 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_7
timestamp 1680363874
transform -1 0 912 0 1 4370
box -8 -3 34 105
use FILL  FILL_373
timestamp 1680363874
transform 1 0 912 0 1 4370
box -8 -3 16 105
use FILL  FILL_374
timestamp 1680363874
transform 1 0 920 0 1 4370
box -8 -3 16 105
use FILL  FILL_378
timestamp 1680363874
transform 1 0 928 0 1 4370
box -8 -3 16 105
use FILL  FILL_380
timestamp 1680363874
transform 1 0 936 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1680363874
transform 1 0 944 0 1 4370
box -8 -3 34 105
use OAI22X1  OAI22X1_33
timestamp 1680363874
transform -1 0 1016 0 1 4370
box -8 -3 46 105
use FILL  FILL_382
timestamp 1680363874
transform 1 0 1016 0 1 4370
box -8 -3 16 105
use FILL  FILL_383
timestamp 1680363874
transform 1 0 1024 0 1 4370
box -8 -3 16 105
use FILL  FILL_384
timestamp 1680363874
transform 1 0 1032 0 1 4370
box -8 -3 16 105
use FILL  FILL_385
timestamp 1680363874
transform 1 0 1040 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_34
timestamp 1680363874
transform 1 0 1048 0 1 4370
box -8 -3 46 105
use FILL  FILL_386
timestamp 1680363874
transform 1 0 1088 0 1 4370
box -8 -3 16 105
use FILL  FILL_387
timestamp 1680363874
transform 1 0 1096 0 1 4370
box -8 -3 16 105
use FILL  FILL_388
timestamp 1680363874
transform 1 0 1104 0 1 4370
box -8 -3 16 105
use FILL  FILL_389
timestamp 1680363874
transform 1 0 1112 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_38
timestamp 1680363874
transform 1 0 1120 0 1 4370
box -8 -3 46 105
use FILL  FILL_397
timestamp 1680363874
transform 1 0 1160 0 1 4370
box -8 -3 16 105
use FILL  FILL_404
timestamp 1680363874
transform 1 0 1168 0 1 4370
box -8 -3 16 105
use FILL  FILL_406
timestamp 1680363874
transform 1 0 1176 0 1 4370
box -8 -3 16 105
use FILL  FILL_407
timestamp 1680363874
transform 1 0 1184 0 1 4370
box -8 -3 16 105
use FILL  FILL_408
timestamp 1680363874
transform 1 0 1192 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1680363874
transform -1 0 1216 0 1 4370
box -9 -3 26 105
use FILL  FILL_409
timestamp 1680363874
transform 1 0 1216 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_39
timestamp 1680363874
transform 1 0 1224 0 1 4370
box -8 -3 46 105
use FILL  FILL_414
timestamp 1680363874
transform 1 0 1264 0 1 4370
box -8 -3 16 105
use FILL  FILL_421
timestamp 1680363874
transform 1 0 1272 0 1 4370
box -8 -3 16 105
use FILL  FILL_422
timestamp 1680363874
transform 1 0 1280 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1680363874
transform -1 0 1384 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_45
timestamp 1680363874
transform -1 0 1400 0 1 4370
box -9 -3 26 105
use FILL  FILL_423
timestamp 1680363874
transform 1 0 1400 0 1 4370
box -8 -3 16 105
use FILL  FILL_431
timestamp 1680363874
transform 1 0 1408 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_42
timestamp 1680363874
transform 1 0 1416 0 1 4370
box -8 -3 46 105
use INVX2  INVX2_46
timestamp 1680363874
transform -1 0 1472 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1680363874
transform 1 0 1472 0 1 4370
box -8 -3 104 105
use FILL  FILL_433
timestamp 1680363874
transform 1 0 1568 0 1 4370
box -8 -3 16 105
use FILL  FILL_442
timestamp 1680363874
transform 1 0 1576 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_47
timestamp 1680363874
transform -1 0 1600 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1680363874
transform 1 0 1600 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_48
timestamp 1680363874
transform -1 0 1712 0 1 4370
box -9 -3 26 105
use FILL  FILL_443
timestamp 1680363874
transform 1 0 1712 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_19
timestamp 1680363874
transform -1 0 1760 0 1 4370
box -8 -3 46 105
use FILL  FILL_444
timestamp 1680363874
transform 1 0 1760 0 1 4370
box -8 -3 16 105
use FILL  FILL_453
timestamp 1680363874
transform 1 0 1768 0 1 4370
box -8 -3 16 105
use FILL  FILL_454
timestamp 1680363874
transform 1 0 1776 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_43
timestamp 1680363874
transform -1 0 1824 0 1 4370
box -8 -3 46 105
use FILL  FILL_455
timestamp 1680363874
transform 1 0 1824 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_44
timestamp 1680363874
transform -1 0 1872 0 1 4370
box -8 -3 46 105
use FILL  FILL_456
timestamp 1680363874
transform 1 0 1872 0 1 4370
box -8 -3 16 105
use FILL  FILL_457
timestamp 1680363874
transform 1 0 1880 0 1 4370
box -8 -3 16 105
use FILL  FILL_458
timestamp 1680363874
transform 1 0 1888 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_51
timestamp 1680363874
transform -1 0 1912 0 1 4370
box -9 -3 26 105
use FILL  FILL_459
timestamp 1680363874
transform 1 0 1912 0 1 4370
box -8 -3 16 105
use FILL  FILL_460
timestamp 1680363874
transform 1 0 1920 0 1 4370
box -8 -3 16 105
use FILL  FILL_461
timestamp 1680363874
transform 1 0 1928 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_20
timestamp 1680363874
transform 1 0 1936 0 1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1680363874
transform 1 0 1976 0 1 4370
box -8 -3 104 105
use FILL  FILL_462
timestamp 1680363874
transform 1 0 2072 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_564
timestamp 1680363874
transform 1 0 2092 0 1 4375
box -3 -3 3 3
use AOI22X1  AOI22X1_21
timestamp 1680363874
transform -1 0 2120 0 1 4370
box -8 -3 46 105
use FILL  FILL_463
timestamp 1680363874
transform 1 0 2120 0 1 4370
box -8 -3 16 105
use FILL  FILL_464
timestamp 1680363874
transform 1 0 2128 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_565
timestamp 1680363874
transform 1 0 2156 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_59
timestamp 1680363874
transform 1 0 2136 0 1 4370
box -8 -3 104 105
use FILL  FILL_465
timestamp 1680363874
transform 1 0 2232 0 1 4370
box -8 -3 16 105
use FILL  FILL_466
timestamp 1680363874
transform 1 0 2240 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_52
timestamp 1680363874
transform 1 0 2248 0 1 4370
box -9 -3 26 105
use FILL  FILL_467
timestamp 1680363874
transform 1 0 2264 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1680363874
transform 1 0 2272 0 1 4370
box -8 -3 104 105
use FILL  FILL_468
timestamp 1680363874
transform 1 0 2368 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_45
timestamp 1680363874
transform 1 0 2376 0 1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1680363874
transform 1 0 2416 0 1 4370
box -8 -3 104 105
use FILL  FILL_469
timestamp 1680363874
transform 1 0 2512 0 1 4370
box -8 -3 16 105
use FILL  FILL_470
timestamp 1680363874
transform 1 0 2520 0 1 4370
box -8 -3 16 105
use FILL  FILL_471
timestamp 1680363874
transform 1 0 2528 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1680363874
transform -1 0 2552 0 1 4370
box -9 -3 26 105
use FILL  FILL_472
timestamp 1680363874
transform 1 0 2552 0 1 4370
box -8 -3 16 105
use FILL  FILL_473
timestamp 1680363874
transform 1 0 2560 0 1 4370
box -8 -3 16 105
use FILL  FILL_474
timestamp 1680363874
transform 1 0 2568 0 1 4370
box -8 -3 16 105
use FILL  FILL_502
timestamp 1680363874
transform 1 0 2576 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1680363874
transform 1 0 2584 0 1 4370
box -8 -3 104 105
use AOI22X1  AOI22X1_26
timestamp 1680363874
transform 1 0 2680 0 1 4370
box -8 -3 46 105
use FILL  FILL_509
timestamp 1680363874
transform 1 0 2720 0 1 4370
box -8 -3 16 105
use FILL  FILL_510
timestamp 1680363874
transform 1 0 2728 0 1 4370
box -8 -3 16 105
use FILL  FILL_511
timestamp 1680363874
transform 1 0 2736 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_566
timestamp 1680363874
transform 1 0 2756 0 1 4375
box -3 -3 3 3
use FILL  FILL_512
timestamp 1680363874
transform 1 0 2744 0 1 4370
box -8 -3 16 105
use FILL  FILL_513
timestamp 1680363874
transform 1 0 2752 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_567
timestamp 1680363874
transform 1 0 2828 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1680363874
transform 1 0 2852 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_66
timestamp 1680363874
transform 1 0 2760 0 1 4370
box -8 -3 104 105
use FILL  FILL_514
timestamp 1680363874
transform 1 0 2856 0 1 4370
box -8 -3 16 105
use FILL  FILL_515
timestamp 1680363874
transform 1 0 2864 0 1 4370
box -8 -3 16 105
use FILL  FILL_516
timestamp 1680363874
transform 1 0 2872 0 1 4370
box -8 -3 16 105
use FILL  FILL_517
timestamp 1680363874
transform 1 0 2880 0 1 4370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1680363874
transform 1 0 2888 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_29
timestamp 1680363874
transform 1 0 2896 0 1 4370
box -8 -3 46 105
use FILL  FILL_519
timestamp 1680363874
transform 1 0 2936 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_59
timestamp 1680363874
transform 1 0 2944 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1680363874
transform -1 0 3056 0 1 4370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1680363874
transform -1 0 3152 0 1 4370
box -8 -3 104 105
use FILL  FILL_520
timestamp 1680363874
transform 1 0 3152 0 1 4370
box -8 -3 16 105
use FILL  FILL_521
timestamp 1680363874
transform 1 0 3160 0 1 4370
box -8 -3 16 105
use FILL  FILL_522
timestamp 1680363874
transform 1 0 3168 0 1 4370
box -8 -3 16 105
use FILL  FILL_523
timestamp 1680363874
transform 1 0 3176 0 1 4370
box -8 -3 16 105
use FILL  FILL_524
timestamp 1680363874
transform 1 0 3184 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_48
timestamp 1680363874
transform 1 0 3192 0 1 4370
box -8 -3 46 105
use FILL  FILL_525
timestamp 1680363874
transform 1 0 3232 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_30
timestamp 1680363874
transform -1 0 3280 0 1 4370
box -8 -3 46 105
use INVX2  INVX2_60
timestamp 1680363874
transform 1 0 3280 0 1 4370
box -9 -3 26 105
use FILL  FILL_526
timestamp 1680363874
transform 1 0 3296 0 1 4370
box -8 -3 16 105
use FILL  FILL_527
timestamp 1680363874
transform 1 0 3304 0 1 4370
box -8 -3 16 105
use FILL  FILL_546
timestamp 1680363874
transform 1 0 3312 0 1 4370
box -8 -3 16 105
use FILL  FILL_548
timestamp 1680363874
transform 1 0 3320 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_33
timestamp 1680363874
transform 1 0 3328 0 1 4370
box -8 -3 46 105
use FILL  FILL_549
timestamp 1680363874
transform 1 0 3368 0 1 4370
box -8 -3 16 105
use FILL  FILL_550
timestamp 1680363874
transform 1 0 3376 0 1 4370
box -8 -3 16 105
use FILL  FILL_551
timestamp 1680363874
transform 1 0 3384 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_569
timestamp 1680363874
transform 1 0 3476 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_71
timestamp 1680363874
transform -1 0 3488 0 1 4370
box -8 -3 104 105
use FILL  FILL_552
timestamp 1680363874
transform 1 0 3488 0 1 4370
box -8 -3 16 105
use FILL  FILL_558
timestamp 1680363874
transform 1 0 3496 0 1 4370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1680363874
transform 1 0 3504 0 1 4370
box -8 -3 16 105
use FILL  FILL_560
timestamp 1680363874
transform 1 0 3512 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_34
timestamp 1680363874
transform 1 0 3520 0 1 4370
box -8 -3 46 105
use FILL  FILL_561
timestamp 1680363874
transform 1 0 3560 0 1 4370
box -8 -3 16 105
use FILL  FILL_562
timestamp 1680363874
transform 1 0 3568 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_62
timestamp 1680363874
transform 1 0 3576 0 1 4370
box -9 -3 26 105
use M3_M2  M3_M2_570
timestamp 1680363874
transform 1 0 3676 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_73
timestamp 1680363874
transform -1 0 3688 0 1 4370
box -8 -3 104 105
use FILL  FILL_563
timestamp 1680363874
transform 1 0 3688 0 1 4370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1680363874
transform 1 0 3696 0 1 4370
box -8 -3 16 105
use FILL  FILL_565
timestamp 1680363874
transform 1 0 3704 0 1 4370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1680363874
transform 1 0 3712 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_63
timestamp 1680363874
transform 1 0 3720 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1680363874
transform -1 0 3832 0 1 4370
box -8 -3 104 105
use FILL  FILL_567
timestamp 1680363874
transform 1 0 3832 0 1 4370
box -8 -3 16 105
use FILL  FILL_568
timestamp 1680363874
transform 1 0 3840 0 1 4370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1680363874
transform 1 0 3848 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_35
timestamp 1680363874
transform -1 0 3896 0 1 4370
box -8 -3 46 105
use FILL  FILL_570
timestamp 1680363874
transform 1 0 3896 0 1 4370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1680363874
transform 1 0 3904 0 1 4370
box -8 -3 16 105
use FILL  FILL_572
timestamp 1680363874
transform 1 0 3912 0 1 4370
box -8 -3 16 105
use FILL  FILL_583
timestamp 1680363874
transform 1 0 3920 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_38
timestamp 1680363874
transform -1 0 3968 0 1 4370
box -8 -3 46 105
use FILL  FILL_584
timestamp 1680363874
transform 1 0 3968 0 1 4370
box -8 -3 16 105
use FILL  FILL_592
timestamp 1680363874
transform 1 0 3976 0 1 4370
box -8 -3 16 105
use FILL  FILL_594
timestamp 1680363874
transform 1 0 3984 0 1 4370
box -8 -3 16 105
use FILL  FILL_595
timestamp 1680363874
transform 1 0 3992 0 1 4370
box -8 -3 16 105
use FILL  FILL_596
timestamp 1680363874
transform 1 0 4000 0 1 4370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1680363874
transform 1 0 4008 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_571
timestamp 1680363874
transform 1 0 4028 0 1 4375
box -3 -3 3 3
use INVX2  INVX2_67
timestamp 1680363874
transform -1 0 4032 0 1 4370
box -9 -3 26 105
use FILL  FILL_599
timestamp 1680363874
transform 1 0 4032 0 1 4370
box -8 -3 16 105
use FILL  FILL_600
timestamp 1680363874
transform 1 0 4040 0 1 4370
box -8 -3 16 105
use FILL  FILL_601
timestamp 1680363874
transform 1 0 4048 0 1 4370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1680363874
transform 1 0 4056 0 1 4370
box -8 -3 16 105
use FILL  FILL_603
timestamp 1680363874
transform 1 0 4064 0 1 4370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1680363874
transform 1 0 4072 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_572
timestamp 1680363874
transform 1 0 4124 0 1 4375
box -3 -3 3 3
use AOI22X1  AOI22X1_39
timestamp 1680363874
transform -1 0 4120 0 1 4370
box -8 -3 46 105
use FILL  FILL_605
timestamp 1680363874
transform 1 0 4120 0 1 4370
box -8 -3 16 105
use FILL  FILL_606
timestamp 1680363874
transform 1 0 4128 0 1 4370
box -8 -3 16 105
use FILL  FILL_607
timestamp 1680363874
transform 1 0 4136 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_41
timestamp 1680363874
transform 1 0 4144 0 1 4370
box -8 -3 46 105
use FILL  FILL_615
timestamp 1680363874
transform 1 0 4184 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1680363874
transform -1 0 4288 0 1 4370
box -8 -3 104 105
use FILL  FILL_616
timestamp 1680363874
transform 1 0 4288 0 1 4370
box -8 -3 16 105
use FILL  FILL_631
timestamp 1680363874
transform 1 0 4296 0 1 4370
box -8 -3 16 105
use FILL  FILL_632
timestamp 1680363874
transform 1 0 4304 0 1 4370
box -8 -3 16 105
use FILL  FILL_633
timestamp 1680363874
transform 1 0 4312 0 1 4370
box -8 -3 16 105
use FILL  FILL_634
timestamp 1680363874
transform 1 0 4320 0 1 4370
box -8 -3 16 105
use FILL  FILL_635
timestamp 1680363874
transform 1 0 4328 0 1 4370
box -8 -3 16 105
use FILL  FILL_636
timestamp 1680363874
transform 1 0 4336 0 1 4370
box -8 -3 16 105
use FILL  FILL_638
timestamp 1680363874
transform 1 0 4344 0 1 4370
box -8 -3 16 105
use FILL  FILL_639
timestamp 1680363874
transform 1 0 4352 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_68
timestamp 1680363874
transform -1 0 4376 0 1 4370
box -9 -3 26 105
use FILL  FILL_640
timestamp 1680363874
transform 1 0 4376 0 1 4370
box -8 -3 16 105
use FILL  FILL_641
timestamp 1680363874
transform 1 0 4384 0 1 4370
box -8 -3 16 105
use FILL  FILL_643
timestamp 1680363874
transform 1 0 4392 0 1 4370
box -8 -3 16 105
use FILL  FILL_645
timestamp 1680363874
transform 1 0 4400 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1680363874
transform -1 0 4448 0 1 4370
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1680363874
transform 1 0 4448 0 1 4370
box -8 -3 46 105
use FILL  FILL_646
timestamp 1680363874
transform 1 0 4488 0 1 4370
box -8 -3 16 105
use FILL  FILL_647
timestamp 1680363874
transform 1 0 4496 0 1 4370
box -8 -3 16 105
use FILL  FILL_648
timestamp 1680363874
transform 1 0 4504 0 1 4370
box -8 -3 16 105
use FILL  FILL_649
timestamp 1680363874
transform 1 0 4512 0 1 4370
box -8 -3 16 105
use FILL  FILL_650
timestamp 1680363874
transform 1 0 4520 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1680363874
transform 1 0 4528 0 1 4370
box -9 -3 26 105
use FILL  FILL_651
timestamp 1680363874
transform 1 0 4544 0 1 4370
box -8 -3 16 105
use FILL  FILL_657
timestamp 1680363874
transform 1 0 4552 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_44
timestamp 1680363874
transform 1 0 4560 0 1 4370
box -8 -3 46 105
use FILL  FILL_658
timestamp 1680363874
transform 1 0 4600 0 1 4370
box -8 -3 16 105
use FILL  FILL_659
timestamp 1680363874
transform 1 0 4608 0 1 4370
box -8 -3 16 105
use FILL  FILL_660
timestamp 1680363874
transform 1 0 4616 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1680363874
transform 1 0 4624 0 1 4370
box -9 -3 26 105
use M3_M2  M3_M2_573
timestamp 1680363874
transform 1 0 4676 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1680363874
transform 1 0 4724 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_79
timestamp 1680363874
transform -1 0 4736 0 1 4370
box -8 -3 104 105
use FILL  FILL_661
timestamp 1680363874
transform 1 0 4736 0 1 4370
box -8 -3 16 105
use FILL  FILL_662
timestamp 1680363874
transform 1 0 4744 0 1 4370
box -8 -3 16 105
use FILL  FILL_663
timestamp 1680363874
transform 1 0 4752 0 1 4370
box -8 -3 16 105
use FILL  FILL_664
timestamp 1680363874
transform 1 0 4760 0 1 4370
box -8 -3 16 105
use FILL  FILL_665
timestamp 1680363874
transform 1 0 4768 0 1 4370
box -8 -3 16 105
use FILL  FILL_666
timestamp 1680363874
transform 1 0 4776 0 1 4370
box -8 -3 16 105
use FILL  FILL_667
timestamp 1680363874
transform 1 0 4784 0 1 4370
box -8 -3 16 105
use FILL  FILL_668
timestamp 1680363874
transform 1 0 4792 0 1 4370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_7
timestamp 1680363874
transform 1 0 4827 0 1 4370
box -10 -3 10 3
use M3_M2  M3_M2_595
timestamp 1680363874
transform 1 0 172 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1680363874
transform 1 0 132 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1680363874
transform 1 0 116 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1680363874
transform 1 0 188 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_689
timestamp 1680363874
transform 1 0 156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1680363874
transform 1 0 172 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1680363874
transform 1 0 188 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1680363874
transform 1 0 204 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1680363874
transform 1 0 68 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1680363874
transform 1 0 132 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_701
timestamp 1680363874
transform 1 0 132 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_813
timestamp 1680363874
transform 1 0 180 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1680363874
transform 1 0 196 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_702
timestamp 1680363874
transform 1 0 180 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1680363874
transform 1 0 196 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1680363874
transform 1 0 228 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_693
timestamp 1680363874
transform 1 0 220 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_625
timestamp 1680363874
transform 1 0 284 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_694
timestamp 1680363874
transform 1 0 236 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1680363874
transform 1 0 284 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_626
timestamp 1680363874
transform 1 0 372 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_695
timestamp 1680363874
transform 1 0 356 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1680363874
transform 1 0 372 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1680363874
transform 1 0 364 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1680363874
transform 1 0 372 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1680363874
transform 1 0 380 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_703
timestamp 1680363874
transform 1 0 356 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_697
timestamp 1680363874
transform 1 0 396 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1680363874
transform 1 0 404 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_704
timestamp 1680363874
transform 1 0 404 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1680363874
transform 1 0 396 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_818
timestamp 1680363874
transform 1 0 428 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1680363874
transform 1 0 452 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1680363874
transform 1 0 476 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1680363874
transform 1 0 476 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_699
timestamp 1680363874
transform 1 0 476 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1680363874
transform 1 0 492 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1680363874
transform 1 0 468 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_598
timestamp 1680363874
transform 1 0 524 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1680363874
transform 1 0 540 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_701
timestamp 1680363874
transform 1 0 588 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1680363874
transform 1 0 500 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1680363874
transform 1 0 508 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1680363874
transform 1 0 540 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_706
timestamp 1680363874
transform 1 0 492 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1680363874
transform 1 0 468 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1680363874
transform 1 0 588 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1680363874
transform 1 0 588 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_702
timestamp 1680363874
transform 1 0 604 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1680363874
transform 1 0 604 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1680363874
transform 1 0 628 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_703
timestamp 1680363874
transform 1 0 628 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_659
timestamp 1680363874
transform 1 0 636 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1680363874
transform 1 0 644 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1680363874
transform 1 0 652 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1680363874
transform 1 0 620 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1680363874
transform 1 0 636 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1680363874
transform 1 0 612 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1680363874
transform 1 0 636 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1680363874
transform 1 0 620 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1680363874
transform 1 0 652 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1680363874
transform 1 0 684 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_706
timestamp 1680363874
transform 1 0 684 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1680363874
transform 1 0 692 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1680363874
transform 1 0 708 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1680363874
transform 1 0 700 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1680363874
transform 1 0 708 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1680363874
transform 1 0 676 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1680363874
transform 1 0 692 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_600
timestamp 1680363874
transform 1 0 796 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1680363874
transform 1 0 788 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1680363874
transform 1 0 772 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1680363874
transform 1 0 780 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_710
timestamp 1680363874
transform 1 0 796 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1680363874
transform 1 0 796 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_709
timestamp 1680363874
transform 1 0 812 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_946
timestamp 1680363874
transform 1 0 820 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_631
timestamp 1680363874
transform 1 0 844 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1680363874
transform 1 0 836 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_711
timestamp 1680363874
transform 1 0 852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1680363874
transform 1 0 836 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_710
timestamp 1680363874
transform 1 0 852 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_712
timestamp 1680363874
transform 1 0 860 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1680363874
transform 1 0 868 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_632
timestamp 1680363874
transform 1 0 884 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_829
timestamp 1680363874
transform 1 0 892 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_748
timestamp 1680363874
transform 1 0 892 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_713
timestamp 1680363874
transform 1 0 916 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1680363874
transform 1 0 924 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_575
timestamp 1680363874
transform 1 0 964 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1680363874
transform 1 0 972 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1680363874
transform 1 0 972 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_714
timestamp 1680363874
transform 1 0 956 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1680363874
transform 1 0 972 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1680363874
transform 1 0 964 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1680363874
transform 1 0 980 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_711
timestamp 1680363874
transform 1 0 956 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1680363874
transform 1 0 1004 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1680363874
transform 1 0 1004 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1680363874
transform 1 0 1012 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1680363874
transform 1 0 1052 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_716
timestamp 1680363874
transform 1 0 1012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1680363874
transform 1 0 1020 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1680363874
transform 1 0 1036 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1680363874
transform 1 0 1052 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1680363874
transform 1 0 1012 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1680363874
transform 1 0 1028 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_687
timestamp 1680363874
transform 1 0 1036 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1680363874
transform 1 0 1044 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_712
timestamp 1680363874
transform 1 0 1020 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_720
timestamp 1680363874
transform 1 0 1076 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1680363874
transform 1 0 1092 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1680363874
transform 1 0 1076 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1680363874
transform 1 0 1100 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1680363874
transform 1 0 1092 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1680363874
transform 1 0 1116 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1680363874
transform 1 0 1124 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1680363874
transform 1 0 1156 0 1 4345
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1680363874
transform 1 0 1156 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1680363874
transform 1 0 1180 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_723
timestamp 1680363874
transform 1 0 1212 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1680363874
transform 1 0 1244 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_766
timestamp 1680363874
transform 1 0 1252 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1680363874
transform 1 0 1252 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1680363874
transform 1 0 1316 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1680363874
transform 1 0 1300 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_724
timestamp 1680363874
transform 1 0 1284 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1680363874
transform 1 0 1300 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1680363874
transform 1 0 1308 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_726
timestamp 1680363874
transform 1 0 1316 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1680363874
transform 1 0 1324 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_688
timestamp 1680363874
transform 1 0 1284 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_839
timestamp 1680363874
transform 1 0 1292 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1680363874
transform 1 0 1308 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1680363874
transform 1 0 1292 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1680363874
transform 1 0 1324 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1680363874
transform 1 0 1380 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_728
timestamp 1680363874
transform 1 0 1364 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1680363874
transform 1 0 1380 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1680363874
transform 1 0 1356 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_776
timestamp 1680363874
transform 1 0 1356 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1680363874
transform 1 0 1396 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1680363874
transform 1 0 1388 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_580
timestamp 1680363874
transform 1 0 1420 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1680363874
transform 1 0 1452 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1680363874
transform 1 0 1500 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_730
timestamp 1680363874
transform 1 0 1476 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1680363874
transform 1 0 1500 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_713
timestamp 1680363874
transform 1 0 1524 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_844
timestamp 1680363874
transform 1 0 1612 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1680363874
transform 1 0 1628 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1680363874
transform 1 0 1636 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_845
timestamp 1680363874
transform 1 0 1636 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_638
timestamp 1680363874
transform 1 0 1676 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1680363874
transform 1 0 1652 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1680363874
transform 1 0 1700 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1680363874
transform 1 0 1732 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1680363874
transform 1 0 1740 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1680363874
transform 1 0 1748 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_714
timestamp 1680363874
transform 1 0 1700 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1680363874
transform 1 0 1740 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_733
timestamp 1680363874
transform 1 0 1764 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1680363874
transform 1 0 1772 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_639
timestamp 1680363874
transform 1 0 1804 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_735
timestamp 1680363874
transform 1 0 1788 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1680363874
transform 1 0 1804 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1680363874
transform 1 0 1796 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1680363874
transform 1 0 1812 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1680363874
transform 1 0 1828 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1680363874
transform 1 0 1844 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_750
timestamp 1680363874
transform 1 0 1844 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1680363874
transform 1 0 1940 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1680363874
transform 1 0 1940 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1680363874
transform 1 0 1916 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1680363874
transform 1 0 1956 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_716
timestamp 1680363874
transform 1 0 1916 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1680363874
transform 1 0 1956 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_855
timestamp 1680363874
transform 1 0 1972 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1680363874
transform 1 0 1972 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1680363874
transform 1 0 1988 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_739
timestamp 1680363874
transform 1 0 1988 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1680363874
transform 1 0 1996 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1680363874
transform 1 0 2012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1680363874
transform 1 0 2004 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1680363874
transform 1 0 2020 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1680363874
transform 1 0 2028 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1680363874
transform 1 0 2028 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1680363874
transform 1 0 1996 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1680363874
transform 1 0 2044 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1680363874
transform 1 0 2140 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1680363874
transform 1 0 2108 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1680363874
transform 1 0 2140 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1680363874
transform 1 0 2060 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1680363874
transform 1 0 2116 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1680363874
transform 1 0 2156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1680363874
transform 1 0 2180 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1680363874
transform 1 0 2172 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1680363874
transform 1 0 2188 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1680363874
transform 1 0 2204 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_720
timestamp 1680363874
transform 1 0 2204 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_745
timestamp 1680363874
transform 1 0 2220 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1680363874
transform 1 0 2228 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_605
timestamp 1680363874
transform 1 0 2276 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_747
timestamp 1680363874
transform 1 0 2276 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1680363874
transform 1 0 2252 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1680363874
transform 1 0 2268 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1680363874
transform 1 0 2284 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1680363874
transform 1 0 2308 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_585
timestamp 1680363874
transform 1 0 2332 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1680363874
transform 1 0 2356 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1680363874
transform 1 0 2396 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1680363874
transform 1 0 2396 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1680363874
transform 1 0 2412 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_748
timestamp 1680363874
transform 1 0 2372 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1680363874
transform 1 0 2380 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1680363874
transform 1 0 2396 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1680363874
transform 1 0 2404 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1680363874
transform 1 0 2364 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_768
timestamp 1680363874
transform 1 0 2364 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_869
timestamp 1680363874
transform 1 0 2388 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1680363874
transform 1 0 2420 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_777
timestamp 1680363874
transform 1 0 2412 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1680363874
transform 1 0 2436 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_752
timestamp 1680363874
transform 1 0 2436 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1680363874
transform 1 0 2484 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_871
timestamp 1680363874
transform 1 0 2460 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_607
timestamp 1680363874
transform 1 0 2556 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_753
timestamp 1680363874
transform 1 0 2524 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1680363874
transform 1 0 2532 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_754
timestamp 1680363874
transform 1 0 2556 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1680363874
transform 1 0 2524 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1680363874
transform 1 0 2532 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1680363874
transform 1 0 2548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1680363874
transform 1 0 2564 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_752
timestamp 1680363874
transform 1 0 2524 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1680363874
transform 1 0 2532 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1680363874
transform 1 0 2564 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1680363874
transform 1 0 2596 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1680363874
transform 1 0 2604 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1680363874
transform 1 0 2612 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1680363874
transform 1 0 2604 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_876
timestamp 1680363874
transform 1 0 2620 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1680363874
transform 1 0 2652 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1680363874
transform 1 0 2684 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1680363874
transform 1 0 2676 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_756
timestamp 1680363874
transform 1 0 2652 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1680363874
transform 1 0 2660 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1680363874
transform 1 0 2716 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1680363874
transform 1 0 2676 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1680363874
transform 1 0 2684 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1680363874
transform 1 0 2708 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1680363874
transform 1 0 2716 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1680363874
transform 1 0 2644 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1680363874
transform 1 0 2660 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1680363874
transform 1 0 2676 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1680363874
transform 1 0 2684 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1680363874
transform 1 0 2700 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1680363874
transform 1 0 2708 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_882
timestamp 1680363874
transform 1 0 2716 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1680363874
transform 1 0 2676 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1680363874
transform 1 0 2716 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1680363874
transform 1 0 2708 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1680363874
transform 1 0 2788 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1680363874
transform 1 0 2804 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1680363874
transform 1 0 2764 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1680363874
transform 1 0 2748 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1680363874
transform 1 0 2756 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_762
timestamp 1680363874
transform 1 0 2764 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1680363874
transform 1 0 2772 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1680363874
transform 1 0 2788 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_670
timestamp 1680363874
transform 1 0 2796 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_883
timestamp 1680363874
transform 1 0 2740 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1680363874
transform 1 0 2756 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_692
timestamp 1680363874
transform 1 0 2772 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_885
timestamp 1680363874
transform 1 0 2780 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1680363874
transform 1 0 2796 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1680363874
transform 1 0 2740 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1680363874
transform 1 0 2732 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1680363874
transform 1 0 2780 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1680363874
transform 1 0 2820 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1680363874
transform 1 0 2868 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_765
timestamp 1680363874
transform 1 0 2820 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1680363874
transform 1 0 2828 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1680363874
transform 1 0 2844 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_671
timestamp 1680363874
transform 1 0 2852 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_768
timestamp 1680363874
transform 1 0 2860 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1680363874
transform 1 0 2868 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1680363874
transform 1 0 2892 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1680363874
transform 1 0 2900 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1680363874
transform 1 0 2836 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1680363874
transform 1 0 2852 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1680363874
transform 1 0 2868 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1680363874
transform 1 0 2884 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_726
timestamp 1680363874
transform 1 0 2836 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1680363874
transform 1 0 2868 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_891
timestamp 1680363874
transform 1 0 2916 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_754
timestamp 1680363874
transform 1 0 2916 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1680363874
transform 1 0 2964 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1680363874
transform 1 0 2948 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1680363874
transform 1 0 3028 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1680363874
transform 1 0 2940 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1680363874
transform 1 0 2948 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1680363874
transform 1 0 2980 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1680363874
transform 1 0 2940 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1680363874
transform 1 0 2980 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_895
timestamp 1680363874
transform 1 0 3044 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1680363874
transform 1 0 3068 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_773
timestamp 1680363874
transform 1 0 3084 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_673
timestamp 1680363874
transform 1 0 3092 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1680363874
transform 1 0 3100 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1680363874
transform 1 0 3092 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1680363874
transform 1 0 3116 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1680363874
transform 1 0 3180 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_775
timestamp 1680363874
transform 1 0 3156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1680363874
transform 1 0 3172 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1680363874
transform 1 0 3156 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_898
timestamp 1680363874
transform 1 0 3164 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1680363874
transform 1 0 3180 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_674
timestamp 1680363874
transform 1 0 3212 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1680363874
transform 1 0 3244 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1680363874
transform 1 0 3260 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_777
timestamp 1680363874
transform 1 0 3292 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1680363874
transform 1 0 3212 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1680363874
transform 1 0 3268 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_612
timestamp 1680363874
transform 1 0 3316 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1680363874
transform 1 0 3308 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_778
timestamp 1680363874
transform 1 0 3324 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1680363874
transform 1 0 3340 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1680363874
transform 1 0 3356 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1680363874
transform 1 0 3316 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1680363874
transform 1 0 3348 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1680363874
transform 1 0 3324 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1680363874
transform 1 0 3316 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1680363874
transform 1 0 3356 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_904
timestamp 1680363874
transform 1 0 3364 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_730
timestamp 1680363874
transform 1 0 3364 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1680363874
transform 1 0 3460 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_781
timestamp 1680363874
transform 1 0 3460 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1680363874
transform 1 0 3412 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_695
timestamp 1680363874
transform 1 0 3460 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1680363874
transform 1 0 3428 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1680363874
transform 1 0 3476 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_782
timestamp 1680363874
transform 1 0 3476 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1680363874
transform 1 0 3476 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_756
timestamp 1680363874
transform 1 0 3476 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1680363874
transform 1 0 3500 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1680363874
transform 1 0 3524 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1680363874
transform 1 0 3492 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_783
timestamp 1680363874
transform 1 0 3524 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1680363874
transform 1 0 3532 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1680363874
transform 1 0 3500 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1680363874
transform 1 0 3516 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1680363874
transform 1 0 3532 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_757
timestamp 1680363874
transform 1 0 3524 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1680363874
transform 1 0 3636 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1680363874
transform 1 0 3564 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1680363874
transform 1 0 3564 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_785
timestamp 1680363874
transform 1 0 3636 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1680363874
transform 1 0 3548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1680363874
transform 1 0 3556 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1680363874
transform 1 0 3588 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_731
timestamp 1680363874
transform 1 0 3548 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1680363874
transform 1 0 3588 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1680363874
transform 1 0 3604 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1680363874
transform 1 0 3556 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1680363874
transform 1 0 3612 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1680363874
transform 1 0 3620 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1680363874
transform 1 0 3668 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1680363874
transform 1 0 3660 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_786
timestamp 1680363874
transform 1 0 3660 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_678
timestamp 1680363874
transform 1 0 3668 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_913
timestamp 1680363874
transform 1 0 3668 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1680363874
transform 1 0 3700 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1680363874
transform 1 0 3716 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_734
timestamp 1680363874
transform 1 0 3700 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_687
timestamp 1680363874
transform 1 0 3740 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1680363874
transform 1 0 3740 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1680363874
transform 1 0 3756 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_591
timestamp 1680363874
transform 1 0 3876 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1680363874
transform 1 0 3900 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1680363874
transform 1 0 3892 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1680363874
transform 1 0 3836 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1680363874
transform 1 0 3780 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1680363874
transform 1 0 3796 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1680363874
transform 1 0 3884 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1680363874
transform 1 0 3900 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1680363874
transform 1 0 3788 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1680363874
transform 1 0 3804 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1680363874
transform 1 0 3860 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_697
timestamp 1680363874
transform 1 0 3884 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_921
timestamp 1680363874
transform 1 0 3900 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_735
timestamp 1680363874
transform 1 0 3860 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1680363874
transform 1 0 3900 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1680363874
transform 1 0 3948 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1680363874
transform 1 0 3980 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_922
timestamp 1680363874
transform 1 0 3996 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1680363874
transform 1 0 4020 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_679
timestamp 1680363874
transform 1 0 4044 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1680363874
transform 1 0 4052 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1680363874
transform 1 0 4044 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1680363874
transform 1 0 4060 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_737
timestamp 1680363874
transform 1 0 4060 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_794
timestamp 1680363874
transform 1 0 4076 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_618
timestamp 1680363874
transform 1 0 4084 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1680363874
transform 1 0 4116 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1680363874
transform 1 0 4132 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_795
timestamp 1680363874
transform 1 0 4108 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1680363874
transform 1 0 4124 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1680363874
transform 1 0 4148 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1680363874
transform 1 0 4140 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1680363874
transform 1 0 4100 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1680363874
transform 1 0 4116 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1680363874
transform 1 0 4132 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1680363874
transform 1 0 4140 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_760
timestamp 1680363874
transform 1 0 4100 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1680363874
transform 1 0 4140 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1680363874
transform 1 0 4188 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_797
timestamp 1680363874
transform 1 0 4156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1680363874
transform 1 0 4172 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1680363874
transform 1 0 4156 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1680363874
transform 1 0 4180 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1680363874
transform 1 0 4180 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_931
timestamp 1680363874
transform 1 0 4196 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_655
timestamp 1680363874
transform 1 0 4204 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1680363874
transform 1 0 4212 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1680363874
transform 1 0 4236 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_799
timestamp 1680363874
transform 1 0 4244 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1680363874
transform 1 0 4276 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_800
timestamp 1680363874
transform 1 0 4300 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1680363874
transform 1 0 4316 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1680363874
transform 1 0 4332 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1680363874
transform 1 0 4340 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1680363874
transform 1 0 4308 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1680363874
transform 1 0 4324 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_740
timestamp 1680363874
transform 1 0 4308 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1680363874
transform 1 0 4324 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_934
timestamp 1680363874
transform 1 0 4340 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1680363874
transform 1 0 4364 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1680363874
transform 1 0 4372 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_741
timestamp 1680363874
transform 1 0 4340 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1680363874
transform 1 0 4372 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1680363874
transform 1 0 4396 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_805
timestamp 1680363874
transform 1 0 4404 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_681
timestamp 1680363874
transform 1 0 4412 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1680363874
transform 1 0 4452 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1680363874
transform 1 0 4460 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1680363874
transform 1 0 4436 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_682
timestamp 1680363874
transform 1 0 4444 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1680363874
transform 1 0 4460 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1680363874
transform 1 0 4444 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1680363874
transform 1 0 4484 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1680363874
transform 1 0 4540 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_742
timestamp 1680363874
transform 1 0 4444 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1680363874
transform 1 0 4484 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_808
timestamp 1680363874
transform 1 0 4556 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1680363874
transform 1 0 4572 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1680363874
transform 1 0 4676 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1680363874
transform 1 0 4580 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1680363874
transform 1 0 4588 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1680363874
transform 1 0 4596 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_744
timestamp 1680363874
transform 1 0 4580 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1680363874
transform 1 0 4612 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1680363874
transform 1 0 4628 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_699
timestamp 1680363874
transform 1 0 4676 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1680363874
transform 1 0 4628 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_943
timestamp 1680363874
transform 1 0 4692 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1680363874
transform 1 0 4780 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_700
timestamp 1680363874
transform 1 0 4708 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1680363874
transform 1 0 4748 0 1 4325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_8
timestamp 1680363874
transform 1 0 24 0 1 4270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_50
timestamp 1680363874
transform -1 0 168 0 -1 4370
box -8 -3 104 105
use OAI22X1  OAI22X1_23
timestamp 1680363874
transform 1 0 168 0 -1 4370
box -8 -3 46 105
use FILL  FILL_324
timestamp 1680363874
transform 1 0 208 0 -1 4370
box -8 -3 16 105
use FILL  FILL_325
timestamp 1680363874
transform 1 0 216 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1680363874
transform 1 0 224 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_39
timestamp 1680363874
transform 1 0 320 0 -1 4370
box -9 -3 26 105
use FILL  FILL_326
timestamp 1680363874
transform 1 0 336 0 -1 4370
box -8 -3 16 105
use FILL  FILL_327
timestamp 1680363874
transform 1 0 344 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_24
timestamp 1680363874
transform 1 0 352 0 -1 4370
box -8 -3 46 105
use FILL  FILL_328
timestamp 1680363874
transform 1 0 392 0 -1 4370
box -8 -3 16 105
use FILL  FILL_329
timestamp 1680363874
transform 1 0 400 0 -1 4370
box -8 -3 16 105
use FILL  FILL_331
timestamp 1680363874
transform 1 0 408 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_41
timestamp 1680363874
transform 1 0 416 0 -1 4370
box -9 -3 26 105
use FILL  FILL_333
timestamp 1680363874
transform 1 0 432 0 -1 4370
box -8 -3 16 105
use FILL  FILL_335
timestamp 1680363874
transform 1 0 440 0 -1 4370
box -8 -3 16 105
use FILL  FILL_344
timestamp 1680363874
transform 1 0 448 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_27
timestamp 1680363874
transform -1 0 496 0 -1 4370
box -8 -3 46 105
use FILL  FILL_345
timestamp 1680363874
transform 1 0 496 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1680363874
transform -1 0 600 0 -1 4370
box -8 -3 104 105
use FILL  FILL_346
timestamp 1680363874
transform 1 0 600 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_29
timestamp 1680363874
transform 1 0 608 0 -1 4370
box -8 -3 46 105
use FILL  FILL_348
timestamp 1680363874
transform 1 0 648 0 -1 4370
box -8 -3 16 105
use FILL  FILL_350
timestamp 1680363874
transform 1 0 656 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_31
timestamp 1680363874
transform 1 0 664 0 -1 4370
box -8 -3 46 105
use FILL  FILL_353
timestamp 1680363874
transform 1 0 704 0 -1 4370
box -8 -3 16 105
use FILL  FILL_354
timestamp 1680363874
transform 1 0 712 0 -1 4370
box -8 -3 16 105
use FILL  FILL_355
timestamp 1680363874
transform 1 0 720 0 -1 4370
box -8 -3 16 105
use FILL  FILL_356
timestamp 1680363874
transform 1 0 728 0 -1 4370
box -8 -3 16 105
use FILL  FILL_357
timestamp 1680363874
transform 1 0 736 0 -1 4370
box -8 -3 16 105
use FILL  FILL_358
timestamp 1680363874
transform 1 0 744 0 -1 4370
box -8 -3 16 105
use FILL  FILL_359
timestamp 1680363874
transform 1 0 752 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1680363874
transform 1 0 760 0 -1 4370
box -8 -3 34 105
use FILL  FILL_361
timestamp 1680363874
transform 1 0 792 0 -1 4370
box -8 -3 16 105
use FILL  FILL_363
timestamp 1680363874
transform 1 0 800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_365
timestamp 1680363874
transform 1 0 808 0 -1 4370
box -8 -3 16 105
use FILL  FILL_367
timestamp 1680363874
transform 1 0 816 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1680363874
transform 1 0 824 0 -1 4370
box -8 -3 34 105
use FILL  FILL_369
timestamp 1680363874
transform 1 0 856 0 -1 4370
box -8 -3 16 105
use FILL  FILL_371
timestamp 1680363874
transform 1 0 864 0 -1 4370
box -8 -3 16 105
use FILL  FILL_375
timestamp 1680363874
transform 1 0 872 0 -1 4370
box -8 -3 16 105
use FILL  FILL_376
timestamp 1680363874
transform 1 0 880 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1680363874
transform 1 0 888 0 -1 4370
box -8 -3 34 105
use FILL  FILL_377
timestamp 1680363874
transform 1 0 920 0 -1 4370
box -8 -3 16 105
use FILL  FILL_379
timestamp 1680363874
transform 1 0 928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_381
timestamp 1680363874
transform 1 0 936 0 -1 4370
box -8 -3 16 105
use FILL  FILL_390
timestamp 1680363874
transform 1 0 944 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_35
timestamp 1680363874
transform 1 0 952 0 -1 4370
box -8 -3 46 105
use FILL  FILL_391
timestamp 1680363874
transform 1 0 992 0 -1 4370
box -8 -3 16 105
use FILL  FILL_392
timestamp 1680363874
transform 1 0 1000 0 -1 4370
box -8 -3 16 105
use FILL  FILL_393
timestamp 1680363874
transform 1 0 1008 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_36
timestamp 1680363874
transform 1 0 1016 0 -1 4370
box -8 -3 46 105
use FILL  FILL_394
timestamp 1680363874
transform 1 0 1056 0 -1 4370
box -8 -3 16 105
use FILL  FILL_395
timestamp 1680363874
transform 1 0 1064 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_37
timestamp 1680363874
transform 1 0 1072 0 -1 4370
box -8 -3 46 105
use FILL  FILL_396
timestamp 1680363874
transform 1 0 1112 0 -1 4370
box -8 -3 16 105
use FILL  FILL_398
timestamp 1680363874
transform 1 0 1120 0 -1 4370
box -8 -3 16 105
use FILL  FILL_399
timestamp 1680363874
transform 1 0 1128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_400
timestamp 1680363874
transform 1 0 1136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_401
timestamp 1680363874
transform 1 0 1144 0 -1 4370
box -8 -3 16 105
use FILL  FILL_402
timestamp 1680363874
transform 1 0 1152 0 -1 4370
box -8 -3 16 105
use FILL  FILL_403
timestamp 1680363874
transform 1 0 1160 0 -1 4370
box -8 -3 16 105
use FILL  FILL_405
timestamp 1680363874
transform 1 0 1168 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1680363874
transform 1 0 1176 0 -1 4370
box -9 -3 26 105
use FILL  FILL_410
timestamp 1680363874
transform 1 0 1192 0 -1 4370
box -8 -3 16 105
use FILL  FILL_411
timestamp 1680363874
transform 1 0 1200 0 -1 4370
box -8 -3 16 105
use FILL  FILL_412
timestamp 1680363874
transform 1 0 1208 0 -1 4370
box -8 -3 16 105
use FILL  FILL_413
timestamp 1680363874
transform 1 0 1216 0 -1 4370
box -8 -3 16 105
use FILL  FILL_415
timestamp 1680363874
transform 1 0 1224 0 -1 4370
box -8 -3 16 105
use FILL  FILL_416
timestamp 1680363874
transform 1 0 1232 0 -1 4370
box -8 -3 16 105
use FILL  FILL_417
timestamp 1680363874
transform 1 0 1240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_418
timestamp 1680363874
transform 1 0 1248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_419
timestamp 1680363874
transform 1 0 1256 0 -1 4370
box -8 -3 16 105
use FILL  FILL_420
timestamp 1680363874
transform 1 0 1264 0 -1 4370
box -8 -3 16 105
use FILL  FILL_424
timestamp 1680363874
transform 1 0 1272 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_40
timestamp 1680363874
transform -1 0 1320 0 -1 4370
box -8 -3 46 105
use FILL  FILL_425
timestamp 1680363874
transform 1 0 1320 0 -1 4370
box -8 -3 16 105
use FILL  FILL_426
timestamp 1680363874
transform 1 0 1328 0 -1 4370
box -8 -3 16 105
use FILL  FILL_427
timestamp 1680363874
transform 1 0 1336 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_41
timestamp 1680363874
transform -1 0 1384 0 -1 4370
box -8 -3 46 105
use FILL  FILL_428
timestamp 1680363874
transform 1 0 1384 0 -1 4370
box -8 -3 16 105
use FILL  FILL_429
timestamp 1680363874
transform 1 0 1392 0 -1 4370
box -8 -3 16 105
use FILL  FILL_430
timestamp 1680363874
transform 1 0 1400 0 -1 4370
box -8 -3 16 105
use FILL  FILL_432
timestamp 1680363874
transform 1 0 1408 0 -1 4370
box -8 -3 16 105
use FILL  FILL_434
timestamp 1680363874
transform 1 0 1416 0 -1 4370
box -8 -3 16 105
use FILL  FILL_435
timestamp 1680363874
transform 1 0 1424 0 -1 4370
box -8 -3 16 105
use FILL  FILL_436
timestamp 1680363874
transform 1 0 1432 0 -1 4370
box -8 -3 16 105
use FILL  FILL_437
timestamp 1680363874
transform 1 0 1440 0 -1 4370
box -8 -3 16 105
use FILL  FILL_438
timestamp 1680363874
transform 1 0 1448 0 -1 4370
box -8 -3 16 105
use FILL  FILL_439
timestamp 1680363874
transform 1 0 1456 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1680363874
transform 1 0 1464 0 -1 4370
box -8 -3 104 105
use FILL  FILL_440
timestamp 1680363874
transform 1 0 1560 0 -1 4370
box -8 -3 16 105
use FILL  FILL_441
timestamp 1680363874
transform 1 0 1568 0 -1 4370
box -8 -3 16 105
use FILL  FILL_445
timestamp 1680363874
transform 1 0 1576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_446
timestamp 1680363874
transform 1 0 1584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_447
timestamp 1680363874
transform 1 0 1592 0 -1 4370
box -8 -3 16 105
use FILL  FILL_448
timestamp 1680363874
transform 1 0 1600 0 -1 4370
box -8 -3 16 105
use FILL  FILL_449
timestamp 1680363874
transform 1 0 1608 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1680363874
transform -1 0 1632 0 -1 4370
box -9 -3 26 105
use FILL  FILL_450
timestamp 1680363874
transform 1 0 1632 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1680363874
transform 1 0 1640 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_50
timestamp 1680363874
transform -1 0 1752 0 -1 4370
box -9 -3 26 105
use FILL  FILL_451
timestamp 1680363874
transform 1 0 1752 0 -1 4370
box -8 -3 16 105
use FILL  FILL_452
timestamp 1680363874
transform 1 0 1760 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1680363874
transform 1 0 1768 0 -1 4370
box -9 -3 26 105
use OAI22X1  OAI22X1_46
timestamp 1680363874
transform -1 0 1824 0 -1 4370
box -8 -3 46 105
use FILL  FILL_475
timestamp 1680363874
transform 1 0 1824 0 -1 4370
box -8 -3 16 105
use FILL  FILL_476
timestamp 1680363874
transform 1 0 1832 0 -1 4370
box -8 -3 16 105
use FILL  FILL_477
timestamp 1680363874
transform 1 0 1840 0 -1 4370
box -8 -3 16 105
use FILL  FILL_478
timestamp 1680363874
transform 1 0 1848 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1680363874
transform -1 0 1952 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_55
timestamp 1680363874
transform -1 0 1968 0 -1 4370
box -9 -3 26 105
use FILL  FILL_479
timestamp 1680363874
transform 1 0 1968 0 -1 4370
box -8 -3 16 105
use FILL  FILL_480
timestamp 1680363874
transform 1 0 1976 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_22
timestamp 1680363874
transform -1 0 2024 0 -1 4370
box -8 -3 46 105
use INVX2  INVX2_56
timestamp 1680363874
transform 1 0 2024 0 -1 4370
box -9 -3 26 105
use FILL  FILL_481
timestamp 1680363874
transform 1 0 2040 0 -1 4370
box -8 -3 16 105
use FILL  FILL_482
timestamp 1680363874
transform 1 0 2048 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1680363874
transform -1 0 2152 0 -1 4370
box -8 -3 104 105
use FILL  FILL_483
timestamp 1680363874
transform 1 0 2152 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_47
timestamp 1680363874
transform 1 0 2160 0 -1 4370
box -8 -3 46 105
use FILL  FILL_484
timestamp 1680363874
transform 1 0 2200 0 -1 4370
box -8 -3 16 105
use FILL  FILL_485
timestamp 1680363874
transform 1 0 2208 0 -1 4370
box -8 -3 16 105
use FILL  FILL_486
timestamp 1680363874
transform 1 0 2216 0 -1 4370
box -8 -3 16 105
use FILL  FILL_487
timestamp 1680363874
transform 1 0 2224 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_23
timestamp 1680363874
transform -1 0 2272 0 -1 4370
box -8 -3 46 105
use FILL  FILL_488
timestamp 1680363874
transform 1 0 2272 0 -1 4370
box -8 -3 16 105
use FILL  FILL_489
timestamp 1680363874
transform 1 0 2280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_490
timestamp 1680363874
transform 1 0 2288 0 -1 4370
box -8 -3 16 105
use FILL  FILL_491
timestamp 1680363874
transform 1 0 2296 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1680363874
transform -1 0 2320 0 -1 4370
box -9 -3 26 105
use FILL  FILL_492
timestamp 1680363874
transform 1 0 2320 0 -1 4370
box -8 -3 16 105
use FILL  FILL_493
timestamp 1680363874
transform 1 0 2328 0 -1 4370
box -8 -3 16 105
use FILL  FILL_494
timestamp 1680363874
transform 1 0 2336 0 -1 4370
box -8 -3 16 105
use FILL  FILL_495
timestamp 1680363874
transform 1 0 2344 0 -1 4370
box -8 -3 16 105
use FILL  FILL_496
timestamp 1680363874
transform 1 0 2352 0 -1 4370
box -8 -3 16 105
use FILL  FILL_497
timestamp 1680363874
transform 1 0 2360 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_24
timestamp 1680363874
transform -1 0 2408 0 -1 4370
box -8 -3 46 105
use FILL  FILL_498
timestamp 1680363874
transform 1 0 2408 0 -1 4370
box -8 -3 16 105
use FILL  FILL_499
timestamp 1680363874
transform 1 0 2416 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1680363874
transform 1 0 2424 0 -1 4370
box -8 -3 104 105
use FILL  FILL_500
timestamp 1680363874
transform 1 0 2520 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_781
timestamp 1680363874
transform 1 0 2564 0 1 4275
box -3 -3 3 3
use AOI22X1  AOI22X1_25
timestamp 1680363874
transform -1 0 2568 0 -1 4370
box -8 -3 46 105
use FILL  FILL_501
timestamp 1680363874
transform 1 0 2568 0 -1 4370
box -8 -3 16 105
use FILL  FILL_503
timestamp 1680363874
transform 1 0 2576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1680363874
transform 1 0 2584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_505
timestamp 1680363874
transform 1 0 2592 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_58
timestamp 1680363874
transform 1 0 2600 0 -1 4370
box -9 -3 26 105
use FILL  FILL_506
timestamp 1680363874
transform 1 0 2616 0 -1 4370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1680363874
transform 1 0 2624 0 -1 4370
box -8 -3 16 105
use FILL  FILL_508
timestamp 1680363874
transform 1 0 2632 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_27
timestamp 1680363874
transform 1 0 2640 0 -1 4370
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1680363874
transform 1 0 2680 0 -1 4370
box -8 -3 46 105
use FILL  FILL_528
timestamp 1680363874
transform 1 0 2720 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_49
timestamp 1680363874
transform -1 0 2768 0 -1 4370
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1680363874
transform -1 0 2808 0 -1 4370
box -8 -3 46 105
use FILL  FILL_529
timestamp 1680363874
transform 1 0 2808 0 -1 4370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1680363874
transform 1 0 2816 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_782
timestamp 1680363874
transform 1 0 2844 0 1 4275
box -3 -3 3 3
use OAI22X1  OAI22X1_51
timestamp 1680363874
transform -1 0 2864 0 -1 4370
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1680363874
transform -1 0 2904 0 -1 4370
box -8 -3 46 105
use FILL  FILL_531
timestamp 1680363874
transform 1 0 2904 0 -1 4370
box -8 -3 16 105
use FILL  FILL_532
timestamp 1680363874
transform 1 0 2912 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1680363874
transform 1 0 2920 0 -1 4370
box -9 -3 26 105
use FILL  FILL_533
timestamp 1680363874
transform 1 0 2936 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_783
timestamp 1680363874
transform 1 0 2988 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1680363874
transform -1 0 3040 0 -1 4370
box -8 -3 104 105
use FILL  FILL_534
timestamp 1680363874
transform 1 0 3040 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_784
timestamp 1680363874
transform 1 0 3060 0 1 4275
box -3 -3 3 3
use FILL  FILL_535
timestamp 1680363874
transform 1 0 3048 0 -1 4370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1680363874
transform 1 0 3056 0 -1 4370
box -8 -3 16 105
use FILL  FILL_537
timestamp 1680363874
transform 1 0 3064 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_785
timestamp 1680363874
transform 1 0 3100 0 1 4275
box -3 -3 3 3
use AOI22X1  AOI22X1_32
timestamp 1680363874
transform 1 0 3072 0 -1 4370
box -8 -3 46 105
use FILL  FILL_538
timestamp 1680363874
transform 1 0 3112 0 -1 4370
box -8 -3 16 105
use FILL  FILL_539
timestamp 1680363874
transform 1 0 3120 0 -1 4370
box -8 -3 16 105
use FILL  FILL_540
timestamp 1680363874
transform 1 0 3128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_541
timestamp 1680363874
transform 1 0 3136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_542
timestamp 1680363874
transform 1 0 3144 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_52
timestamp 1680363874
transform -1 0 3192 0 -1 4370
box -8 -3 46 105
use FILL  FILL_543
timestamp 1680363874
transform 1 0 3192 0 -1 4370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1680363874
transform 1 0 3200 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_786
timestamp 1680363874
transform 1 0 3300 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_70
timestamp 1680363874
transform -1 0 3304 0 -1 4370
box -8 -3 104 105
use FILL  FILL_545
timestamp 1680363874
transform 1 0 3304 0 -1 4370
box -8 -3 16 105
use FILL  FILL_547
timestamp 1680363874
transform 1 0 3312 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_787
timestamp 1680363874
transform 1 0 3332 0 1 4275
box -3 -3 3 3
use OAI22X1  OAI22X1_53
timestamp 1680363874
transform 1 0 3320 0 -1 4370
box -8 -3 46 105
use FILL  FILL_553
timestamp 1680363874
transform 1 0 3360 0 -1 4370
box -8 -3 16 105
use FILL  FILL_554
timestamp 1680363874
transform 1 0 3368 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_788
timestamp 1680363874
transform 1 0 3388 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_72
timestamp 1680363874
transform -1 0 3472 0 -1 4370
box -8 -3 104 105
use FILL  FILL_555
timestamp 1680363874
transform 1 0 3472 0 -1 4370
box -8 -3 16 105
use FILL  FILL_556
timestamp 1680363874
transform 1 0 3480 0 -1 4370
box -8 -3 16 105
use FILL  FILL_557
timestamp 1680363874
transform 1 0 3488 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_36
timestamp 1680363874
transform 1 0 3496 0 -1 4370
box -8 -3 46 105
use INVX2  INVX2_64
timestamp 1680363874
transform 1 0 3536 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1680363874
transform -1 0 3648 0 -1 4370
box -8 -3 104 105
use FILL  FILL_573
timestamp 1680363874
transform 1 0 3648 0 -1 4370
box -8 -3 16 105
use FILL  FILL_574
timestamp 1680363874
transform 1 0 3656 0 -1 4370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1680363874
transform 1 0 3664 0 -1 4370
box -8 -3 16 105
use FILL  FILL_576
timestamp 1680363874
transform 1 0 3672 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1680363874
transform 1 0 3680 0 -1 4370
box -8 -3 46 105
use FILL  FILL_577
timestamp 1680363874
transform 1 0 3720 0 -1 4370
box -8 -3 16 105
use FILL  FILL_578
timestamp 1680363874
transform 1 0 3728 0 -1 4370
box -8 -3 16 105
use FILL  FILL_579
timestamp 1680363874
transform 1 0 3736 0 -1 4370
box -8 -3 16 105
use FILL  FILL_580
timestamp 1680363874
transform 1 0 3744 0 -1 4370
box -8 -3 16 105
use FILL  FILL_581
timestamp 1680363874
transform 1 0 3752 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_54
timestamp 1680363874
transform 1 0 3760 0 -1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1680363874
transform -1 0 3896 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_65
timestamp 1680363874
transform 1 0 3896 0 -1 4370
box -9 -3 26 105
use FILL  FILL_582
timestamp 1680363874
transform 1 0 3912 0 -1 4370
box -8 -3 16 105
use FILL  FILL_585
timestamp 1680363874
transform 1 0 3920 0 -1 4370
box -8 -3 16 105
use FILL  FILL_586
timestamp 1680363874
transform 1 0 3928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_587
timestamp 1680363874
transform 1 0 3936 0 -1 4370
box -8 -3 16 105
use FILL  FILL_588
timestamp 1680363874
transform 1 0 3944 0 -1 4370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1680363874
transform 1 0 3952 0 -1 4370
box -8 -3 16 105
use FILL  FILL_590
timestamp 1680363874
transform 1 0 3960 0 -1 4370
box -8 -3 16 105
use FILL  FILL_591
timestamp 1680363874
transform 1 0 3968 0 -1 4370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1680363874
transform 1 0 3976 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_66
timestamp 1680363874
transform 1 0 3984 0 -1 4370
box -9 -3 26 105
use FILL  FILL_597
timestamp 1680363874
transform 1 0 4000 0 -1 4370
box -8 -3 16 105
use FILL  FILL_608
timestamp 1680363874
transform 1 0 4008 0 -1 4370
box -8 -3 16 105
use FILL  FILL_609
timestamp 1680363874
transform 1 0 4016 0 -1 4370
box -8 -3 16 105
use FILL  FILL_610
timestamp 1680363874
transform 1 0 4024 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_55
timestamp 1680363874
transform 1 0 4032 0 -1 4370
box -8 -3 46 105
use FILL  FILL_611
timestamp 1680363874
transform 1 0 4072 0 -1 4370
box -8 -3 16 105
use FILL  FILL_612
timestamp 1680363874
transform 1 0 4080 0 -1 4370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1680363874
transform 1 0 4088 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_40
timestamp 1680363874
transform 1 0 4096 0 -1 4370
box -8 -3 46 105
use FILL  FILL_614
timestamp 1680363874
transform 1 0 4136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_617
timestamp 1680363874
transform 1 0 4144 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_56
timestamp 1680363874
transform 1 0 4152 0 -1 4370
box -8 -3 46 105
use FILL  FILL_618
timestamp 1680363874
transform 1 0 4192 0 -1 4370
box -8 -3 16 105
use FILL  FILL_619
timestamp 1680363874
transform 1 0 4200 0 -1 4370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1680363874
transform 1 0 4208 0 -1 4370
box -8 -3 16 105
use FILL  FILL_621
timestamp 1680363874
transform 1 0 4216 0 -1 4370
box -8 -3 16 105
use FILL  FILL_622
timestamp 1680363874
transform 1 0 4224 0 -1 4370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1680363874
transform 1 0 4232 0 -1 4370
box -8 -3 16 105
use FILL  FILL_624
timestamp 1680363874
transform 1 0 4240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_625
timestamp 1680363874
transform 1 0 4248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_626
timestamp 1680363874
transform 1 0 4256 0 -1 4370
box -8 -3 16 105
use FILL  FILL_627
timestamp 1680363874
transform 1 0 4264 0 -1 4370
box -8 -3 16 105
use FILL  FILL_628
timestamp 1680363874
transform 1 0 4272 0 -1 4370
box -8 -3 16 105
use FILL  FILL_629
timestamp 1680363874
transform 1 0 4280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_630
timestamp 1680363874
transform 1 0 4288 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_57
timestamp 1680363874
transform 1 0 4296 0 -1 4370
box -8 -3 46 105
use FILL  FILL_637
timestamp 1680363874
transform 1 0 4336 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_58
timestamp 1680363874
transform 1 0 4344 0 -1 4370
box -8 -3 46 105
use FILL  FILL_642
timestamp 1680363874
transform 1 0 4384 0 -1 4370
box -8 -3 16 105
use FILL  FILL_644
timestamp 1680363874
transform 1 0 4392 0 -1 4370
box -8 -3 16 105
use FILL  FILL_652
timestamp 1680363874
transform 1 0 4400 0 -1 4370
box -8 -3 16 105
use FILL  FILL_653
timestamp 1680363874
transform 1 0 4408 0 -1 4370
box -8 -3 16 105
use FILL  FILL_654
timestamp 1680363874
transform 1 0 4416 0 -1 4370
box -8 -3 16 105
use FILL  FILL_655
timestamp 1680363874
transform 1 0 4424 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1680363874
transform 1 0 4432 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1680363874
transform 1 0 4448 0 -1 4370
box -8 -3 104 105
use FILL  FILL_656
timestamp 1680363874
transform 1 0 4544 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_72
timestamp 1680363874
transform 1 0 4552 0 -1 4370
box -9 -3 26 105
use FILL  FILL_669
timestamp 1680363874
transform 1 0 4568 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1680363874
transform 1 0 4576 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1680363874
transform -1 0 4688 0 -1 4370
box -8 -3 104 105
use FILL  FILL_670
timestamp 1680363874
transform 1 0 4688 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1680363874
transform -1 0 4792 0 -1 4370
box -8 -3 104 105
use FILL  FILL_671
timestamp 1680363874
transform 1 0 4792 0 -1 4370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_9
timestamp 1680363874
transform 1 0 4851 0 1 4270
box -10 -3 10 3
use M3_M2  M3_M2_907
timestamp 1680363874
transform 1 0 68 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1076
timestamp 1680363874
transform 1 0 68 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_821
timestamp 1680363874
transform 1 0 188 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1680363874
transform 1 0 172 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_952
timestamp 1680363874
transform 1 0 172 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1680363874
transform 1 0 188 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1680363874
transform 1 0 164 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1680363874
transform 1 0 180 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_954
timestamp 1680363874
transform 1 0 164 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1680363874
transform 1 0 188 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1680363874
transform 1 0 204 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_956
timestamp 1680363874
transform 1 0 204 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1680363874
transform 1 0 236 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1680363874
transform 1 0 268 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_954
timestamp 1680363874
transform 1 0 284 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1680363874
transform 1 0 236 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_957
timestamp 1680363874
transform 1 0 236 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1680363874
transform 1 0 284 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1680363874
transform 1 0 332 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1680363874
transform 1 0 372 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1680363874
transform 1 0 380 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_955
timestamp 1680363874
transform 1 0 364 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1680363874
transform 1 0 380 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1680363874
transform 1 0 356 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_939
timestamp 1680363874
transform 1 0 364 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1082
timestamp 1680363874
transform 1 0 372 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_959
timestamp 1680363874
transform 1 0 372 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1680363874
transform 1 0 380 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1680363874
transform 1 0 428 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_910
timestamp 1680363874
transform 1 0 460 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_957
timestamp 1680363874
transform 1 0 484 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1680363874
transform 1 0 460 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_989
timestamp 1680363874
transform 1 0 460 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_958
timestamp 1680363874
transform 1 0 556 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_823
timestamp 1680363874
transform 1 0 604 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1680363874
transform 1 0 612 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1680363874
transform 1 0 588 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_911
timestamp 1680363874
transform 1 0 596 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_960
timestamp 1680363874
transform 1 0 604 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1680363874
transform 1 0 580 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1680363874
transform 1 0 596 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1680363874
transform 1 0 612 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1680363874
transform 1 0 620 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1680363874
transform 1 0 580 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1680363874
transform 1 0 636 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1680363874
transform 1 0 628 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_961
timestamp 1680363874
transform 1 0 628 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_961
timestamp 1680363874
transform 1 0 620 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1680363874
transform 1 0 636 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1680363874
transform 1 0 676 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1680363874
transform 1 0 676 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_962
timestamp 1680363874
transform 1 0 668 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1680363874
transform 1 0 660 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_941
timestamp 1680363874
transform 1 0 668 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1090
timestamp 1680363874
transform 1 0 676 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_962
timestamp 1680363874
transform 1 0 660 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_963
timestamp 1680363874
transform 1 0 700 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_942
timestamp 1680363874
transform 1 0 692 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1680363874
transform 1 0 740 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1680363874
transform 1 0 732 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_964
timestamp 1680363874
transform 1 0 740 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1680363874
transform 1 0 716 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1680363874
transform 1 0 732 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1680363874
transform 1 0 748 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1680363874
transform 1 0 756 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_799
timestamp 1680363874
transform 1 0 764 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1680363874
transform 1 0 756 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1680363874
transform 1 0 788 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1680363874
transform 1 0 788 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1680363874
transform 1 0 804 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_949
timestamp 1680363874
transform 1 0 796 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1680363874
transform 1 0 780 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_912
timestamp 1680363874
transform 1 0 804 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1680363874
transform 1 0 796 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_990
timestamp 1680363874
transform 1 0 780 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1096
timestamp 1680363874
transform 1 0 804 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1680363874
transform 1 0 820 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_943
timestamp 1680363874
transform 1 0 820 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1680363874
transform 1 0 860 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1680363874
transform 1 0 868 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_913
timestamp 1680363874
transform 1 0 868 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1097
timestamp 1680363874
transform 1 0 852 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1680363874
transform 1 0 860 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1680363874
transform 1 0 892 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_967
timestamp 1680363874
transform 1 0 892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1680363874
transform 1 0 924 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1680363874
transform 1 0 924 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1680363874
transform 1 0 924 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_826
timestamp 1680363874
transform 1 0 964 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1680363874
transform 1 0 980 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1680363874
transform 1 0 996 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_968
timestamp 1680363874
transform 1 0 964 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1680363874
transform 1 0 988 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1680363874
transform 1 0 964 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_944
timestamp 1680363874
transform 1 0 972 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1101
timestamp 1680363874
transform 1 0 980 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1680363874
transform 1 0 996 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_827
timestamp 1680363874
transform 1 0 1020 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_970
timestamp 1680363874
transform 1 0 1012 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_875
timestamp 1680363874
transform 1 0 1036 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1680363874
transform 1 0 1028 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1680363874
transform 1 0 1076 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1680363874
transform 1 0 1092 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1680363874
transform 1 0 1052 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1680363874
transform 1 0 1068 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1680363874
transform 1 0 1076 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1680363874
transform 1 0 1092 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1680363874
transform 1 0 1028 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1680363874
transform 1 0 1044 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1680363874
transform 1 0 1060 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1680363874
transform 1 0 1068 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1680363874
transform 1 0 1084 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1680363874
transform 1 0 1100 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1680363874
transform 1 0 1084 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1680363874
transform 1 0 1044 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1680363874
transform 1 0 1060 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1680363874
transform 1 0 1100 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1680363874
transform 1 0 1116 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_974
timestamp 1680363874
transform 1 0 1124 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1680363874
transform 1 0 1180 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1680363874
transform 1 0 1204 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_965
timestamp 1680363874
transform 1 0 1180 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1680363874
transform 1 0 1228 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1110
timestamp 1680363874
transform 1 0 1228 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1680363874
transform 1 0 1244 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1680363874
transform 1 0 1260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1680363874
transform 1 0 1276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1680363874
transform 1 0 1252 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1680363874
transform 1 0 1268 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_966
timestamp 1680363874
transform 1 0 1252 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1680363874
transform 1 0 1276 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1680363874
transform 1 0 1300 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1113
timestamp 1680363874
transform 1 0 1292 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1680363874
transform 1 0 1300 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_967
timestamp 1680363874
transform 1 0 1292 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_979
timestamp 1680363874
transform 1 0 1340 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_877
timestamp 1680363874
transform 1 0 1364 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_980
timestamp 1680363874
transform 1 0 1356 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1680363874
transform 1 0 1316 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1680363874
transform 1 0 1332 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1680363874
transform 1 0 1348 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_946
timestamp 1680363874
transform 1 0 1356 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1680363874
transform 1 0 1348 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1680363874
transform 1 0 1388 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1680363874
transform 1 0 1380 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_994
timestamp 1680363874
transform 1 0 1388 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1680363874
transform 1 0 1404 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1680363874
transform 1 0 1468 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1680363874
transform 1 0 1468 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1680363874
transform 1 0 1516 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_879
timestamp 1680363874
transform 1 0 1652 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1680363874
transform 1 0 1692 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_983
timestamp 1680363874
transform 1 0 1652 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1680363874
transform 1 0 1684 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1680363874
transform 1 0 1692 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1680363874
transform 1 0 1604 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_970
timestamp 1680363874
transform 1 0 1604 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1680363874
transform 1 0 1644 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1680363874
transform 1 0 1708 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1680363874
transform 1 0 1716 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_986
timestamp 1680363874
transform 1 0 1724 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1680363874
transform 1 0 1708 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1680363874
transform 1 0 1716 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_972
timestamp 1680363874
transform 1 0 1700 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1680363874
transform 1 0 1684 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1680363874
transform 1 0 1716 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1123
timestamp 1680363874
transform 1 0 1732 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_829
timestamp 1680363874
transform 1 0 1748 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1680363874
transform 1 0 1796 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1680363874
transform 1 0 1788 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_987
timestamp 1680363874
transform 1 0 1748 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1680363874
transform 1 0 1764 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_921
timestamp 1680363874
transform 1 0 1772 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1680363874
transform 1 0 1764 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1680363874
transform 1 0 1812 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_989
timestamp 1680363874
transform 1 0 1788 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1680363874
transform 1 0 1796 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1680363874
transform 1 0 1812 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1680363874
transform 1 0 1772 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1680363874
transform 1 0 1780 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_996
timestamp 1680363874
transform 1 0 1780 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1680363874
transform 1 0 1820 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1680363874
transform 1 0 1796 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1126
timestamp 1680363874
transform 1 0 1820 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_831
timestamp 1680363874
transform 1 0 1836 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1680363874
transform 1 0 1836 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1680363874
transform 1 0 1852 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_789
timestamp 1680363874
transform 1 0 1868 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1680363874
transform 1 0 1876 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1680363874
transform 1 0 1868 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1680363874
transform 1 0 1884 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1680363874
transform 1 0 1892 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1680363874
transform 1 0 1868 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1128
timestamp 1680363874
transform 1 0 1892 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_974
timestamp 1680363874
transform 1 0 1884 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1680363874
transform 1 0 1916 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1680363874
transform 1 0 1940 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1680363874
transform 1 0 1932 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1680363874
transform 1 0 1924 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1680363874
transform 1 0 1924 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1680363874
transform 1 0 1932 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1680363874
transform 1 0 1948 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_924
timestamp 1680363874
transform 1 0 1956 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1680363874
transform 1 0 1972 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1680363874
transform 1 0 1940 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1680363874
transform 1 0 1956 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1680363874
transform 1 0 1964 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_975
timestamp 1680363874
transform 1 0 1940 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1680363874
transform 1 0 1932 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_999
timestamp 1680363874
transform 1 0 1996 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_802
timestamp 1680363874
transform 1 0 2012 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1680363874
transform 1 0 2020 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1680363874
transform 1 0 2012 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_998
timestamp 1680363874
transform 1 0 2012 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1680363874
transform 1 0 2036 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1680363874
transform 1 0 2028 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1680363874
transform 1 0 2076 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1680363874
transform 1 0 2084 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1680363874
transform 1 0 2068 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1680363874
transform 1 0 2084 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1680363874
transform 1 0 2060 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1680363874
transform 1 0 2076 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1680363874
transform 1 0 2084 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1680363874
transform 1 0 2116 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_950
timestamp 1680363874
transform 1 0 2148 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1680363874
transform 1 0 2164 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1680363874
transform 1 0 2188 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1680363874
transform 1 0 2196 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1680363874
transform 1 0 2180 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1680363874
transform 1 0 2172 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1680363874
transform 1 0 2204 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1680363874
transform 1 0 2164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1680363874
transform 1 0 2180 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1680363874
transform 1 0 2196 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1680363874
transform 1 0 2204 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1680363874
transform 1 0 2172 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_951
timestamp 1680363874
transform 1 0 2180 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1137
timestamp 1680363874
transform 1 0 2212 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_976
timestamp 1680363874
transform 1 0 2212 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1680363874
transform 1 0 2260 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1680363874
transform 1 0 2236 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_1138
timestamp 1680363874
transform 1 0 2228 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1680363874
transform 1 0 2244 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1680363874
transform 1 0 2260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1680363874
transform 1 0 2252 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1680363874
transform 1 0 2268 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_887
timestamp 1680363874
transform 1 0 2348 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1680363874
transform 1 0 2348 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1680363874
transform 1 0 2380 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1680363874
transform 1 0 2300 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1680363874
transform 1 0 2340 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1680363874
transform 1 0 2396 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1680363874
transform 1 0 2404 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1012
timestamp 1680363874
transform 1 0 2404 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1680363874
transform 1 0 2404 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_1000
timestamp 1680363874
transform 1 0 2436 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1013
timestamp 1680363874
transform 1 0 2460 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_925
timestamp 1680363874
transform 1 0 2468 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1680363874
transform 1 0 2500 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1680363874
transform 1 0 2524 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1143
timestamp 1680363874
transform 1 0 2524 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1680363874
transform 1 0 2612 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1680363874
transform 1 0 2572 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1680363874
transform 1 0 2620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1680363874
transform 1 0 2540 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1680363874
transform 1 0 2636 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_849
timestamp 1680363874
transform 1 0 2652 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1680363874
transform 1 0 2676 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1680363874
transform 1 0 2692 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1680363874
transform 1 0 2676 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1680363874
transform 1 0 2660 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1680363874
transform 1 0 2676 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1680363874
transform 1 0 2652 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1680363874
transform 1 0 2700 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1018
timestamp 1680363874
transform 1 0 2692 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_977
timestamp 1680363874
transform 1 0 2676 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1019
timestamp 1680363874
transform 1 0 2716 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1680363874
transform 1 0 2748 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1680363874
transform 1 0 2756 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1020
timestamp 1680363874
transform 1 0 2748 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1680363874
transform 1 0 2732 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1680363874
transform 1 0 2740 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1680363874
transform 1 0 2756 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1680363874
transform 1 0 2764 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_978
timestamp 1680363874
transform 1 0 2764 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1680363874
transform 1 0 2812 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1680363874
transform 1 0 2812 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_852
timestamp 1680363874
transform 1 0 2828 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1022
timestamp 1680363874
transform 1 0 2828 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1680363874
transform 1 0 2844 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1680363874
transform 1 0 2852 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1680363874
transform 1 0 2916 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1680363874
transform 1 0 2892 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1680363874
transform 1 0 2908 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1680363874
transform 1 0 2956 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1680363874
transform 1 0 2852 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1680363874
transform 1 0 2868 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1680363874
transform 1 0 2876 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1680363874
transform 1 0 2908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1680363874
transform 1 0 2836 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1680363874
transform 1 0 2844 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1680363874
transform 1 0 2868 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1680363874
transform 1 0 2956 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1680363874
transform 1 0 2836 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1680363874
transform 1 0 2972 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1680363874
transform 1 0 3028 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1680363874
transform 1 0 3052 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1680363874
transform 1 0 3076 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1680363874
transform 1 0 3068 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1680363874
transform 1 0 3052 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_980
timestamp 1680363874
transform 1 0 3044 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1680363874
transform 1 0 3060 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1028
timestamp 1680363874
transform 1 0 3076 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_896
timestamp 1680363874
transform 1 0 3092 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1680363874
transform 1 0 3180 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1680363874
transform 1 0 3132 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1680363874
transform 1 0 3172 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1680363874
transform 1 0 3156 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1029
timestamp 1680363874
transform 1 0 3156 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1680363874
transform 1 0 3180 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1680363874
transform 1 0 3196 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1030
timestamp 1680363874
transform 1 0 3196 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_927
timestamp 1680363874
transform 1 0 3212 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1680363874
transform 1 0 3244 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1680363874
transform 1 0 3252 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1031
timestamp 1680363874
transform 1 0 3244 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1680363874
transform 1 0 3260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1680363874
transform 1 0 3276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1680363874
transform 1 0 3244 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1680363874
transform 1 0 3252 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1680363874
transform 1 0 3268 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_981
timestamp 1680363874
transform 1 0 3276 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1680363874
transform 1 0 3292 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1680363874
transform 1 0 3332 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1034
timestamp 1680363874
transform 1 0 3300 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1680363874
transform 1 0 3316 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1680363874
transform 1 0 3332 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1680363874
transform 1 0 3308 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1680363874
transform 1 0 3324 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1680363874
transform 1 0 3332 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_982
timestamp 1680363874
transform 1 0 3300 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1680363874
transform 1 0 3356 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1037
timestamp 1680363874
transform 1 0 3412 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_814
timestamp 1680363874
transform 1 0 3532 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1680363874
transform 1 0 3524 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1680363874
transform 1 0 3564 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1038
timestamp 1680363874
transform 1 0 3524 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1680363874
transform 1 0 3556 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1680363874
transform 1 0 3564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1680363874
transform 1 0 3476 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1680363874
transform 1 0 3588 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1680363874
transform 1 0 3636 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1041
timestamp 1680363874
transform 1 0 3620 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_929
timestamp 1680363874
transform 1 0 3628 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1042
timestamp 1680363874
transform 1 0 3636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1680363874
transform 1 0 3612 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1680363874
transform 1 0 3628 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1680363874
transform 1 0 3652 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_815
timestamp 1680363874
transform 1 0 3716 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1680363874
transform 1 0 3724 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1680363874
transform 1 0 3764 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1680363874
transform 1 0 3676 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1680363874
transform 1 0 3724 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1680363874
transform 1 0 3748 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1044
timestamp 1680363874
transform 1 0 3756 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1680363874
transform 1 0 3764 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1680363874
transform 1 0 3676 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_983
timestamp 1680363874
transform 1 0 3772 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1680363874
transform 1 0 3804 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1046
timestamp 1680363874
transform 1 0 3804 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_837
timestamp 1680363874
transform 1 0 3844 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1680363874
transform 1 0 3820 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1047
timestamp 1680363874
transform 1 0 3828 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1680363874
transform 1 0 3844 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1680363874
transform 1 0 3812 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1680363874
transform 1 0 3820 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1680363874
transform 1 0 3836 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_796
timestamp 1680363874
transform 1 0 3908 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1680363874
transform 1 0 3884 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1680363874
transform 1 0 3876 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1680363874
transform 1 0 3892 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1049
timestamp 1680363874
transform 1 0 3884 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1680363874
transform 1 0 3892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1680363874
transform 1 0 3908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1680363874
transform 1 0 3876 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1680363874
transform 1 0 3900 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_1002
timestamp 1680363874
transform 1 0 3892 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1052
timestamp 1680363874
transform 1 0 3940 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1680363874
transform 1 0 3964 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1053
timestamp 1680363874
transform 1 0 3996 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1680363874
transform 1 0 4028 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1680363874
transform 1 0 4076 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_862
timestamp 1680363874
transform 1 0 4092 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1680363874
transform 1 0 4108 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1055
timestamp 1680363874
transform 1 0 4116 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_817
timestamp 1680363874
transform 1 0 4164 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1056
timestamp 1680363874
transform 1 0 4164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1680363874
transform 1 0 4164 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_818
timestamp 1680363874
transform 1 0 4188 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1680363874
transform 1 0 4196 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1680363874
transform 1 0 4292 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1680363874
transform 1 0 4324 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1680363874
transform 1 0 4276 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1680363874
transform 1 0 4316 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1057
timestamp 1680363874
transform 1 0 4196 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1680363874
transform 1 0 4212 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1680363874
transform 1 0 4276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1680363874
transform 1 0 4188 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1680363874
transform 1 0 4204 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_984
timestamp 1680363874
transform 1 0 4204 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1680363874
transform 1 0 4300 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1060
timestamp 1680363874
transform 1 0 4308 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1680363874
transform 1 0 4316 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1680363874
transform 1 0 4228 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_1003
timestamp 1680363874
transform 1 0 4212 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1680363874
transform 1 0 4244 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1680363874
transform 1 0 4332 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1680363874
transform 1 0 4348 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1680363874
transform 1 0 4340 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1680363874
transform 1 0 4364 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1062
timestamp 1680363874
transform 1 0 4348 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1680363874
transform 1 0 4356 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1680363874
transform 1 0 4364 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1680363874
transform 1 0 4380 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1680363874
transform 1 0 4388 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1680363874
transform 1 0 4348 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1680363874
transform 1 0 4356 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1680363874
transform 1 0 4372 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_985
timestamp 1680363874
transform 1 0 4372 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1680363874
transform 1 0 4420 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1680363874
transform 1 0 4452 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1066
timestamp 1680363874
transform 1 0 4420 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1680363874
transform 1 0 4436 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1680363874
transform 1 0 4452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1680363874
transform 1 0 4428 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_936
timestamp 1680363874
transform 1 0 4492 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1069
timestamp 1680363874
transform 1 0 4500 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1680363874
transform 1 0 4516 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1680363874
transform 1 0 4492 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1680363874
transform 1 0 4508 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_905
timestamp 1680363874
transform 1 0 4548 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1680363874
transform 1 0 4540 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1071
timestamp 1680363874
transform 1 0 4548 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1680363874
transform 1 0 4548 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_986
timestamp 1680363874
transform 1 0 4548 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1072
timestamp 1680363874
transform 1 0 4572 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1680363874
transform 1 0 4588 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1680363874
transform 1 0 4564 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1680363874
transform 1 0 4580 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_987
timestamp 1680363874
transform 1 0 4580 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1680363874
transform 1 0 4564 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1680363874
transform 1 0 4620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1680363874
transform 1 0 4596 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1680363874
transform 1 0 4604 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1680363874
transform 1 0 4628 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1680363874
transform 1 0 4636 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_1006
timestamp 1680363874
transform 1 0 4612 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1680363874
transform 1 0 4628 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1680363874
transform 1 0 4692 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1680363874
transform 1 0 4748 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1075
timestamp 1680363874
transform 1 0 4756 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1680363874
transform 1 0 4780 0 1 4205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_10
timestamp 1680363874
transform 1 0 48 0 1 4170
box -10 -3 10 3
use FILL  FILL_672
timestamp 1680363874
transform 1 0 72 0 1 4170
box -8 -3 16 105
use FILL  FILL_673
timestamp 1680363874
transform 1 0 80 0 1 4170
box -8 -3 16 105
use FILL  FILL_674
timestamp 1680363874
transform 1 0 88 0 1 4170
box -8 -3 16 105
use FILL  FILL_675
timestamp 1680363874
transform 1 0 96 0 1 4170
box -8 -3 16 105
use FILL  FILL_676
timestamp 1680363874
transform 1 0 104 0 1 4170
box -8 -3 16 105
use FILL  FILL_677
timestamp 1680363874
transform 1 0 112 0 1 4170
box -8 -3 16 105
use FILL  FILL_678
timestamp 1680363874
transform 1 0 120 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1680363874
transform 1 0 128 0 1 4170
box -9 -3 26 105
use FILL  FILL_679
timestamp 1680363874
transform 1 0 144 0 1 4170
box -8 -3 16 105
use FILL  FILL_680
timestamp 1680363874
transform 1 0 152 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_59
timestamp 1680363874
transform 1 0 160 0 1 4170
box -8 -3 46 105
use FILL  FILL_681
timestamp 1680363874
transform 1 0 200 0 1 4170
box -8 -3 16 105
use FILL  FILL_682
timestamp 1680363874
transform 1 0 208 0 1 4170
box -8 -3 16 105
use FILL  FILL_683
timestamp 1680363874
transform 1 0 216 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1680363874
transform 1 0 224 0 1 4170
box -8 -3 104 105
use FILL  FILL_684
timestamp 1680363874
transform 1 0 320 0 1 4170
box -8 -3 16 105
use FILL  FILL_685
timestamp 1680363874
transform 1 0 328 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_75
timestamp 1680363874
transform 1 0 336 0 1 4170
box -9 -3 26 105
use OAI22X1  OAI22X1_60
timestamp 1680363874
transform 1 0 352 0 1 4170
box -8 -3 46 105
use FILL  FILL_686
timestamp 1680363874
transform 1 0 392 0 1 4170
box -8 -3 16 105
use FILL  FILL_687
timestamp 1680363874
transform 1 0 400 0 1 4170
box -8 -3 16 105
use FILL  FILL_688
timestamp 1680363874
transform 1 0 408 0 1 4170
box -8 -3 16 105
use FILL  FILL_689
timestamp 1680363874
transform 1 0 416 0 1 4170
box -8 -3 16 105
use FILL  FILL_690
timestamp 1680363874
transform 1 0 424 0 1 4170
box -8 -3 16 105
use FILL  FILL_691
timestamp 1680363874
transform 1 0 432 0 1 4170
box -8 -3 16 105
use FILL  FILL_698
timestamp 1680363874
transform 1 0 440 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1680363874
transform 1 0 448 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_79
timestamp 1680363874
transform 1 0 544 0 1 4170
box -9 -3 26 105
use FILL  FILL_700
timestamp 1680363874
transform 1 0 560 0 1 4170
box -8 -3 16 105
use FILL  FILL_701
timestamp 1680363874
transform 1 0 568 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_63
timestamp 1680363874
transform 1 0 576 0 1 4170
box -8 -3 46 105
use FILL  FILL_702
timestamp 1680363874
transform 1 0 616 0 1 4170
box -8 -3 16 105
use FILL  FILL_703
timestamp 1680363874
transform 1 0 624 0 1 4170
box -8 -3 16 105
use FILL  FILL_704
timestamp 1680363874
transform 1 0 632 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_64
timestamp 1680363874
transform 1 0 640 0 1 4170
box -8 -3 46 105
use FILL  FILL_705
timestamp 1680363874
transform 1 0 680 0 1 4170
box -8 -3 16 105
use FILL  FILL_721
timestamp 1680363874
transform 1 0 688 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1008
timestamp 1680363874
transform 1 0 708 0 1 4175
box -3 -3 3 3
use FILL  FILL_722
timestamp 1680363874
transform 1 0 696 0 1 4170
box -8 -3 16 105
use FILL  FILL_723
timestamp 1680363874
transform 1 0 704 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_68
timestamp 1680363874
transform 1 0 712 0 1 4170
box -8 -3 46 105
use FILL  FILL_724
timestamp 1680363874
transform 1 0 752 0 1 4170
box -8 -3 16 105
use FILL  FILL_729
timestamp 1680363874
transform 1 0 760 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_10
timestamp 1680363874
transform 1 0 768 0 1 4170
box -8 -3 34 105
use FILL  FILL_730
timestamp 1680363874
transform 1 0 800 0 1 4170
box -8 -3 16 105
use FILL  FILL_733
timestamp 1680363874
transform 1 0 808 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_12
timestamp 1680363874
transform 1 0 816 0 1 4170
box -8 -3 34 105
use M3_M2  M3_M2_1009
timestamp 1680363874
transform 1 0 860 0 1 4175
box -3 -3 3 3
use FILL  FILL_735
timestamp 1680363874
transform 1 0 848 0 1 4170
box -8 -3 16 105
use FILL  FILL_736
timestamp 1680363874
transform 1 0 856 0 1 4170
box -8 -3 16 105
use FILL  FILL_741
timestamp 1680363874
transform 1 0 864 0 1 4170
box -8 -3 16 105
use FILL  FILL_743
timestamp 1680363874
transform 1 0 872 0 1 4170
box -8 -3 16 105
use FILL  FILL_745
timestamp 1680363874
transform 1 0 880 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_13
timestamp 1680363874
transform 1 0 888 0 1 4170
box -8 -3 34 105
use FILL  FILL_747
timestamp 1680363874
transform 1 0 920 0 1 4170
box -8 -3 16 105
use FILL  FILL_749
timestamp 1680363874
transform 1 0 928 0 1 4170
box -8 -3 16 105
use FILL  FILL_751
timestamp 1680363874
transform 1 0 936 0 1 4170
box -8 -3 16 105
use FILL  FILL_753
timestamp 1680363874
transform 1 0 944 0 1 4170
box -8 -3 16 105
use FILL  FILL_755
timestamp 1680363874
transform 1 0 952 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_70
timestamp 1680363874
transform 1 0 960 0 1 4170
box -8 -3 46 105
use FILL  FILL_757
timestamp 1680363874
transform 1 0 1000 0 1 4170
box -8 -3 16 105
use FILL  FILL_759
timestamp 1680363874
transform 1 0 1008 0 1 4170
box -8 -3 16 105
use FILL  FILL_761
timestamp 1680363874
transform 1 0 1016 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_72
timestamp 1680363874
transform 1 0 1024 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_74
timestamp 1680363874
transform 1 0 1064 0 1 4170
box -8 -3 46 105
use FILL  FILL_763
timestamp 1680363874
transform 1 0 1104 0 1 4170
box -8 -3 16 105
use FILL  FILL_770
timestamp 1680363874
transform 1 0 1112 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1680363874
transform -1 0 1216 0 1 4170
box -8 -3 104 105
use FILL  FILL_771
timestamp 1680363874
transform 1 0 1216 0 1 4170
box -8 -3 16 105
use FILL  FILL_772
timestamp 1680363874
transform 1 0 1224 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_75
timestamp 1680363874
transform 1 0 1232 0 1 4170
box -8 -3 46 105
use FILL  FILL_773
timestamp 1680363874
transform 1 0 1272 0 1 4170
box -8 -3 16 105
use FILL  FILL_774
timestamp 1680363874
transform 1 0 1280 0 1 4170
box -8 -3 16 105
use FILL  FILL_775
timestamp 1680363874
transform 1 0 1288 0 1 4170
box -8 -3 16 105
use FILL  FILL_776
timestamp 1680363874
transform 1 0 1296 0 1 4170
box -8 -3 16 105
use FILL  FILL_782
timestamp 1680363874
transform 1 0 1304 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_77
timestamp 1680363874
transform 1 0 1312 0 1 4170
box -8 -3 46 105
use FILL  FILL_784
timestamp 1680363874
transform 1 0 1352 0 1 4170
box -8 -3 16 105
use FILL  FILL_785
timestamp 1680363874
transform 1 0 1360 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_82
timestamp 1680363874
transform -1 0 1384 0 1 4170
box -9 -3 26 105
use FILL  FILL_786
timestamp 1680363874
transform 1 0 1384 0 1 4170
box -8 -3 16 105
use FILL  FILL_787
timestamp 1680363874
transform 1 0 1392 0 1 4170
box -8 -3 16 105
use FILL  FILL_788
timestamp 1680363874
transform 1 0 1400 0 1 4170
box -8 -3 16 105
use FILL  FILL_789
timestamp 1680363874
transform 1 0 1408 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_83
timestamp 1680363874
transform -1 0 1432 0 1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1680363874
transform -1 0 1528 0 1 4170
box -8 -3 104 105
use FILL  FILL_790
timestamp 1680363874
transform 1 0 1528 0 1 4170
box -8 -3 16 105
use FILL  FILL_791
timestamp 1680363874
transform 1 0 1536 0 1 4170
box -8 -3 16 105
use FILL  FILL_792
timestamp 1680363874
transform 1 0 1544 0 1 4170
box -8 -3 16 105
use FILL  FILL_793
timestamp 1680363874
transform 1 0 1552 0 1 4170
box -8 -3 16 105
use FILL  FILL_794
timestamp 1680363874
transform 1 0 1560 0 1 4170
box -8 -3 16 105
use FILL  FILL_795
timestamp 1680363874
transform 1 0 1568 0 1 4170
box -8 -3 16 105
use FILL  FILL_796
timestamp 1680363874
transform 1 0 1576 0 1 4170
box -8 -3 16 105
use FILL  FILL_797
timestamp 1680363874
transform 1 0 1584 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1680363874
transform 1 0 1592 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_84
timestamp 1680363874
transform -1 0 1704 0 1 4170
box -9 -3 26 105
use FILL  FILL_798
timestamp 1680363874
transform 1 0 1704 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1010
timestamp 1680363874
transform 1 0 1732 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_85
timestamp 1680363874
transform 1 0 1712 0 1 4170
box -9 -3 26 105
use FILL  FILL_799
timestamp 1680363874
transform 1 0 1728 0 1 4170
box -8 -3 16 105
use FILL  FILL_800
timestamp 1680363874
transform 1 0 1736 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1011
timestamp 1680363874
transform 1 0 1788 0 1 4175
box -3 -3 3 3
use AOI22X1  AOI22X1_45
timestamp 1680363874
transform -1 0 1784 0 1 4170
box -8 -3 46 105
use FILL  FILL_801
timestamp 1680363874
transform 1 0 1784 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_46
timestamp 1680363874
transform -1 0 1832 0 1 4170
box -8 -3 46 105
use FILL  FILL_802
timestamp 1680363874
transform 1 0 1832 0 1 4170
box -8 -3 16 105
use FILL  FILL_803
timestamp 1680363874
transform 1 0 1840 0 1 4170
box -8 -3 16 105
use FILL  FILL_804
timestamp 1680363874
transform 1 0 1848 0 1 4170
box -8 -3 16 105
use FILL  FILL_813
timestamp 1680363874
transform 1 0 1856 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_47
timestamp 1680363874
transform -1 0 1904 0 1 4170
box -8 -3 46 105
use FILL  FILL_814
timestamp 1680363874
transform 1 0 1904 0 1 4170
box -8 -3 16 105
use FILL  FILL_815
timestamp 1680363874
transform 1 0 1912 0 1 4170
box -8 -3 16 105
use FILL  FILL_816
timestamp 1680363874
transform 1 0 1920 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_48
timestamp 1680363874
transform 1 0 1928 0 1 4170
box -8 -3 46 105
use FILL  FILL_821
timestamp 1680363874
transform 1 0 1968 0 1 4170
box -8 -3 16 105
use FILL  FILL_822
timestamp 1680363874
transform 1 0 1976 0 1 4170
box -8 -3 16 105
use FILL  FILL_823
timestamp 1680363874
transform 1 0 1984 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1012
timestamp 1680363874
transform 1 0 2020 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_87
timestamp 1680363874
transform 1 0 1992 0 1 4170
box -9 -3 26 105
use FILL  FILL_824
timestamp 1680363874
transform 1 0 2008 0 1 4170
box -8 -3 16 105
use FILL  FILL_825
timestamp 1680363874
transform 1 0 2016 0 1 4170
box -8 -3 16 105
use FILL  FILL_826
timestamp 1680363874
transform 1 0 2024 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1013
timestamp 1680363874
transform 1 0 2044 0 1 4175
box -3 -3 3 3
use FILL  FILL_827
timestamp 1680363874
transform 1 0 2032 0 1 4170
box -8 -3 16 105
use FILL  FILL_830
timestamp 1680363874
transform 1 0 2040 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1014
timestamp 1680363874
transform 1 0 2084 0 1 4175
box -3 -3 3 3
use AOI22X1  AOI22X1_49
timestamp 1680363874
transform -1 0 2088 0 1 4170
box -8 -3 46 105
use FILL  FILL_831
timestamp 1680363874
transform 1 0 2088 0 1 4170
box -8 -3 16 105
use FILL  FILL_832
timestamp 1680363874
transform 1 0 2096 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_88
timestamp 1680363874
transform 1 0 2104 0 1 4170
box -9 -3 26 105
use FILL  FILL_833
timestamp 1680363874
transform 1 0 2120 0 1 4170
box -8 -3 16 105
use FILL  FILL_834
timestamp 1680363874
transform 1 0 2128 0 1 4170
box -8 -3 16 105
use FILL  FILL_835
timestamp 1680363874
transform 1 0 2136 0 1 4170
box -8 -3 16 105
use FILL  FILL_836
timestamp 1680363874
transform 1 0 2144 0 1 4170
box -8 -3 16 105
use FILL  FILL_837
timestamp 1680363874
transform 1 0 2152 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1680363874
transform -1 0 2200 0 1 4170
box -8 -3 46 105
use FILL  FILL_838
timestamp 1680363874
transform 1 0 2200 0 1 4170
box -8 -3 16 105
use FILL  FILL_839
timestamp 1680363874
transform 1 0 2208 0 1 4170
box -8 -3 16 105
use FILL  FILL_840
timestamp 1680363874
transform 1 0 2216 0 1 4170
box -8 -3 16 105
use FILL  FILL_841
timestamp 1680363874
transform 1 0 2224 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_81
timestamp 1680363874
transform 1 0 2232 0 1 4170
box -8 -3 46 105
use FILL  FILL_842
timestamp 1680363874
transform 1 0 2272 0 1 4170
box -8 -3 16 105
use FILL  FILL_847
timestamp 1680363874
transform 1 0 2280 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1680363874
transform 1 0 2288 0 1 4170
box -8 -3 104 105
use FILL  FILL_848
timestamp 1680363874
transform 1 0 2384 0 1 4170
box -8 -3 16 105
use FILL  FILL_849
timestamp 1680363874
transform 1 0 2392 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_90
timestamp 1680363874
transform 1 0 2400 0 1 4170
box -9 -3 26 105
use FILL  FILL_850
timestamp 1680363874
transform 1 0 2416 0 1 4170
box -8 -3 16 105
use FILL  FILL_859
timestamp 1680363874
transform 1 0 2424 0 1 4170
box -8 -3 16 105
use FILL  FILL_860
timestamp 1680363874
transform 1 0 2432 0 1 4170
box -8 -3 16 105
use FILL  FILL_861
timestamp 1680363874
transform 1 0 2440 0 1 4170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1680363874
transform 1 0 2448 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_91
timestamp 1680363874
transform -1 0 2472 0 1 4170
box -9 -3 26 105
use FILL  FILL_863
timestamp 1680363874
transform 1 0 2472 0 1 4170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1680363874
transform 1 0 2480 0 1 4170
box -8 -3 16 105
use FILL  FILL_865
timestamp 1680363874
transform 1 0 2488 0 1 4170
box -8 -3 16 105
use FILL  FILL_866
timestamp 1680363874
transform 1 0 2496 0 1 4170
box -8 -3 16 105
use FILL  FILL_867
timestamp 1680363874
transform 1 0 2504 0 1 4170
box -8 -3 16 105
use FILL  FILL_868
timestamp 1680363874
transform 1 0 2512 0 1 4170
box -8 -3 16 105
use FILL  FILL_869
timestamp 1680363874
transform 1 0 2520 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1680363874
transform 1 0 2528 0 1 4170
box -8 -3 104 105
use FILL  FILL_870
timestamp 1680363874
transform 1 0 2624 0 1 4170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1680363874
transform 1 0 2632 0 1 4170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1680363874
transform 1 0 2640 0 1 4170
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1680363874
transform 1 0 2648 0 1 4170
box -8 -3 40 105
use FILL  FILL_883
timestamp 1680363874
transform 1 0 2680 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_93
timestamp 1680363874
transform -1 0 2704 0 1 4170
box -9 -3 26 105
use FILL  FILL_884
timestamp 1680363874
transform 1 0 2704 0 1 4170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1680363874
transform 1 0 2712 0 1 4170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1680363874
transform 1 0 2720 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1680363874
transform -1 0 2768 0 1 4170
box -8 -3 46 105
use FILL  FILL_887
timestamp 1680363874
transform 1 0 2768 0 1 4170
box -8 -3 16 105
use FILL  FILL_892
timestamp 1680363874
transform 1 0 2776 0 1 4170
box -8 -3 16 105
use FILL  FILL_894
timestamp 1680363874
transform 1 0 2784 0 1 4170
box -8 -3 16 105
use FILL  FILL_895
timestamp 1680363874
transform 1 0 2792 0 1 4170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1680363874
transform 1 0 2800 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_94
timestamp 1680363874
transform 1 0 2808 0 1 4170
box -9 -3 26 105
use FILL  FILL_897
timestamp 1680363874
transform 1 0 2824 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_53
timestamp 1680363874
transform 1 0 2832 0 1 4170
box -8 -3 46 105
use M3_M2  M3_M2_1015
timestamp 1680363874
transform 1 0 2964 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_101
timestamp 1680363874
transform -1 0 2968 0 1 4170
box -8 -3 104 105
use FILL  FILL_898
timestamp 1680363874
transform 1 0 2968 0 1 4170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1680363874
transform 1 0 2976 0 1 4170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1680363874
transform 1 0 2984 0 1 4170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1680363874
transform 1 0 2992 0 1 4170
box -8 -3 16 105
use FILL  FILL_909
timestamp 1680363874
transform 1 0 3000 0 1 4170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1680363874
transform 1 0 3008 0 1 4170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1680363874
transform 1 0 3016 0 1 4170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1680363874
transform 1 0 3024 0 1 4170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1680363874
transform 1 0 3032 0 1 4170
box -8 -3 16 105
use FILL  FILL_917
timestamp 1680363874
transform 1 0 3040 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_95
timestamp 1680363874
transform 1 0 3048 0 1 4170
box -9 -3 26 105
use FILL  FILL_919
timestamp 1680363874
transform 1 0 3064 0 1 4170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1680363874
transform 1 0 3072 0 1 4170
box -8 -3 16 105
use FILL  FILL_921
timestamp 1680363874
transform 1 0 3080 0 1 4170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1680363874
transform 1 0 3088 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1680363874
transform -1 0 3192 0 1 4170
box -8 -3 104 105
use FILL  FILL_924
timestamp 1680363874
transform 1 0 3192 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_96
timestamp 1680363874
transform -1 0 3216 0 1 4170
box -9 -3 26 105
use FILL  FILL_925
timestamp 1680363874
transform 1 0 3216 0 1 4170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1680363874
transform 1 0 3224 0 1 4170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1680363874
transform 1 0 3232 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_54
timestamp 1680363874
transform -1 0 3280 0 1 4170
box -8 -3 46 105
use FILL  FILL_928
timestamp 1680363874
transform 1 0 3280 0 1 4170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1680363874
transform 1 0 3288 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_55
timestamp 1680363874
transform 1 0 3296 0 1 4170
box -8 -3 46 105
use FILL  FILL_930
timestamp 1680363874
transform 1 0 3336 0 1 4170
box -8 -3 16 105
use FILL  FILL_931
timestamp 1680363874
transform 1 0 3344 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_97
timestamp 1680363874
transform 1 0 3352 0 1 4170
box -9 -3 26 105
use FILL  FILL_932
timestamp 1680363874
transform 1 0 3368 0 1 4170
box -8 -3 16 105
use FILL  FILL_933
timestamp 1680363874
transform 1 0 3376 0 1 4170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1680363874
transform 1 0 3384 0 1 4170
box -8 -3 16 105
use FILL  FILL_935
timestamp 1680363874
transform 1 0 3392 0 1 4170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1680363874
transform 1 0 3400 0 1 4170
box -8 -3 16 105
use FILL  FILL_937
timestamp 1680363874
transform 1 0 3408 0 1 4170
box -8 -3 16 105
use FILL  FILL_938
timestamp 1680363874
transform 1 0 3416 0 1 4170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1680363874
transform 1 0 3424 0 1 4170
box -8 -3 16 105
use FILL  FILL_940
timestamp 1680363874
transform 1 0 3432 0 1 4170
box -8 -3 16 105
use FILL  FILL_941
timestamp 1680363874
transform 1 0 3440 0 1 4170
box -8 -3 16 105
use FILL  FILL_942
timestamp 1680363874
transform 1 0 3448 0 1 4170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1680363874
transform 1 0 3456 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1680363874
transform 1 0 3464 0 1 4170
box -8 -3 104 105
use FILL  FILL_954
timestamp 1680363874
transform 1 0 3560 0 1 4170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1680363874
transform 1 0 3568 0 1 4170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1680363874
transform 1 0 3576 0 1 4170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1680363874
transform 1 0 3584 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_100
timestamp 1680363874
transform 1 0 3592 0 1 4170
box -9 -3 26 105
use OAI22X1  OAI22X1_85
timestamp 1680363874
transform 1 0 3608 0 1 4170
box -8 -3 46 105
use FILL  FILL_958
timestamp 1680363874
transform 1 0 3648 0 1 4170
box -8 -3 16 105
use FILL  FILL_959
timestamp 1680363874
transform 1 0 3656 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1016
timestamp 1680363874
transform 1 0 3708 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_107
timestamp 1680363874
transform 1 0 3664 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_101
timestamp 1680363874
transform -1 0 3776 0 1 4170
box -9 -3 26 105
use FILL  FILL_960
timestamp 1680363874
transform 1 0 3776 0 1 4170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1680363874
transform 1 0 3784 0 1 4170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1680363874
transform 1 0 3792 0 1 4170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1680363874
transform 1 0 3800 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_57
timestamp 1680363874
transform -1 0 3848 0 1 4170
box -8 -3 46 105
use FILL  FILL_964
timestamp 1680363874
transform 1 0 3848 0 1 4170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1680363874
transform 1 0 3856 0 1 4170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1680363874
transform 1 0 3864 0 1 4170
box -8 -3 16 105
use FILL  FILL_984
timestamp 1680363874
transform 1 0 3872 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_86
timestamp 1680363874
transform 1 0 3880 0 1 4170
box -8 -3 46 105
use FILL  FILL_986
timestamp 1680363874
transform 1 0 3920 0 1 4170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1680363874
transform 1 0 3928 0 1 4170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1680363874
transform 1 0 3936 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1680363874
transform -1 0 4040 0 1 4170
box -8 -3 104 105
use FILL  FILL_996
timestamp 1680363874
transform 1 0 4040 0 1 4170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1680363874
transform 1 0 4048 0 1 4170
box -8 -3 16 105
use FILL  FILL_998
timestamp 1680363874
transform 1 0 4056 0 1 4170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1680363874
transform 1 0 4064 0 1 4170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1680363874
transform 1 0 4072 0 1 4170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1680363874
transform 1 0 4080 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_102
timestamp 1680363874
transform -1 0 4104 0 1 4170
box -9 -3 26 105
use FILL  FILL_1002
timestamp 1680363874
transform 1 0 4104 0 1 4170
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1680363874
transform 1 0 4112 0 1 4170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1680363874
transform 1 0 4120 0 1 4170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1680363874
transform 1 0 4128 0 1 4170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1680363874
transform 1 0 4136 0 1 4170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1680363874
transform 1 0 4144 0 1 4170
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1680363874
transform 1 0 4152 0 1 4170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1680363874
transform 1 0 4160 0 1 4170
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1680363874
transform 1 0 4168 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_60
timestamp 1680363874
transform -1 0 4216 0 1 4170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1680363874
transform 1 0 4216 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_103
timestamp 1680363874
transform -1 0 4328 0 1 4170
box -9 -3 26 105
use FILL  FILL_1011
timestamp 1680363874
transform 1 0 4328 0 1 4170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1680363874
transform 1 0 4336 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_61
timestamp 1680363874
transform -1 0 4384 0 1 4170
box -8 -3 46 105
use FILL  FILL_1013
timestamp 1680363874
transform 1 0 4384 0 1 4170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1680363874
transform 1 0 4392 0 1 4170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1680363874
transform 1 0 4400 0 1 4170
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1680363874
transform 1 0 4408 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_62
timestamp 1680363874
transform 1 0 4416 0 1 4170
box -8 -3 46 105
use FILL  FILL_1026
timestamp 1680363874
transform 1 0 4456 0 1 4170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1680363874
transform 1 0 4464 0 1 4170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1680363874
transform 1 0 4472 0 1 4170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1680363874
transform 1 0 4480 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_88
timestamp 1680363874
transform 1 0 4488 0 1 4170
box -8 -3 46 105
use FILL  FILL_1034
timestamp 1680363874
transform 1 0 4528 0 1 4170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1680363874
transform 1 0 4536 0 1 4170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1680363874
transform 1 0 4544 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_64
timestamp 1680363874
transform 1 0 4552 0 1 4170
box -8 -3 46 105
use FILL  FILL_1040
timestamp 1680363874
transform 1 0 4592 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_65
timestamp 1680363874
transform -1 0 4640 0 1 4170
box -8 -3 46 105
use FILL  FILL_1041
timestamp 1680363874
transform 1 0 4640 0 1 4170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1680363874
transform 1 0 4648 0 1 4170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1680363874
transform 1 0 4656 0 1 4170
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1680363874
transform 1 0 4664 0 1 4170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1680363874
transform 1 0 4672 0 1 4170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1680363874
transform 1 0 4680 0 1 4170
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1680363874
transform 1 0 4688 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1680363874
transform -1 0 4792 0 1 4170
box -8 -3 104 105
use FILL  FILL_1059
timestamp 1680363874
transform 1 0 4792 0 1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_11
timestamp 1680363874
transform 1 0 4827 0 1 4170
box -10 -3 10 3
use M3_M2  M3_M2_1052
timestamp 1680363874
transform 1 0 132 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1680363874
transform 1 0 68 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1192
timestamp 1680363874
transform 1 0 156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1680363874
transform 1 0 172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1680363874
transform 1 0 68 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1680363874
transform 1 0 132 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1680363874
transform 1 0 180 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1680363874
transform 1 0 188 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1680363874
transform 1 0 220 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1680363874
transform 1 0 212 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1195
timestamp 1680363874
transform 1 0 220 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1680363874
transform 1 0 236 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1680363874
transform 1 0 244 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1680363874
transform 1 0 212 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1680363874
transform 1 0 228 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1174
timestamp 1680363874
transform 1 0 228 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1680363874
transform 1 0 316 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1198
timestamp 1680363874
transform 1 0 268 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1680363874
transform 1 0 252 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1680363874
transform 1 0 316 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1680363874
transform 1 0 260 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1199
timestamp 1680363874
transform 1 0 372 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1680363874
transform 1 0 412 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1680363874
transform 1 0 412 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1680363874
transform 1 0 428 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1680363874
transform 1 0 404 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1680363874
transform 1 0 420 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1141
timestamp 1680363874
transform 1 0 404 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1202
timestamp 1680363874
transform 1 0 484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1680363874
transform 1 0 500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1680363874
transform 1 0 508 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1680363874
transform 1 0 476 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1680363874
transform 1 0 476 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1680363874
transform 1 0 508 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1680363874
transform 1 0 564 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1680363874
transform 1 0 556 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1680363874
transform 1 0 540 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1680363874
transform 1 0 556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1680363874
transform 1 0 572 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1680363874
transform 1 0 580 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1680363874
transform 1 0 540 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1680363874
transform 1 0 548 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1680363874
transform 1 0 564 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1123
timestamp 1680363874
transform 1 0 572 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1680363874
transform 1 0 548 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1680363874
transform 1 0 580 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1680363874
transform 1 0 588 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1680363874
transform 1 0 604 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1680363874
transform 1 0 652 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1680363874
transform 1 0 628 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1680363874
transform 1 0 644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1680363874
transform 1 0 652 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1680363874
transform 1 0 620 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1680363874
transform 1 0 636 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1124
timestamp 1680363874
transform 1 0 644 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1308
timestamp 1680363874
transform 1 0 652 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1179
timestamp 1680363874
transform 1 0 652 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1211
timestamp 1680363874
transform 1 0 684 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1680363874
transform 1 0 708 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1104
timestamp 1680363874
transform 1 0 716 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1680363874
transform 1 0 724 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1680363874
transform 1 0 732 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1680363874
transform 1 0 700 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1680363874
transform 1 0 708 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1310
timestamp 1680363874
transform 1 0 716 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1144
timestamp 1680363874
transform 1 0 700 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1680363874
transform 1 0 740 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1680363874
transform 1 0 732 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1680363874
transform 1 0 788 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1680363874
transform 1 0 772 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1215
timestamp 1680363874
transform 1 0 788 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1680363874
transform 1 0 772 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1127
timestamp 1680363874
transform 1 0 780 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1680363874
transform 1 0 804 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1411
timestamp 1680363874
transform 1 0 804 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1020
timestamp 1680363874
transform 1 0 820 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1680363874
transform 1 0 836 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1680363874
transform 1 0 860 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1680363874
transform 1 0 852 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1216
timestamp 1680363874
transform 1 0 852 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1680363874
transform 1 0 860 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1680363874
transform 1 0 868 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1680363874
transform 1 0 908 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1313
timestamp 1680363874
transform 1 0 892 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1180
timestamp 1680363874
transform 1 0 892 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1680363874
transform 1 0 924 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1680363874
transform 1 0 924 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1680363874
transform 1 0 932 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1038
timestamp 1680363874
transform 1 0 996 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1680363874
transform 1 0 972 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1219
timestamp 1680363874
transform 1 0 964 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1680363874
transform 1 0 980 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1107
timestamp 1680363874
transform 1 0 988 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1221
timestamp 1680363874
transform 1 0 996 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1680363874
transform 1 0 972 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1128
timestamp 1680363874
transform 1 0 980 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1315
timestamp 1680363874
transform 1 0 988 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1063
timestamp 1680363874
transform 1 0 1012 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1222
timestamp 1680363874
transform 1 0 1028 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1680363874
transform 1 0 1044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1680363874
transform 1 0 1020 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1680363874
transform 1 0 1052 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1317
timestamp 1680363874
transform 1 0 1052 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1181
timestamp 1680363874
transform 1 0 1044 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1224
timestamp 1680363874
transform 1 0 1100 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1109
timestamp 1680363874
transform 1 0 1108 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1680363874
transform 1 0 1100 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1680363874
transform 1 0 1132 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1680363874
transform 1 0 1204 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1680363874
transform 1 0 1188 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1225
timestamp 1680363874
transform 1 0 1132 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1680363874
transform 1 0 1148 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1680363874
transform 1 0 1164 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1680363874
transform 1 0 1116 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1680363874
transform 1 0 1140 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1146
timestamp 1680363874
transform 1 0 1116 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1680363874
transform 1 0 1148 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1320
timestamp 1680363874
transform 1 0 1188 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1182
timestamp 1680363874
transform 1 0 1140 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1680363874
transform 1 0 1188 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1680363874
transform 1 0 1300 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1228
timestamp 1680363874
transform 1 0 1292 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1680363874
transform 1 0 1276 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1680363874
transform 1 0 1284 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1680363874
transform 1 0 1284 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1323
timestamp 1680363874
transform 1 0 1300 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1680363874
transform 1 0 1308 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1205
timestamp 1680363874
transform 1 0 1308 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1680363874
transform 1 0 1324 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1680363874
transform 1 0 1348 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1680363874
transform 1 0 1332 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1230
timestamp 1680363874
transform 1 0 1332 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1110
timestamp 1680363874
transform 1 0 1340 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1231
timestamp 1680363874
transform 1 0 1348 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1680363874
transform 1 0 1324 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1680363874
transform 1 0 1340 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1130
timestamp 1680363874
transform 1 0 1348 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1680363874
transform 1 0 1324 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1680363874
transform 1 0 1340 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1680363874
transform 1 0 1372 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1680363874
transform 1 0 1444 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1680363874
transform 1 0 1396 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1232
timestamp 1680363874
transform 1 0 1444 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1680363874
transform 1 0 1364 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1680363874
transform 1 0 1396 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1068
timestamp 1680363874
transform 1 0 1476 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1680363874
transform 1 0 1516 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1233
timestamp 1680363874
transform 1 0 1476 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1680363874
transform 1 0 1500 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1680363874
transform 1 0 1588 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1234
timestamp 1680363874
transform 1 0 1572 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1680363874
transform 1 0 1588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1680363874
transform 1 0 1500 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1680363874
transform 1 0 1556 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1680363874
transform 1 0 1564 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1680363874
transform 1 0 1564 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1680363874
transform 1 0 1588 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1331
timestamp 1680363874
transform 1 0 1628 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1680363874
transform 1 0 1668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1680363874
transform 1 0 1700 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1680363874
transform 1 0 1724 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1680363874
transform 1 0 1788 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1680363874
transform 1 0 1804 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1334
timestamp 1680363874
transform 1 0 1804 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1680363874
transform 1 0 1852 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1238
timestamp 1680363874
transform 1 0 1828 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1680363874
transform 1 0 1844 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1680363874
transform 1 0 1852 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1680363874
transform 1 0 1820 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1680363874
transform 1 0 1836 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1150
timestamp 1680363874
transform 1 0 1844 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1680363874
transform 1 0 1820 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1680363874
transform 1 0 1860 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1241
timestamp 1680363874
transform 1 0 1900 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1680363874
transform 1 0 1892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1680363874
transform 1 0 1908 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1680363874
transform 1 0 1908 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1680363874
transform 1 0 1892 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1680363874
transform 1 0 1908 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1242
timestamp 1680363874
transform 1 0 1932 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1680363874
transform 1 0 2020 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1680363874
transform 1 0 1940 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1680363874
transform 1 0 1996 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1133
timestamp 1680363874
transform 1 0 2020 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1680363874
transform 1 0 2036 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1680363874
transform 1 0 2060 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1680363874
transform 1 0 2244 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1680363874
transform 1 0 2172 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1680363874
transform 1 0 2252 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1680363874
transform 1 0 2060 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1680363874
transform 1 0 2148 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1680363874
transform 1 0 2156 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1680363874
transform 1 0 2172 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1113
timestamp 1680363874
transform 1 0 2196 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1680363874
transform 1 0 2260 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1680363874
transform 1 0 2108 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1680363874
transform 1 0 2148 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1680363874
transform 1 0 2156 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1680363874
transform 1 0 2196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1680363874
transform 1 0 2252 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1152
timestamp 1680363874
transform 1 0 2060 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1680363874
transform 1 0 2148 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1680363874
transform 1 0 2204 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1680363874
transform 1 0 2252 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1680363874
transform 1 0 2268 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1680363874
transform 1 0 2284 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1680363874
transform 1 0 2316 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1680363874
transform 1 0 2300 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1680363874
transform 1 0 2300 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1247
timestamp 1680363874
transform 1 0 2308 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1680363874
transform 1 0 2300 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1680363874
transform 1 0 2316 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1074
timestamp 1680363874
transform 1 0 2388 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1248
timestamp 1680363874
transform 1 0 2372 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1680363874
transform 1 0 2388 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1680363874
transform 1 0 2396 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1680363874
transform 1 0 2364 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1680363874
transform 1 0 2380 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1026
timestamp 1680363874
transform 1 0 2476 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1251
timestamp 1680363874
transform 1 0 2436 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1116
timestamp 1680363874
transform 1 0 2524 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1350
timestamp 1680363874
transform 1 0 2460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1680363874
transform 1 0 2516 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1680363874
transform 1 0 2524 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1154
timestamp 1680363874
transform 1 0 2436 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1680363874
transform 1 0 2556 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1252
timestamp 1680363874
transform 1 0 2556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1680363874
transform 1 0 2548 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1680363874
transform 1 0 2540 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1680363874
transform 1 0 2548 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1253
timestamp 1680363874
transform 1 0 2580 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1680363874
transform 1 0 2572 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1076
timestamp 1680363874
transform 1 0 2636 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1680363874
transform 1 0 2740 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1254
timestamp 1680363874
transform 1 0 2660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1680363874
transform 1 0 2692 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1680363874
transform 1 0 2740 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1027
timestamp 1680363874
transform 1 0 2788 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1680363874
transform 1 0 2868 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1255
timestamp 1680363874
transform 1 0 2796 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1117
timestamp 1680363874
transform 1 0 2844 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1680363874
transform 1 0 2884 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1256
timestamp 1680363874
transform 1 0 2884 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1680363874
transform 1 0 2836 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1680363874
transform 1 0 2876 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1029
timestamp 1680363874
transform 1 0 2940 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1257
timestamp 1680363874
transform 1 0 2924 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1680363874
transform 1 0 2940 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1680363874
transform 1 0 2916 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1188
timestamp 1680363874
transform 1 0 2916 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1680363874
transform 1 0 2988 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1680363874
transform 1 0 3004 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1680363874
transform 1 0 2980 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1680363874
transform 1 0 2980 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1361
timestamp 1680363874
transform 1 0 2996 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1680363874
transform 1 0 3012 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1157
timestamp 1680363874
transform 1 0 3012 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1680363874
transform 1 0 2996 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1680363874
transform 1 0 3044 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1680363874
transform 1 0 3068 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1261
timestamp 1680363874
transform 1 0 3044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1680363874
transform 1 0 3052 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1190
timestamp 1680363874
transform 1 0 3036 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1680363874
transform 1 0 3052 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1680363874
transform 1 0 3076 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1680363874
transform 1 0 3060 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1680363874
transform 1 0 3092 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1680363874
transform 1 0 3084 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1680363874
transform 1 0 3092 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1680363874
transform 1 0 3108 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1209
timestamp 1680363874
transform 1 0 3108 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1680363874
transform 1 0 3140 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1366
timestamp 1680363874
transform 1 0 3140 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1680363874
transform 1 0 3148 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1191
timestamp 1680363874
transform 1 0 3148 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1680363874
transform 1 0 3252 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1680363874
transform 1 0 3252 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1137
timestamp 1680363874
transform 1 0 3212 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1368
timestamp 1680363874
transform 1 0 3228 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1158
timestamp 1680363874
transform 1 0 3228 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1680363874
transform 1 0 3236 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1680363874
transform 1 0 3268 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1369
timestamp 1680363874
transform 1 0 3268 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1159
timestamp 1680363874
transform 1 0 3268 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1370
timestamp 1680363874
transform 1 0 3292 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1030
timestamp 1680363874
transform 1 0 3332 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1680363874
transform 1 0 3356 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1680363874
transform 1 0 3420 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1265
timestamp 1680363874
transform 1 0 3308 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1680363874
transform 1 0 3316 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1680363874
transform 1 0 3332 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1160
timestamp 1680363874
transform 1 0 3300 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1680363874
transform 1 0 3300 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1680363874
transform 1 0 3340 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1268
timestamp 1680363874
transform 1 0 3356 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1680363874
transform 1 0 3324 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1680363874
transform 1 0 3340 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1680363874
transform 1 0 3404 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1680363874
transform 1 0 3436 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1680363874
transform 1 0 3444 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1161
timestamp 1680363874
transform 1 0 3340 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1680363874
transform 1 0 3404 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1680363874
transform 1 0 3444 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1680363874
transform 1 0 3316 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1680363874
transform 1 0 3348 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1680363874
transform 1 0 3436 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1680363874
transform 1 0 3476 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1269
timestamp 1680363874
transform 1 0 3484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1680363874
transform 1 0 3492 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1121
timestamp 1680363874
transform 1 0 3516 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1680363874
transform 1 0 3532 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1680363874
transform 1 0 3532 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1271
timestamp 1680363874
transform 1 0 3532 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1680363874
transform 1 0 3484 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1680363874
transform 1 0 3500 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1680363874
transform 1 0 3516 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1680363874
transform 1 0 3524 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1164
timestamp 1680363874
transform 1 0 3484 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1680363874
transform 1 0 3492 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1680363874
transform 1 0 3524 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1680363874
transform 1 0 3516 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1272
timestamp 1680363874
transform 1 0 3548 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1086
timestamp 1680363874
transform 1 0 3596 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1273
timestamp 1680363874
transform 1 0 3596 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1680363874
transform 1 0 3572 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1680363874
transform 1 0 3588 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1680363874
transform 1 0 3572 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1680363874
transform 1 0 3604 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1382
timestamp 1680363874
transform 1 0 3644 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1196
timestamp 1680363874
transform 1 0 3644 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1680363874
transform 1 0 3636 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1680363874
transform 1 0 3660 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1274
timestamp 1680363874
transform 1 0 3660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1680363874
transform 1 0 3684 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1680363874
transform 1 0 3740 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1197
timestamp 1680363874
transform 1 0 3692 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1680363874
transform 1 0 3676 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1680363874
transform 1 0 3764 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1275
timestamp 1680363874
transform 1 0 3764 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1680363874
transform 1 0 3796 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1680363874
transform 1 0 3844 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1089
timestamp 1680363874
transform 1 0 3868 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1680363874
transform 1 0 3908 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1680363874
transform 1 0 3908 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1387
timestamp 1680363874
transform 1 0 3916 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1680363874
transform 1 0 3932 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1091
timestamp 1680363874
transform 1 0 4004 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1277
timestamp 1680363874
transform 1 0 4004 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1680363874
transform 1 0 3988 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1032
timestamp 1680363874
transform 1 0 4028 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1680363874
transform 1 0 4044 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1680363874
transform 1 0 4172 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1680363874
transform 1 0 4228 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1680363874
transform 1 0 4268 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1680363874
transform 1 0 4204 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1680363874
transform 1 0 4172 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1680363874
transform 1 0 4196 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1278
timestamp 1680363874
transform 1 0 4028 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1680363874
transform 1 0 4044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1680363874
transform 1 0 4132 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1680363874
transform 1 0 4148 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1680363874
transform 1 0 4164 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1680363874
transform 1 0 4172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1680363874
transform 1 0 4012 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1680363874
transform 1 0 4076 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1680363874
transform 1 0 4124 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1680363874
transform 1 0 4140 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1680363874
transform 1 0 4156 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1680363874
transform 1 0 4268 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1680363874
transform 1 0 4180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1680363874
transform 1 0 4188 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1680363874
transform 1 0 4220 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1168
timestamp 1680363874
transform 1 0 4180 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1680363874
transform 1 0 4220 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1680363874
transform 1 0 4308 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1680363874
transform 1 0 4324 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1680363874
transform 1 0 4348 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1285
timestamp 1680363874
transform 1 0 4308 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1122
timestamp 1680363874
transform 1 0 4388 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1397
timestamp 1680363874
transform 1 0 4356 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1170
timestamp 1680363874
transform 1 0 4356 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1680363874
transform 1 0 4388 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1413
timestamp 1680363874
transform 1 0 4396 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1201
timestamp 1680363874
transform 1 0 4356 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1680363874
transform 1 0 4380 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1680363874
transform 1 0 4420 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1680363874
transform 1 0 4412 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1680363874
transform 1 0 4444 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1286
timestamp 1680363874
transform 1 0 4428 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1680363874
transform 1 0 4444 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1680363874
transform 1 0 4412 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1680363874
transform 1 0 4420 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1680363874
transform 1 0 4436 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1680363874
transform 1 0 4452 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1680363874
transform 1 0 4460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1680363874
transform 1 0 4412 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1198
timestamp 1680363874
transform 1 0 4420 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1680363874
transform 1 0 4476 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1403
timestamp 1680363874
transform 1 0 4500 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1680363874
transform 1 0 4524 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1680363874
transform 1 0 4532 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1680363874
transform 1 0 4556 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1680363874
transform 1 0 4604 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1680363874
transform 1 0 4636 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1289
timestamp 1680363874
transform 1 0 4596 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1680363874
transform 1 0 4604 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1680363874
transform 1 0 4620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1680363874
transform 1 0 4628 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1680363874
transform 1 0 4588 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1680363874
transform 1 0 4604 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1406
timestamp 1680363874
transform 1 0 4612 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1680363874
transform 1 0 4628 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1203
timestamp 1680363874
transform 1 0 4628 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1680363874
transform 1 0 4788 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1293
timestamp 1680363874
transform 1 0 4708 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1680363874
transform 1 0 4692 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1680363874
transform 1 0 4732 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1140
timestamp 1680363874
transform 1 0 4756 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1680363874
transform 1 0 4788 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1172
timestamp 1680363874
transform 1 0 4692 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1680363874
transform 1 0 4732 0 1 4115
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_12
timestamp 1680363874
transform 1 0 24 0 1 4070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_83
timestamp 1680363874
transform -1 0 168 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_76
timestamp 1680363874
transform 1 0 168 0 -1 4170
box -9 -3 26 105
use FILL  FILL_692
timestamp 1680363874
transform 1 0 184 0 -1 4170
box -8 -3 16 105
use FILL  FILL_693
timestamp 1680363874
transform 1 0 192 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_61
timestamp 1680363874
transform 1 0 200 0 -1 4170
box -8 -3 46 105
use INVX2  INVX2_77
timestamp 1680363874
transform 1 0 240 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1680363874
transform 1 0 256 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_78
timestamp 1680363874
transform 1 0 352 0 -1 4170
box -9 -3 26 105
use FILL  FILL_694
timestamp 1680363874
transform 1 0 368 0 -1 4170
box -8 -3 16 105
use FILL  FILL_695
timestamp 1680363874
transform 1 0 376 0 -1 4170
box -8 -3 16 105
use FILL  FILL_696
timestamp 1680363874
transform 1 0 384 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_62
timestamp 1680363874
transform 1 0 392 0 -1 4170
box -8 -3 46 105
use FILL  FILL_697
timestamp 1680363874
transform 1 0 432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_699
timestamp 1680363874
transform 1 0 440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_706
timestamp 1680363874
transform 1 0 448 0 -1 4170
box -8 -3 16 105
use FILL  FILL_707
timestamp 1680363874
transform 1 0 456 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_65
timestamp 1680363874
transform -1 0 504 0 -1 4170
box -8 -3 46 105
use FILL  FILL_708
timestamp 1680363874
transform 1 0 504 0 -1 4170
box -8 -3 16 105
use FILL  FILL_709
timestamp 1680363874
transform 1 0 512 0 -1 4170
box -8 -3 16 105
use FILL  FILL_710
timestamp 1680363874
transform 1 0 520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_711
timestamp 1680363874
transform 1 0 528 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_66
timestamp 1680363874
transform 1 0 536 0 -1 4170
box -8 -3 46 105
use FILL  FILL_712
timestamp 1680363874
transform 1 0 576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_713
timestamp 1680363874
transform 1 0 584 0 -1 4170
box -8 -3 16 105
use FILL  FILL_714
timestamp 1680363874
transform 1 0 592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_715
timestamp 1680363874
transform 1 0 600 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1215
timestamp 1680363874
transform 1 0 628 0 1 4075
box -3 -3 3 3
use OAI22X1  OAI22X1_67
timestamp 1680363874
transform 1 0 608 0 -1 4170
box -8 -3 46 105
use FILL  FILL_716
timestamp 1680363874
transform 1 0 648 0 -1 4170
box -8 -3 16 105
use FILL  FILL_717
timestamp 1680363874
transform 1 0 656 0 -1 4170
box -8 -3 16 105
use FILL  FILL_718
timestamp 1680363874
transform 1 0 664 0 -1 4170
box -8 -3 16 105
use FILL  FILL_719
timestamp 1680363874
transform 1 0 672 0 -1 4170
box -8 -3 16 105
use FILL  FILL_720
timestamp 1680363874
transform 1 0 680 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_69
timestamp 1680363874
transform 1 0 688 0 -1 4170
box -8 -3 46 105
use FILL  FILL_725
timestamp 1680363874
transform 1 0 728 0 -1 4170
box -8 -3 16 105
use FILL  FILL_726
timestamp 1680363874
transform 1 0 736 0 -1 4170
box -8 -3 16 105
use FILL  FILL_727
timestamp 1680363874
transform 1 0 744 0 -1 4170
box -8 -3 16 105
use FILL  FILL_728
timestamp 1680363874
transform 1 0 752 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1680363874
transform 1 0 760 0 -1 4170
box -8 -3 34 105
use FILL  FILL_731
timestamp 1680363874
transform 1 0 792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_732
timestamp 1680363874
transform 1 0 800 0 -1 4170
box -8 -3 16 105
use FILL  FILL_734
timestamp 1680363874
transform 1 0 808 0 -1 4170
box -8 -3 16 105
use FILL  FILL_737
timestamp 1680363874
transform 1 0 816 0 -1 4170
box -8 -3 16 105
use FILL  FILL_738
timestamp 1680363874
transform 1 0 824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_739
timestamp 1680363874
transform 1 0 832 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_80
timestamp 1680363874
transform -1 0 856 0 -1 4170
box -9 -3 26 105
use FILL  FILL_740
timestamp 1680363874
transform 1 0 856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_742
timestamp 1680363874
transform 1 0 864 0 -1 4170
box -8 -3 16 105
use FILL  FILL_744
timestamp 1680363874
transform 1 0 872 0 -1 4170
box -8 -3 16 105
use FILL  FILL_746
timestamp 1680363874
transform 1 0 880 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_14
timestamp 1680363874
transform 1 0 888 0 -1 4170
box -8 -3 34 105
use FILL  FILL_748
timestamp 1680363874
transform 1 0 920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_750
timestamp 1680363874
transform 1 0 928 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1216
timestamp 1680363874
transform 1 0 948 0 1 4075
box -3 -3 3 3
use FILL  FILL_752
timestamp 1680363874
transform 1 0 936 0 -1 4170
box -8 -3 16 105
use FILL  FILL_754
timestamp 1680363874
transform 1 0 944 0 -1 4170
box -8 -3 16 105
use FILL  FILL_756
timestamp 1680363874
transform 1 0 952 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_71
timestamp 1680363874
transform 1 0 960 0 -1 4170
box -8 -3 46 105
use FILL  FILL_758
timestamp 1680363874
transform 1 0 1000 0 -1 4170
box -8 -3 16 105
use FILL  FILL_760
timestamp 1680363874
transform 1 0 1008 0 -1 4170
box -8 -3 16 105
use FILL  FILL_762
timestamp 1680363874
transform 1 0 1016 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_73
timestamp 1680363874
transform 1 0 1024 0 -1 4170
box -8 -3 46 105
use FILL  FILL_764
timestamp 1680363874
transform 1 0 1064 0 -1 4170
box -8 -3 16 105
use FILL  FILL_765
timestamp 1680363874
transform 1 0 1072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_766
timestamp 1680363874
transform 1 0 1080 0 -1 4170
box -8 -3 16 105
use FILL  FILL_767
timestamp 1680363874
transform 1 0 1088 0 -1 4170
box -8 -3 16 105
use FILL  FILL_768
timestamp 1680363874
transform 1 0 1096 0 -1 4170
box -8 -3 16 105
use FILL  FILL_769
timestamp 1680363874
transform 1 0 1104 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_76
timestamp 1680363874
transform 1 0 1112 0 -1 4170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1680363874
transform 1 0 1152 0 -1 4170
box -8 -3 104 105
use FILL  FILL_777
timestamp 1680363874
transform 1 0 1248 0 -1 4170
box -8 -3 16 105
use FILL  FILL_778
timestamp 1680363874
transform 1 0 1256 0 -1 4170
box -8 -3 16 105
use FILL  FILL_779
timestamp 1680363874
transform 1 0 1264 0 -1 4170
box -8 -3 16 105
use FILL  FILL_780
timestamp 1680363874
transform 1 0 1272 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_81
timestamp 1680363874
transform -1 0 1296 0 -1 4170
box -9 -3 26 105
use FILL  FILL_781
timestamp 1680363874
transform 1 0 1296 0 -1 4170
box -8 -3 16 105
use FILL  FILL_783
timestamp 1680363874
transform 1 0 1304 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_78
timestamp 1680363874
transform 1 0 1312 0 -1 4170
box -8 -3 46 105
use FILL  FILL_805
timestamp 1680363874
transform 1 0 1352 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1680363874
transform -1 0 1456 0 -1 4170
box -8 -3 104 105
use FILL  FILL_806
timestamp 1680363874
transform 1 0 1456 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1680363874
transform 1 0 1464 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_86
timestamp 1680363874
transform -1 0 1576 0 -1 4170
box -9 -3 26 105
use M3_M2  M3_M2_1217
timestamp 1680363874
transform 1 0 1660 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_92
timestamp 1680363874
transform 1 0 1576 0 -1 4170
box -8 -3 104 105
use FILL  FILL_807
timestamp 1680363874
transform 1 0 1672 0 -1 4170
box -8 -3 16 105
use FILL  FILL_808
timestamp 1680363874
transform 1 0 1680 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1680363874
transform 1 0 1688 0 -1 4170
box -8 -3 104 105
use FILL  FILL_809
timestamp 1680363874
transform 1 0 1784 0 -1 4170
box -8 -3 16 105
use FILL  FILL_810
timestamp 1680363874
transform 1 0 1792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_811
timestamp 1680363874
transform 1 0 1800 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_79
timestamp 1680363874
transform -1 0 1848 0 -1 4170
box -8 -3 46 105
use FILL  FILL_812
timestamp 1680363874
transform 1 0 1848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_817
timestamp 1680363874
transform 1 0 1856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_818
timestamp 1680363874
transform 1 0 1864 0 -1 4170
box -8 -3 16 105
use FILL  FILL_819
timestamp 1680363874
transform 1 0 1872 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_80
timestamp 1680363874
transform -1 0 1920 0 -1 4170
box -8 -3 46 105
use FILL  FILL_820
timestamp 1680363874
transform 1 0 1920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_828
timestamp 1680363874
transform 1 0 1928 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1680363874
transform -1 0 2032 0 -1 4170
box -8 -3 104 105
use FILL  FILL_829
timestamp 1680363874
transform 1 0 2032 0 -1 4170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1680363874
transform 1 0 2040 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1680363874
transform 1 0 2048 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_89
timestamp 1680363874
transform 1 0 2144 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1680363874
transform 1 0 2160 0 -1 4170
box -8 -3 104 105
use FILL  FILL_844
timestamp 1680363874
transform 1 0 2256 0 -1 4170
box -8 -3 16 105
use FILL  FILL_845
timestamp 1680363874
transform 1 0 2264 0 -1 4170
box -8 -3 16 105
use FILL  FILL_846
timestamp 1680363874
transform 1 0 2272 0 -1 4170
box -8 -3 16 105
use FILL  FILL_851
timestamp 1680363874
transform 1 0 2280 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_82
timestamp 1680363874
transform -1 0 2328 0 -1 4170
box -8 -3 46 105
use FILL  FILL_852
timestamp 1680363874
transform 1 0 2328 0 -1 4170
box -8 -3 16 105
use FILL  FILL_853
timestamp 1680363874
transform 1 0 2336 0 -1 4170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1680363874
transform 1 0 2344 0 -1 4170
box -8 -3 16 105
use FILL  FILL_855
timestamp 1680363874
transform 1 0 2352 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_51
timestamp 1680363874
transform -1 0 2400 0 -1 4170
box -8 -3 46 105
use FILL  FILL_856
timestamp 1680363874
transform 1 0 2400 0 -1 4170
box -8 -3 16 105
use FILL  FILL_857
timestamp 1680363874
transform 1 0 2408 0 -1 4170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1680363874
transform 1 0 2416 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1680363874
transform 1 0 2424 0 -1 4170
box -8 -3 104 105
use FILL  FILL_871
timestamp 1680363874
transform 1 0 2520 0 -1 4170
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1680363874
transform -1 0 2560 0 -1 4170
box -8 -3 40 105
use FILL  FILL_872
timestamp 1680363874
transform 1 0 2560 0 -1 4170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1680363874
transform 1 0 2568 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_92
timestamp 1680363874
transform 1 0 2576 0 -1 4170
box -9 -3 26 105
use FILL  FILL_874
timestamp 1680363874
transform 1 0 2592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1680363874
transform 1 0 2600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_876
timestamp 1680363874
transform 1 0 2608 0 -1 4170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1680363874
transform 1 0 2616 0 -1 4170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1680363874
transform 1 0 2624 0 -1 4170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1680363874
transform 1 0 2632 0 -1 4170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1680363874
transform 1 0 2640 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1680363874
transform 1 0 2648 0 -1 4170
box -8 -3 104 105
use FILL  FILL_888
timestamp 1680363874
transform 1 0 2744 0 -1 4170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1680363874
transform 1 0 2752 0 -1 4170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1680363874
transform 1 0 2760 0 -1 4170
box -8 -3 16 105
use FILL  FILL_891
timestamp 1680363874
transform 1 0 2768 0 -1 4170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1680363874
transform 1 0 2776 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1680363874
transform 1 0 2784 0 -1 4170
box -8 -3 104 105
use FILL  FILL_899
timestamp 1680363874
transform 1 0 2880 0 -1 4170
box -8 -3 16 105
use FILL  FILL_900
timestamp 1680363874
transform 1 0 2888 0 -1 4170
box -8 -3 16 105
use FILL  FILL_901
timestamp 1680363874
transform 1 0 2896 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_83
timestamp 1680363874
transform -1 0 2944 0 -1 4170
box -8 -3 46 105
use FILL  FILL_902
timestamp 1680363874
transform 1 0 2944 0 -1 4170
box -8 -3 16 105
use FILL  FILL_903
timestamp 1680363874
transform 1 0 2952 0 -1 4170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1680363874
transform 1 0 2960 0 -1 4170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1680363874
transform 1 0 2968 0 -1 4170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1680363874
transform 1 0 2976 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_84
timestamp 1680363874
transform -1 0 3024 0 -1 4170
box -8 -3 46 105
use FILL  FILL_914
timestamp 1680363874
transform 1 0 3024 0 -1 4170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1680363874
transform 1 0 3032 0 -1 4170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1680363874
transform 1 0 3040 0 -1 4170
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1680363874
transform 1 0 3048 0 -1 4170
box -8 -3 40 105
use FILL  FILL_922
timestamp 1680363874
transform 1 0 3080 0 -1 4170
box -8 -3 16 105
use FILL  FILL_944
timestamp 1680363874
transform 1 0 3088 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1218
timestamp 1680363874
transform 1 0 3116 0 1 4075
box -3 -3 3 3
use AND2X2  AND2X2_3
timestamp 1680363874
transform 1 0 3096 0 -1 4170
box -8 -3 40 105
use FILL  FILL_945
timestamp 1680363874
transform 1 0 3128 0 -1 4170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1680363874
transform 1 0 3136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1680363874
transform 1 0 3144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1680363874
transform 1 0 3152 0 -1 4170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1680363874
transform 1 0 3160 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1219
timestamp 1680363874
transform 1 0 3244 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_104
timestamp 1680363874
transform -1 0 3264 0 -1 4170
box -8 -3 104 105
use FILL  FILL_950
timestamp 1680363874
transform 1 0 3264 0 -1 4170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1680363874
transform 1 0 3272 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_98
timestamp 1680363874
transform -1 0 3296 0 -1 4170
box -9 -3 26 105
use FILL  FILL_952
timestamp 1680363874
transform 1 0 3296 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_56
timestamp 1680363874
transform -1 0 3344 0 -1 4170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1680363874
transform 1 0 3344 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_99
timestamp 1680363874
transform -1 0 3456 0 -1 4170
box -9 -3 26 105
use FILL  FILL_953
timestamp 1680363874
transform 1 0 3456 0 -1 4170
box -8 -3 16 105
use FILL  FILL_965
timestamp 1680363874
transform 1 0 3464 0 -1 4170
box -8 -3 16 105
use FILL  FILL_966
timestamp 1680363874
transform 1 0 3472 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_58
timestamp 1680363874
transform -1 0 3520 0 -1 4170
box -8 -3 46 105
use FILL  FILL_967
timestamp 1680363874
transform 1 0 3520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1680363874
transform 1 0 3528 0 -1 4170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1680363874
transform 1 0 3536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1680363874
transform 1 0 3544 0 -1 4170
box -8 -3 16 105
use FILL  FILL_971
timestamp 1680363874
transform 1 0 3552 0 -1 4170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1680363874
transform 1 0 3560 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_59
timestamp 1680363874
transform -1 0 3608 0 -1 4170
box -8 -3 46 105
use FILL  FILL_973
timestamp 1680363874
transform 1 0 3608 0 -1 4170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1680363874
transform 1 0 3616 0 -1 4170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1680363874
transform 1 0 3624 0 -1 4170
box -8 -3 16 105
use FILL  FILL_976
timestamp 1680363874
transform 1 0 3632 0 -1 4170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1680363874
transform 1 0 3640 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1680363874
transform 1 0 3648 0 -1 4170
box -8 -3 104 105
use FILL  FILL_978
timestamp 1680363874
transform 1 0 3744 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1680363874
transform 1 0 3752 0 -1 4170
box -8 -3 104 105
use FILL  FILL_979
timestamp 1680363874
transform 1 0 3848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1680363874
transform 1 0 3856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1680363874
transform 1 0 3864 0 -1 4170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1680363874
transform 1 0 3872 0 -1 4170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1680363874
transform 1 0 3880 0 -1 4170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1680363874
transform 1 0 3888 0 -1 4170
box -8 -3 16 105
use FILL  FILL_989
timestamp 1680363874
transform 1 0 3896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1680363874
transform 1 0 3904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1680363874
transform 1 0 3912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_992
timestamp 1680363874
transform 1 0 3920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1680363874
transform 1 0 3928 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1680363874
transform 1 0 3936 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1680363874
transform 1 0 3944 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1220
timestamp 1680363874
transform 1 0 3980 0 1 4075
box -3 -3 3 3
use INVX2  INVX2_104
timestamp 1680363874
transform 1 0 3952 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1017
timestamp 1680363874
transform 1 0 3968 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1680363874
transform 1 0 3976 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_0
timestamp 1680363874
transform 1 0 3984 0 -1 4170
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1680363874
transform 1 0 4008 0 -1 4170
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1680363874
transform 1 0 4032 0 -1 4170
box -8 -3 104 105
use OAI22X1  OAI22X1_87
timestamp 1680363874
transform -1 0 4168 0 -1 4170
box -8 -3 46 105
use INVX2  INVX2_105
timestamp 1680363874
transform 1 0 4168 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1680363874
transform -1 0 4280 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1019
timestamp 1680363874
transform 1 0 4280 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1680363874
transform 1 0 4288 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1680363874
transform 1 0 4296 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1021
timestamp 1680363874
transform 1 0 4392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1680363874
transform 1 0 4400 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1680363874
transform 1 0 4408 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_63
timestamp 1680363874
transform 1 0 4416 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1027
timestamp 1680363874
transform 1 0 4456 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1680363874
transform 1 0 4464 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1680363874
transform 1 0 4472 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1680363874
transform 1 0 4480 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1680363874
transform 1 0 4488 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1680363874
transform 1 0 4496 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_89
timestamp 1680363874
transform 1 0 4504 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1039
timestamp 1680363874
transform 1 0 4544 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1680363874
transform 1 0 4552 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1680363874
transform 1 0 4560 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1680363874
transform 1 0 4568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1680363874
transform 1 0 4576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1680363874
transform 1 0 4584 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_66
timestamp 1680363874
transform -1 0 4632 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1047
timestamp 1680363874
transform 1 0 4632 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1680363874
transform 1 0 4640 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1680363874
transform 1 0 4648 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1680363874
transform 1 0 4656 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1680363874
transform 1 0 4664 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1680363874
transform 1 0 4672 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_106
timestamp 1680363874
transform 1 0 4680 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1680363874
transform 1 0 4696 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1060
timestamp 1680363874
transform 1 0 4792 0 -1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_13
timestamp 1680363874
transform 1 0 4851 0 1 4070
box -10 -3 10 3
use M2_M1  M2_M1_1430
timestamp 1680363874
transform 1 0 76 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1680363874
transform 1 0 132 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1680363874
transform 1 0 156 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1680363874
transform 1 0 172 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1331
timestamp 1680363874
transform 1 0 132 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1529
timestamp 1680363874
transform 1 0 188 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1680363874
transform 1 0 228 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1680363874
transform 1 0 212 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1432
timestamp 1680363874
transform 1 0 212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1680363874
transform 1 0 228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1680363874
transform 1 0 244 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1680363874
transform 1 0 220 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1680363874
transform 1 0 236 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1332
timestamp 1680363874
transform 1 0 220 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1680363874
transform 1 0 252 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1680363874
transform 1 0 276 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1241
timestamp 1680363874
transform 1 0 420 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1434
timestamp 1680363874
transform 1 0 348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1680363874
transform 1 0 380 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1680363874
transform 1 0 444 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1680363874
transform 1 0 300 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1303
timestamp 1680363874
transform 1 0 348 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1680363874
transform 1 0 372 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1680363874
transform 1 0 300 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1680363874
transform 1 0 292 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1680363874
transform 1 0 396 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1305
timestamp 1680363874
transform 1 0 444 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1680363874
transform 1 0 468 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1680363874
transform 1 0 396 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1680363874
transform 1 0 412 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1437
timestamp 1680363874
transform 1 0 492 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1254
timestamp 1680363874
transform 1 0 572 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1438
timestamp 1680363874
transform 1 0 548 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1279
timestamp 1680363874
transform 1 0 556 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1439
timestamp 1680363874
transform 1 0 564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1680363874
transform 1 0 540 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1680363874
transform 1 0 556 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1680363874
transform 1 0 572 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1680363874
transform 1 0 580 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1336
timestamp 1680363874
transform 1 0 540 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1680363874
transform 1 0 580 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1680363874
transform 1 0 572 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1680363874
transform 1 0 620 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1440
timestamp 1680363874
transform 1 0 620 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1680363874
transform 1 0 644 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1680363874
transform 1 0 636 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1307
timestamp 1680363874
transform 1 0 644 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1680363874
transform 1 0 660 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1442
timestamp 1680363874
transform 1 0 660 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1680363874
transform 1 0 652 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1338
timestamp 1680363874
transform 1 0 652 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1680363874
transform 1 0 636 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1443
timestamp 1680363874
transform 1 0 708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1680363874
transform 1 0 684 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1680363874
transform 1 0 700 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1308
timestamp 1680363874
transform 1 0 708 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1680363874
transform 1 0 748 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1444
timestamp 1680363874
transform 1 0 740 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1680363874
transform 1 0 724 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1680363874
transform 1 0 732 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1680363874
transform 1 0 780 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1680363874
transform 1 0 796 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1257
timestamp 1680363874
transform 1 0 804 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1680363874
transform 1 0 804 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1419
timestamp 1680363874
transform 1 0 836 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1680363874
transform 1 0 852 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1680363874
transform 1 0 860 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1371
timestamp 1680363874
transform 1 0 900 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1680363874
transform 1 0 932 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1446
timestamp 1680363874
transform 1 0 940 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1680363874
transform 1 0 932 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1258
timestamp 1680363874
transform 1 0 964 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1421
timestamp 1680363874
transform 1 0 972 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1680363874
transform 1 0 956 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1281
timestamp 1680363874
transform 1 0 964 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1545
timestamp 1680363874
transform 1 0 948 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1339
timestamp 1680363874
transform 1 0 940 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1680363874
transform 1 0 932 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1448
timestamp 1680363874
transform 1 0 980 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1309
timestamp 1680363874
transform 1 0 988 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1546
timestamp 1680363874
transform 1 0 1004 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1242
timestamp 1680363874
transform 1 0 1020 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1680363874
transform 1 0 1028 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1449
timestamp 1680363874
transform 1 0 1020 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1680363874
transform 1 0 1036 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1243
timestamp 1680363874
transform 1 0 1060 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1680363874
transform 1 0 1052 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1547
timestamp 1680363874
transform 1 0 1028 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1680363874
transform 1 0 1044 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1680363874
transform 1 0 1052 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1340
timestamp 1680363874
transform 1 0 1028 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1451
timestamp 1680363874
transform 1 0 1068 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1310
timestamp 1680363874
transform 1 0 1068 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1680363874
transform 1 0 1100 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1680363874
transform 1 0 1100 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1452
timestamp 1680363874
transform 1 0 1108 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1680363874
transform 1 0 1100 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1680363874
transform 1 0 1116 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1311
timestamp 1680363874
transform 1 0 1124 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1453
timestamp 1680363874
transform 1 0 1140 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1680363874
transform 1 0 1196 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1680363874
transform 1 0 1220 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1341
timestamp 1680363874
transform 1 0 1220 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1455
timestamp 1680363874
transform 1 0 1292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1680363874
transform 1 0 1268 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1312
timestamp 1680363874
transform 1 0 1316 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1680363874
transform 1 0 1268 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1456
timestamp 1680363874
transform 1 0 1356 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1680363874
transform 1 0 1372 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1680363874
transform 1 0 1388 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1261
timestamp 1680363874
transform 1 0 1420 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1458
timestamp 1680363874
transform 1 0 1404 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1680363874
transform 1 0 1420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1680363874
transform 1 0 1396 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1680363874
transform 1 0 1412 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1313
timestamp 1680363874
transform 1 0 1420 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1557
timestamp 1680363874
transform 1 0 1428 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1343
timestamp 1680363874
transform 1 0 1412 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1680363874
transform 1 0 1428 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1680363874
transform 1 0 1452 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1680363874
transform 1 0 1556 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1460
timestamp 1680363874
transform 1 0 1492 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1680363874
transform 1 0 1548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1680363874
transform 1 0 1556 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1680363874
transform 1 0 1468 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1344
timestamp 1680363874
transform 1 0 1492 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1559
timestamp 1680363874
transform 1 0 1564 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1263
timestamp 1680363874
transform 1 0 1620 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1680363874
transform 1 0 1612 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1463
timestamp 1680363874
transform 1 0 1620 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1680363874
transform 1 0 1636 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1680363874
transform 1 0 1612 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1314
timestamp 1680363874
transform 1 0 1620 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1561
timestamp 1680363874
transform 1 0 1636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1680363874
transform 1 0 1652 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1264
timestamp 1680363874
transform 1 0 1660 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1680363874
transform 1 0 1668 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1465
timestamp 1680363874
transform 1 0 1716 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1285
timestamp 1680363874
transform 1 0 1740 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1466
timestamp 1680363874
transform 1 0 1748 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1680363874
transform 1 0 1764 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1680363874
transform 1 0 1732 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1680363874
transform 1 0 1740 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1680363874
transform 1 0 1756 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1680363874
transform 1 0 1780 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1315
timestamp 1680363874
transform 1 0 1796 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1469
timestamp 1680363874
transform 1 0 1820 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1680363874
transform 1 0 1836 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1680363874
transform 1 0 1828 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1680363874
transform 1 0 1876 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1680363874
transform 1 0 1892 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1566
timestamp 1680363874
transform 1 0 1940 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1232
timestamp 1680363874
transform 1 0 1996 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1680363874
transform 1 0 2108 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1265
timestamp 1680363874
transform 1 0 2156 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1472
timestamp 1680363874
transform 1 0 2164 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1680363874
transform 1 0 2172 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1473
timestamp 1680363874
transform 1 0 2212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1680363874
transform 1 0 2196 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1680363874
transform 1 0 2204 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1680363874
transform 1 0 2220 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1345
timestamp 1680363874
transform 1 0 2220 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1474
timestamp 1680363874
transform 1 0 2236 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1221
timestamp 1680363874
transform 1 0 2276 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1680363874
transform 1 0 2300 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1680363874
transform 1 0 2316 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1680363874
transform 1 0 2292 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1475
timestamp 1680363874
transform 1 0 2292 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1287
timestamp 1680363874
transform 1 0 2340 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1423
timestamp 1680363874
transform 1 0 2356 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1680363874
transform 1 0 2348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1680363874
transform 1 0 2268 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1316
timestamp 1680363874
transform 1 0 2356 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1477
timestamp 1680363874
transform 1 0 2396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1680363874
transform 1 0 2412 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1680363874
transform 1 0 2404 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1346
timestamp 1680363874
transform 1 0 2404 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1680363874
transform 1 0 2444 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1680363874
transform 1 0 2444 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1223
timestamp 1680363874
transform 1 0 2468 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1479
timestamp 1680363874
transform 1 0 2460 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1680363874
transform 1 0 2460 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1268
timestamp 1680363874
transform 1 0 2516 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1680363874
transform 1 0 2532 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1480
timestamp 1680363874
transform 1 0 2500 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1680363874
transform 1 0 2516 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1680363874
transform 1 0 2532 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1680363874
transform 1 0 2540 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1317
timestamp 1680363874
transform 1 0 2500 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1680363874
transform 1 0 2508 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1680363874
transform 1 0 2524 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1347
timestamp 1680363874
transform 1 0 2524 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1680363874
transform 1 0 2540 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1680363874
transform 1 0 2596 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1680363874
transform 1 0 2572 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1484
timestamp 1680363874
transform 1 0 2580 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1680363874
transform 1 0 2572 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1680363874
transform 1 0 2588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1348
timestamp 1680363874
transform 1 0 2588 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1485
timestamp 1680363874
transform 1 0 2604 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1289
timestamp 1680363874
transform 1 0 2620 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1680363874
transform 1 0 2644 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1486
timestamp 1680363874
transform 1 0 2636 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1680363874
transform 1 0 2644 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1487
timestamp 1680363874
transform 1 0 2668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1680363874
transform 1 0 2716 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1680363874
transform 1 0 2732 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1349
timestamp 1680363874
transform 1 0 2636 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1680363874
transform 1 0 2732 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1488
timestamp 1680363874
transform 1 0 2748 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1245
timestamp 1680363874
transform 1 0 2764 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1489
timestamp 1680363874
transform 1 0 2820 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1680363874
transform 1 0 2772 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1319
timestamp 1680363874
transform 1 0 2820 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1680363874
transform 1 0 2844 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1490
timestamp 1680363874
transform 1 0 2868 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1680363874
transform 1 0 2876 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1351
timestamp 1680363874
transform 1 0 2868 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1491
timestamp 1680363874
transform 1 0 2884 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1680363874
transform 1 0 2892 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1352
timestamp 1680363874
transform 1 0 2892 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1492
timestamp 1680363874
transform 1 0 2940 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1353
timestamp 1680363874
transform 1 0 2948 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1680363874
transform 1 0 2980 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1271
timestamp 1680363874
transform 1 0 2988 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1493
timestamp 1680363874
transform 1 0 2996 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1291
timestamp 1680363874
transform 1 0 3020 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1680363874
transform 1 0 3044 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1425
timestamp 1680363874
transform 1 0 3052 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1680363874
transform 1 0 3020 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1680363874
transform 1 0 3028 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1273
timestamp 1680363874
transform 1 0 3100 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1494
timestamp 1680363874
transform 1 0 3116 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1680363874
transform 1 0 3100 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1680363874
transform 1 0 3132 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1292
timestamp 1680363874
transform 1 0 3132 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1495
timestamp 1680363874
transform 1 0 3140 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1321
timestamp 1680363874
transform 1 0 3140 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1586
timestamp 1680363874
transform 1 0 3148 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1322
timestamp 1680363874
transform 1 0 3156 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1680363874
transform 1 0 3172 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1680363874
transform 1 0 3180 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1680363874
transform 1 0 3196 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1496
timestamp 1680363874
transform 1 0 3188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1680363874
transform 1 0 3172 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1323
timestamp 1680363874
transform 1 0 3188 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1427
timestamp 1680363874
transform 1 0 3204 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1293
timestamp 1680363874
transform 1 0 3204 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1588
timestamp 1680363874
transform 1 0 3204 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1248
timestamp 1680363874
transform 1 0 3252 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1680363874
transform 1 0 3276 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1497
timestamp 1680363874
transform 1 0 3244 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1680363874
transform 1 0 3260 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1294
timestamp 1680363874
transform 1 0 3268 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1499
timestamp 1680363874
transform 1 0 3284 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1680363874
transform 1 0 3244 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1680363874
transform 1 0 3252 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1680363874
transform 1 0 3268 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1680363874
transform 1 0 3276 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1680363874
transform 1 0 3292 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1376
timestamp 1680363874
transform 1 0 3300 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1680363874
transform 1 0 3316 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1680363874
transform 1 0 3372 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1501
timestamp 1680363874
transform 1 0 3324 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1680363874
transform 1 0 3332 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1295
timestamp 1680363874
transform 1 0 3340 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1503
timestamp 1680363874
transform 1 0 3364 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1324
timestamp 1680363874
transform 1 0 3324 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1680363874
transform 1 0 3364 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1593
timestamp 1680363874
transform 1 0 3412 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1680363874
transform 1 0 3436 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1680363874
transform 1 0 3452 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1326
timestamp 1680363874
transform 1 0 3452 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1428
timestamp 1680363874
transform 1 0 3476 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1680363874
transform 1 0 3484 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1354
timestamp 1680363874
transform 1 0 3484 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1680363874
transform 1 0 3516 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1680363874
transform 1 0 3508 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1595
timestamp 1680363874
transform 1 0 3508 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1680363874
transform 1 0 3532 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1680363874
transform 1 0 3516 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1327
timestamp 1680363874
transform 1 0 3532 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1597
timestamp 1680363874
transform 1 0 3548 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1377
timestamp 1680363874
transform 1 0 3596 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1598
timestamp 1680363874
transform 1 0 3652 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1355
timestamp 1680363874
transform 1 0 3652 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1680363874
transform 1 0 3652 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1599
timestamp 1680363874
transform 1 0 3668 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1680363874
transform 1 0 3684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1680363874
transform 1 0 3700 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1680363874
transform 1 0 3716 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1680363874
transform 1 0 3708 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1680363874
transform 1 0 3724 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1356
timestamp 1680363874
transform 1 0 3716 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1680363874
transform 1 0 3708 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1602
timestamp 1680363874
transform 1 0 3740 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1680363874
transform 1 0 3780 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1357
timestamp 1680363874
transform 1 0 3780 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1510
timestamp 1680363874
transform 1 0 3796 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1680363874
transform 1 0 3836 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1380
timestamp 1680363874
transform 1 0 3828 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1680363874
transform 1 0 3852 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1680363874
transform 1 0 3956 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1511
timestamp 1680363874
transform 1 0 3916 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1680363874
transform 1 0 3948 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1680363874
transform 1 0 3956 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1680363874
transform 1 0 3868 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1359
timestamp 1680363874
transform 1 0 3868 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1680363874
transform 1 0 3972 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1514
timestamp 1680363874
transform 1 0 4044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1680363874
transform 1 0 4036 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1680363874
transform 1 0 4060 0 1 3995
box -2 -2 2 2
use M3_M2  M3_M2_1225
timestamp 1680363874
transform 1 0 4140 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1680363874
transform 1 0 4148 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1680363874
transform 1 0 4164 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1515
timestamp 1680363874
transform 1 0 4116 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1297
timestamp 1680363874
transform 1 0 4148 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1516
timestamp 1680363874
transform 1 0 4164 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1680363874
transform 1 0 4148 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1361
timestamp 1680363874
transform 1 0 4148 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1680363874
transform 1 0 4180 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1517
timestamp 1680363874
transform 1 0 4196 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1237
timestamp 1680363874
transform 1 0 4220 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1607
timestamp 1680363874
transform 1 0 4212 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1680363874
transform 1 0 4204 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1680363874
transform 1 0 4284 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1298
timestamp 1680363874
transform 1 0 4308 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1608
timestamp 1680363874
transform 1 0 4308 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1362
timestamp 1680363874
transform 1 0 4308 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1680363874
transform 1 0 4324 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1609
timestamp 1680363874
transform 1 0 4340 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1363
timestamp 1680363874
transform 1 0 4332 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1680363874
transform 1 0 4372 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1680363874
transform 1 0 4356 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1519
timestamp 1680363874
transform 1 0 4356 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1680363874
transform 1 0 4372 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1680363874
transform 1 0 4364 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1680363874
transform 1 0 4388 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1381
timestamp 1680363874
transform 1 0 4380 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1680363874
transform 1 0 4396 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1364
timestamp 1680363874
transform 1 0 4396 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1522
timestamp 1680363874
transform 1 0 4428 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1680363874
transform 1 0 4420 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1328
timestamp 1680363874
transform 1 0 4428 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1680363874
transform 1 0 4444 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1680363874
transform 1 0 4460 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1680363874
transform 1 0 4452 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1523
timestamp 1680363874
transform 1 0 4444 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1680363874
transform 1 0 4460 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1680363874
transform 1 0 4452 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1680363874
transform 1 0 4476 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1680363874
transform 1 0 4484 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1365
timestamp 1680363874
transform 1 0 4476 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1680363874
transform 1 0 4532 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1680363874
transform 1 0 4508 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1680363874
transform 1 0 4564 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1680363874
transform 1 0 4500 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1680363874
transform 1 0 4500 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1680363874
transform 1 0 4564 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1300
timestamp 1680363874
transform 1 0 4588 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1680363874
transform 1 0 4524 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1615
timestamp 1680363874
transform 1 0 4588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1278
timestamp 1680363874
transform 1 0 4604 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1526
timestamp 1680363874
transform 1 0 4604 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1680363874
transform 1 0 4612 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1301
timestamp 1680363874
transform 1 0 4708 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1680363874
transform 1 0 4740 0 1 4015
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_14
timestamp 1680363874
transform 1 0 48 0 1 3970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_117
timestamp 1680363874
transform -1 0 168 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_107
timestamp 1680363874
transform 1 0 168 0 1 3970
box -9 -3 26 105
use FILL  FILL_1061
timestamp 1680363874
transform 1 0 184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1680363874
transform 1 0 192 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_90
timestamp 1680363874
transform 1 0 200 0 1 3970
box -8 -3 46 105
use FILL  FILL_1063
timestamp 1680363874
transform 1 0 240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1680363874
transform 1 0 248 0 1 3970
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1680363874
transform 1 0 256 0 1 3970
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1680363874
transform 1 0 264 0 1 3970
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1680363874
transform 1 0 272 0 1 3970
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1680363874
transform 1 0 280 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1680363874
transform 1 0 288 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_1382
timestamp 1680363874
transform 1 0 460 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_120
timestamp 1680363874
transform 1 0 384 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_109
timestamp 1680363874
transform 1 0 480 0 1 3970
box -9 -3 26 105
use FILL  FILL_1069
timestamp 1680363874
transform 1 0 496 0 1 3970
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1680363874
transform 1 0 504 0 1 3970
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1680363874
transform 1 0 512 0 1 3970
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1680363874
transform 1 0 520 0 1 3970
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1680363874
transform 1 0 528 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_94
timestamp 1680363874
transform 1 0 536 0 1 3970
box -8 -3 46 105
use FILL  FILL_1089
timestamp 1680363874
transform 1 0 576 0 1 3970
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1680363874
transform 1 0 584 0 1 3970
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1680363874
transform 1 0 592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1680363874
transform 1 0 600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1680363874
transform 1 0 608 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_96
timestamp 1680363874
transform 1 0 616 0 1 3970
box -8 -3 46 105
use FILL  FILL_1098
timestamp 1680363874
transform 1 0 656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1680363874
transform 1 0 664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1680363874
transform 1 0 672 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_98
timestamp 1680363874
transform 1 0 680 0 1 3970
box -8 -3 46 105
use FILL  FILL_1105
timestamp 1680363874
transform 1 0 720 0 1 3970
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1680363874
transform 1 0 728 0 1 3970
box -8 -3 32 105
use FILL  FILL_1109
timestamp 1680363874
transform 1 0 752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1680363874
transform 1 0 760 0 1 3970
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1680363874
transform 1 0 768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1680363874
transform 1 0 776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1680363874
transform 1 0 784 0 1 3970
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1680363874
transform 1 0 792 0 1 3970
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1680363874
transform 1 0 800 0 1 3970
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1680363874
transform 1 0 808 0 1 3970
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1680363874
transform 1 0 816 0 1 3970
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1680363874
transform 1 0 824 0 1 3970
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1680363874
transform -1 0 856 0 1 3970
box -8 -3 32 105
use FILL  FILL_1127
timestamp 1680363874
transform 1 0 856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1680363874
transform 1 0 864 0 1 3970
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1680363874
transform 1 0 872 0 1 3970
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1680363874
transform 1 0 880 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_16
timestamp 1680363874
transform -1 0 920 0 1 3970
box -8 -3 34 105
use FILL  FILL_1135
timestamp 1680363874
transform 1 0 920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1680363874
transform 1 0 928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1680363874
transform 1 0 936 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1680363874
transform 1 0 944 0 1 3970
box -8 -3 34 105
use FILL  FILL_1138
timestamp 1680363874
transform 1 0 976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1680363874
transform 1 0 984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1680363874
transform 1 0 992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1680363874
transform 1 0 1000 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_99
timestamp 1680363874
transform 1 0 1008 0 1 3970
box -8 -3 46 105
use FILL  FILL_1142
timestamp 1680363874
transform 1 0 1048 0 1 3970
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1680363874
transform 1 0 1056 0 1 3970
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1680363874
transform 1 0 1064 0 1 3970
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1680363874
transform 1 0 1072 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_100
timestamp 1680363874
transform 1 0 1080 0 1 3970
box -8 -3 46 105
use FILL  FILL_1146
timestamp 1680363874
transform 1 0 1120 0 1 3970
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1680363874
transform 1 0 1128 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1383
timestamp 1680363874
transform 1 0 1204 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_122
timestamp 1680363874
transform -1 0 1232 0 1 3970
box -8 -3 104 105
use FILL  FILL_1148
timestamp 1680363874
transform 1 0 1232 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1384
timestamp 1680363874
transform 1 0 1252 0 1 3975
box -3 -3 3 3
use FILL  FILL_1168
timestamp 1680363874
transform 1 0 1240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1680363874
transform 1 0 1248 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1385
timestamp 1680363874
transform 1 0 1356 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_123
timestamp 1680363874
transform 1 0 1256 0 1 3970
box -8 -3 104 105
use FILL  FILL_1172
timestamp 1680363874
transform 1 0 1352 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1680363874
transform -1 0 1376 0 1 3970
box -9 -3 26 105
use FILL  FILL_1173
timestamp 1680363874
transform 1 0 1376 0 1 3970
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1680363874
transform 1 0 1384 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_105
timestamp 1680363874
transform -1 0 1432 0 1 3970
box -8 -3 46 105
use FILL  FILL_1175
timestamp 1680363874
transform 1 0 1432 0 1 3970
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1680363874
transform 1 0 1440 0 1 3970
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1680363874
transform 1 0 1448 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1680363874
transform 1 0 1456 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_113
timestamp 1680363874
transform -1 0 1568 0 1 3970
box -9 -3 26 105
use FILL  FILL_1178
timestamp 1680363874
transform 1 0 1568 0 1 3970
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1680363874
transform 1 0 1576 0 1 3970
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1680363874
transform 1 0 1584 0 1 3970
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1680363874
transform 1 0 1592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1680363874
transform 1 0 1600 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_19
timestamp 1680363874
transform 1 0 1608 0 1 3970
box -8 -3 34 105
use FILL  FILL_1196
timestamp 1680363874
transform 1 0 1640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1680363874
transform 1 0 1648 0 1 3970
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1680363874
transform 1 0 1656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1680363874
transform 1 0 1664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1680363874
transform 1 0 1672 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_116
timestamp 1680363874
transform -1 0 1696 0 1 3970
box -9 -3 26 105
use FILL  FILL_1206
timestamp 1680363874
transform 1 0 1696 0 1 3970
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1680363874
transform 1 0 1704 0 1 3970
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1680363874
transform 1 0 1712 0 1 3970
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1680363874
transform 1 0 1720 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_67
timestamp 1680363874
transform -1 0 1768 0 1 3970
box -8 -3 46 105
use FILL  FILL_1212
timestamp 1680363874
transform 1 0 1768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1680363874
transform 1 0 1776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1680363874
transform 1 0 1784 0 1 3970
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1680363874
transform 1 0 1792 0 1 3970
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1680363874
transform 1 0 1800 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_109
timestamp 1680363874
transform -1 0 1848 0 1 3970
box -8 -3 46 105
use FILL  FILL_1222
timestamp 1680363874
transform 1 0 1848 0 1 3970
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1680363874
transform 1 0 1856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1680363874
transform 1 0 1864 0 1 3970
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1680363874
transform 1 0 1872 0 1 3970
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1680363874
transform 1 0 1880 0 1 3970
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1680363874
transform 1 0 1888 0 1 3970
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1680363874
transform 1 0 1896 0 1 3970
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1680363874
transform 1 0 1904 0 1 3970
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1680363874
transform 1 0 1912 0 1 3970
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1680363874
transform 1 0 1920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1680363874
transform 1 0 1928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1680363874
transform 1 0 1936 0 1 3970
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1680363874
transform 1 0 1944 0 1 3970
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1680363874
transform 1 0 1952 0 1 3970
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1680363874
transform 1 0 1960 0 1 3970
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1680363874
transform 1 0 1968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1680363874
transform 1 0 1976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1680363874
transform 1 0 1984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1680363874
transform 1 0 1992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1680363874
transform 1 0 2000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1680363874
transform 1 0 2008 0 1 3970
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1680363874
transform 1 0 2016 0 1 3970
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1680363874
transform 1 0 2024 0 1 3970
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1680363874
transform 1 0 2032 0 1 3970
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1680363874
transform 1 0 2040 0 1 3970
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1680363874
transform 1 0 2048 0 1 3970
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1680363874
transform 1 0 2056 0 1 3970
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1680363874
transform 1 0 2064 0 1 3970
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1680363874
transform 1 0 2072 0 1 3970
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1680363874
transform 1 0 2080 0 1 3970
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1680363874
transform 1 0 2088 0 1 3970
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1680363874
transform 1 0 2096 0 1 3970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1680363874
transform 1 0 2104 0 1 3970
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1680363874
transform 1 0 2112 0 1 3970
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1680363874
transform 1 0 2120 0 1 3970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1680363874
transform 1 0 2128 0 1 3970
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1680363874
transform 1 0 2136 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_122
timestamp 1680363874
transform -1 0 2160 0 1 3970
box -9 -3 26 105
use FILL  FILL_1280
timestamp 1680363874
transform 1 0 2160 0 1 3970
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1680363874
transform 1 0 2168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1680363874
transform 1 0 2176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1680363874
transform 1 0 2184 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_72
timestamp 1680363874
transform -1 0 2232 0 1 3970
box -8 -3 46 105
use FILL  FILL_1290
timestamp 1680363874
transform 1 0 2232 0 1 3970
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1680363874
transform 1 0 2240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1680363874
transform 1 0 2248 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1386
timestamp 1680363874
transform 1 0 2276 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_126
timestamp 1680363874
transform 1 0 2256 0 1 3970
box -8 -3 104 105
use FILL  FILL_1302
timestamp 1680363874
transform 1 0 2352 0 1 3970
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1680363874
transform 1 0 2360 0 1 3970
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1680363874
transform 1 0 2368 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1387
timestamp 1680363874
transform 1 0 2396 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_73
timestamp 1680363874
transform -1 0 2416 0 1 3970
box -8 -3 46 105
use FILL  FILL_1305
timestamp 1680363874
transform 1 0 2416 0 1 3970
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1680363874
transform 1 0 2424 0 1 3970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1680363874
transform 1 0 2432 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_123
timestamp 1680363874
transform 1 0 2440 0 1 3970
box -9 -3 26 105
use FILL  FILL_1308
timestamp 1680363874
transform 1 0 2456 0 1 3970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1680363874
transform 1 0 2464 0 1 3970
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1680363874
transform 1 0 2472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1680363874
transform 1 0 2480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1680363874
transform 1 0 2488 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1388
timestamp 1680363874
transform 1 0 2524 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_76
timestamp 1680363874
transform -1 0 2536 0 1 3970
box -8 -3 46 105
use FILL  FILL_1327
timestamp 1680363874
transform 1 0 2536 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1389
timestamp 1680363874
transform 1 0 2556 0 1 3975
box -3 -3 3 3
use FILL  FILL_1328
timestamp 1680363874
transform 1 0 2544 0 1 3970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1680363874
transform 1 0 2552 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_77
timestamp 1680363874
transform -1 0 2600 0 1 3970
box -8 -3 46 105
use FILL  FILL_1330
timestamp 1680363874
transform 1 0 2600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1680363874
transform 1 0 2608 0 1 3970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1680363874
transform 1 0 2616 0 1 3970
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1680363874
transform 1 0 2624 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1390
timestamp 1680363874
transform 1 0 2716 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_127
timestamp 1680363874
transform -1 0 2728 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_126
timestamp 1680363874
transform 1 0 2728 0 1 3970
box -9 -3 26 105
use FILL  FILL_1334
timestamp 1680363874
transform 1 0 2744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1680363874
transform 1 0 2752 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1391
timestamp 1680363874
transform 1 0 2772 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_128
timestamp 1680363874
transform 1 0 2760 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_1392
timestamp 1680363874
transform 1 0 2884 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_127
timestamp 1680363874
transform 1 0 2856 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1680363874
transform 1 0 2872 0 1 3970
box -9 -3 26 105
use FILL  FILL_1336
timestamp 1680363874
transform 1 0 2888 0 1 3970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1680363874
transform 1 0 2896 0 1 3970
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1680363874
transform 1 0 2904 0 1 3970
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1680363874
transform 1 0 2912 0 1 3970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1680363874
transform 1 0 2920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1680363874
transform 1 0 2928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1680363874
transform 1 0 2936 0 1 3970
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1680363874
transform 1 0 2944 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_21
timestamp 1680363874
transform 1 0 2952 0 1 3970
box -8 -3 34 105
use FILL  FILL_1366
timestamp 1680363874
transform 1 0 2984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1680363874
transform 1 0 2992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1680363874
transform 1 0 3000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1680363874
transform 1 0 3008 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1393
timestamp 1680363874
transform 1 0 3028 0 1 3975
box -3 -3 3 3
use FILL  FILL_1370
timestamp 1680363874
transform 1 0 3016 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1680363874
transform 1 0 3024 0 1 3970
box -8 -3 34 105
use FILL  FILL_1376
timestamp 1680363874
transform 1 0 3056 0 1 3970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1680363874
transform 1 0 3064 0 1 3970
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1680363874
transform 1 0 3072 0 1 3970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1680363874
transform 1 0 3080 0 1 3970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1680363874
transform 1 0 3088 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1394
timestamp 1680363874
transform 1 0 3108 0 1 3975
box -3 -3 3 3
use OAI21X1  OAI21X1_24
timestamp 1680363874
transform -1 0 3128 0 1 3970
box -8 -3 34 105
use FILL  FILL_1381
timestamp 1680363874
transform 1 0 3128 0 1 3970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1680363874
transform 1 0 3136 0 1 3970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1680363874
transform 1 0 3144 0 1 3970
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1680363874
transform 1 0 3152 0 1 3970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1680363874
transform 1 0 3160 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1680363874
transform -1 0 3200 0 1 3970
box -8 -3 34 105
use FILL  FILL_1386
timestamp 1680363874
transform 1 0 3200 0 1 3970
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1680363874
transform 1 0 3208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1680363874
transform 1 0 3216 0 1 3970
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1680363874
transform 1 0 3224 0 1 3970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1680363874
transform 1 0 3232 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_78
timestamp 1680363874
transform 1 0 3240 0 1 3970
box -8 -3 46 105
use FILL  FILL_1401
timestamp 1680363874
transform 1 0 3280 0 1 3970
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1680363874
transform 1 0 3288 0 1 3970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1680363874
transform 1 0 3296 0 1 3970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1680363874
transform 1 0 3304 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_131
timestamp 1680363874
transform 1 0 3312 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1680363874
transform -1 0 3424 0 1 3970
box -8 -3 104 105
use FILL  FILL_1405
timestamp 1680363874
transform 1 0 3424 0 1 3970
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1680363874
transform 1 0 3432 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1395
timestamp 1680363874
transform 1 0 3476 0 1 3975
box -3 -3 3 3
use OAI21X1  OAI21X1_27
timestamp 1680363874
transform 1 0 3440 0 1 3970
box -8 -3 34 105
use FILL  FILL_1407
timestamp 1680363874
transform 1 0 3472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1680363874
transform 1 0 3480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1680363874
transform 1 0 3488 0 1 3970
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1680363874
transform 1 0 3496 0 1 3970
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1680363874
transform 1 0 3504 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_28
timestamp 1680363874
transform -1 0 3544 0 1 3970
box -8 -3 34 105
use FILL  FILL_1412
timestamp 1680363874
transform 1 0 3544 0 1 3970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1680363874
transform 1 0 3552 0 1 3970
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1680363874
transform 1 0 3560 0 1 3970
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1680363874
transform 1 0 3568 0 1 3970
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1680363874
transform 1 0 3576 0 1 3970
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1680363874
transform 1 0 3584 0 1 3970
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1680363874
transform 1 0 3592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1680363874
transform 1 0 3600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1680363874
transform 1 0 3608 0 1 3970
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1680363874
transform 1 0 3616 0 1 3970
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1680363874
transform 1 0 3624 0 1 3970
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1680363874
transform 1 0 3632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1680363874
transform 1 0 3640 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_135
timestamp 1680363874
transform 1 0 3648 0 1 3970
box -9 -3 26 105
use FILL  FILL_1445
timestamp 1680363874
transform 1 0 3664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1680363874
transform 1 0 3672 0 1 3970
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1680363874
transform 1 0 3680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1680363874
transform 1 0 3688 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_82
timestamp 1680363874
transform 1 0 3696 0 1 3970
box -8 -3 46 105
use FILL  FILL_1454
timestamp 1680363874
transform 1 0 3736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1680363874
transform 1 0 3744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1680363874
transform 1 0 3752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1680363874
transform 1 0 3760 0 1 3970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1680363874
transform 1 0 3768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1680363874
transform 1 0 3776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1680363874
transform 1 0 3784 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_136
timestamp 1680363874
transform -1 0 3808 0 1 3970
box -9 -3 26 105
use FILL  FILL_1467
timestamp 1680363874
transform 1 0 3808 0 1 3970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1680363874
transform 1 0 3816 0 1 3970
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1680363874
transform 1 0 3824 0 1 3970
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1680363874
transform 1 0 3832 0 1 3970
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1680363874
transform 1 0 3840 0 1 3970
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1680363874
transform 1 0 3848 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1680363874
transform 1 0 3856 0 1 3970
box -8 -3 104 105
use FILL  FILL_1477
timestamp 1680363874
transform 1 0 3952 0 1 3970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1680363874
transform 1 0 3960 0 1 3970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1680363874
transform 1 0 3968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1680363874
transform 1 0 3976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1680363874
transform 1 0 3984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1680363874
transform 1 0 3992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1680363874
transform 1 0 4000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1680363874
transform 1 0 4008 0 1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1680363874
transform -1 0 4040 0 1 3970
box -8 -3 32 105
use FILL  FILL_1496
timestamp 1680363874
transform 1 0 4040 0 1 3970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1680363874
transform 1 0 4048 0 1 3970
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1680363874
transform 1 0 4056 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1680363874
transform -1 0 4160 0 1 3970
box -8 -3 104 105
use NOR2X1  NOR2X1_2
timestamp 1680363874
transform -1 0 4184 0 1 3970
box -8 -3 32 105
use FILL  FILL_1503
timestamp 1680363874
transform 1 0 4184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1680363874
transform 1 0 4192 0 1 3970
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1680363874
transform 1 0 4200 0 1 3970
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1680363874
transform 1 0 4208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1680363874
transform 1 0 4216 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1396
timestamp 1680363874
transform 1 0 4300 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_136
timestamp 1680363874
transform -1 0 4320 0 1 3970
box -8 -3 104 105
use FILL  FILL_1519
timestamp 1680363874
transform 1 0 4320 0 1 3970
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1680363874
transform 1 0 4328 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1397
timestamp 1680363874
transform 1 0 4348 0 1 3975
box -3 -3 3 3
use FILL  FILL_1530
timestamp 1680363874
transform 1 0 4336 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_113
timestamp 1680363874
transform 1 0 4344 0 1 3970
box -8 -3 46 105
use FILL  FILL_1531
timestamp 1680363874
transform 1 0 4384 0 1 3970
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1680363874
transform 1 0 4392 0 1 3970
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1680363874
transform 1 0 4400 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_139
timestamp 1680363874
transform -1 0 4424 0 1 3970
box -9 -3 26 105
use NOR2X1  NOR2X1_3
timestamp 1680363874
transform -1 0 4448 0 1 3970
box -8 -3 32 105
use FILL  FILL_1534
timestamp 1680363874
transform 1 0 4448 0 1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1680363874
transform -1 0 4480 0 1 3970
box -8 -3 32 105
use FILL  FILL_1535
timestamp 1680363874
transform 1 0 4480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1680363874
transform 1 0 4488 0 1 3970
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1680363874
transform 1 0 4496 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1680363874
transform -1 0 4600 0 1 3970
box -8 -3 104 105
use FILL  FILL_1538
timestamp 1680363874
transform 1 0 4600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1680363874
transform 1 0 4608 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1680363874
transform 1 0 4616 0 1 3970
box -9 -3 26 105
use FILL  FILL_1540
timestamp 1680363874
transform 1 0 4632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1680363874
transform 1 0 4640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1680363874
transform 1 0 4648 0 1 3970
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1680363874
transform 1 0 4656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1680363874
transform 1 0 4664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1680363874
transform 1 0 4672 0 1 3970
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1680363874
transform 1 0 4680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1680363874
transform 1 0 4688 0 1 3970
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1680363874
transform 1 0 4696 0 1 3970
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1680363874
transform 1 0 4704 0 1 3970
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1680363874
transform 1 0 4712 0 1 3970
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1680363874
transform 1 0 4720 0 1 3970
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1680363874
transform 1 0 4728 0 1 3970
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1680363874
transform 1 0 4736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1680363874
transform 1 0 4744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1680363874
transform 1 0 4752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1680363874
transform 1 0 4760 0 1 3970
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1680363874
transform 1 0 4768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1680363874
transform 1 0 4776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1680363874
transform 1 0 4784 0 1 3970
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1680363874
transform 1 0 4792 0 1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_15
timestamp 1680363874
transform 1 0 4827 0 1 3970
box -10 -3 10 3
use M3_M2  M3_M2_1398
timestamp 1680363874
transform 1 0 76 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1680363874
transform 1 0 172 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1680363874
transform 1 0 188 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1680363874
transform 1 0 172 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1680363874
transform 1 0 196 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1680363874
transform 1 0 268 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1680363874
transform 1 0 84 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1680363874
transform 1 0 84 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1680363874
transform 1 0 132 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1544
timestamp 1680363874
transform 1 0 132 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1680363874
transform 1 0 196 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1680363874
transform 1 0 244 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1680363874
transform 1 0 300 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1624
timestamp 1680363874
transform 1 0 196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1680363874
transform 1 0 284 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1680363874
transform 1 0 300 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1680363874
transform 1 0 180 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1680363874
transform 1 0 244 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1680363874
transform 1 0 276 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1680363874
transform 1 0 292 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1680363874
transform 1 0 308 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1545
timestamp 1680363874
transform 1 0 220 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1680363874
transform 1 0 180 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1680363874
transform 1 0 356 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1680363874
transform 1 0 388 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1627
timestamp 1680363874
transform 1 0 348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1680363874
transform 1 0 356 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1680363874
transform 1 0 364 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1680363874
transform 1 0 404 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1629
timestamp 1680363874
transform 1 0 372 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1680363874
transform 1 0 388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1680363874
transform 1 0 396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1680363874
transform 1 0 364 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1508
timestamp 1680363874
transform 1 0 372 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1744
timestamp 1680363874
transform 1 0 380 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1546
timestamp 1680363874
transform 1 0 364 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1680363874
transform 1 0 380 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1745
timestamp 1680363874
transform 1 0 396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1547
timestamp 1680363874
transform 1 0 396 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1680363874
transform 1 0 420 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1680363874
transform 1 0 420 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1680363874
transform 1 0 484 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1633
timestamp 1680363874
transform 1 0 452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1680363874
transform 1 0 468 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1680363874
transform 1 0 484 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1680363874
transform 1 0 460 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1630
timestamp 1680363874
transform 1 0 452 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1747
timestamp 1680363874
transform 1 0 492 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1680363874
transform 1 0 508 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1680363874
transform 1 0 524 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1548
timestamp 1680363874
transform 1 0 524 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1680363874
transform 1 0 556 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1638
timestamp 1680363874
transform 1 0 556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1680363874
transform 1 0 572 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1680363874
transform 1 0 580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1680363874
transform 1 0 548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1680363874
transform 1 0 564 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1549
timestamp 1680363874
transform 1 0 580 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1680363874
transform 1 0 572 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1680363874
transform 1 0 564 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1641
timestamp 1680363874
transform 1 0 628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1680363874
transform 1 0 644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1680363874
transform 1 0 620 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1680363874
transform 1 0 628 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1751
timestamp 1680363874
transform 1 0 636 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1588
timestamp 1680363874
transform 1 0 644 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1752
timestamp 1680363874
transform 1 0 668 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1680363874
transform 1 0 692 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1680363874
transform 1 0 732 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1477
timestamp 1680363874
transform 1 0 756 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1854
timestamp 1680363874
transform 1 0 764 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1680363874
transform 1 0 772 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1478
timestamp 1680363874
transform 1 0 788 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1645
timestamp 1680363874
transform 1 0 804 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1510
timestamp 1680363874
transform 1 0 788 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1856
timestamp 1680363874
transform 1 0 812 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1680363874
transform 1 0 836 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1680363874
transform 1 0 836 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1857
timestamp 1680363874
transform 1 0 860 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1680363874
transform 1 0 876 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1511
timestamp 1680363874
transform 1 0 916 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1680363874
transform 1 0 940 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1646
timestamp 1680363874
transform 1 0 940 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1512
timestamp 1680363874
transform 1 0 940 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1680363874
transform 1 0 980 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1680363874
transform 1 0 972 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1647
timestamp 1680363874
transform 1 0 980 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1680363874
transform 1 0 996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1680363874
transform 1 0 972 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1680363874
transform 1 0 988 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1680363874
transform 1 0 1004 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1551
timestamp 1680363874
transform 1 0 996 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1680363874
transform 1 0 1004 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1680363874
transform 1 0 1036 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1680363874
transform 1 0 1068 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1680363874
transform 1 0 1084 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1649
timestamp 1680363874
transform 1 0 1044 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1680363874
transform 1 0 1052 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1680363874
transform 1 0 1068 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1480
timestamp 1680363874
transform 1 0 1076 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1652
timestamp 1680363874
transform 1 0 1084 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1680363874
transform 1 0 1092 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1513
timestamp 1680363874
transform 1 0 1052 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1758
timestamp 1680363874
transform 1 0 1060 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1680363874
transform 1 0 1076 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1552
timestamp 1680363874
transform 1 0 1044 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1680363874
transform 1 0 1052 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1680363874
transform 1 0 1092 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1680363874
transform 1 0 1108 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1680363874
transform 1 0 1140 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1680363874
transform 1 0 1164 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1680363874
transform 1 0 1156 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1680363874
transform 1 0 1132 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1654
timestamp 1680363874
transform 1 0 1140 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1680363874
transform 1 0 1156 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1680363874
transform 1 0 1124 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1680363874
transform 1 0 1148 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1592
timestamp 1680363874
transform 1 0 1148 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1762
timestamp 1680363874
transform 1 0 1164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1680363874
transform 1 0 1172 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1632
timestamp 1680363874
transform 1 0 1172 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1680363874
transform 1 0 1228 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1680363874
transform 1 0 1220 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1657
timestamp 1680363874
transform 1 0 1196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1680363874
transform 1 0 1212 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1680363874
transform 1 0 1204 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1680363874
transform 1 0 1220 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1593
timestamp 1680363874
transform 1 0 1212 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1659
timestamp 1680363874
transform 1 0 1228 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1680363874
transform 1 0 1236 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1633
timestamp 1680363874
transform 1 0 1236 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1661
timestamp 1680363874
transform 1 0 1292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1680363874
transform 1 0 1308 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1680363874
transform 1 0 1284 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1515
timestamp 1680363874
transform 1 0 1292 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1766
timestamp 1680363874
transform 1 0 1300 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1594
timestamp 1680363874
transform 1 0 1308 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1680363874
transform 1 0 1300 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1680363874
transform 1 0 1364 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1663
timestamp 1680363874
transform 1 0 1348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1680363874
transform 1 0 1364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1680363874
transform 1 0 1380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1680363874
transform 1 0 1356 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1680363874
transform 1 0 1372 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1553
timestamp 1680363874
transform 1 0 1372 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1680363874
transform 1 0 1348 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1680363874
transform 1 0 1396 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1680363874
transform 1 0 1388 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1769
timestamp 1680363874
transform 1 0 1396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1445
timestamp 1680363874
transform 1 0 1476 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1666
timestamp 1680363874
transform 1 0 1420 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1680363874
transform 1 0 1436 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1680363874
transform 1 0 1452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1680363874
transform 1 0 1428 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1680363874
transform 1 0 1476 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1596
timestamp 1680363874
transform 1 0 1436 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1680363874
transform 1 0 1428 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1772
timestamp 1680363874
transform 1 0 1556 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1680363874
transform 1 0 1564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1680363874
transform 1 0 1572 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1483
timestamp 1680363874
transform 1 0 1580 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1774
timestamp 1680363874
transform 1 0 1580 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1554
timestamp 1680363874
transform 1 0 1564 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1622
timestamp 1680363874
transform 1 0 1620 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1680363874
transform 1 0 1620 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1680363874
transform 1 0 1628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1680363874
transform 1 0 1636 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1597
timestamp 1680363874
transform 1 0 1636 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1672
timestamp 1680363874
transform 1 0 1676 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1555
timestamp 1680363874
transform 1 0 1676 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1680363874
transform 1 0 1708 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1680363874
transform 1 0 1700 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1673
timestamp 1680363874
transform 1 0 1692 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1598
timestamp 1680363874
transform 1 0 1692 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1776
timestamp 1680363874
transform 1 0 1700 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1484
timestamp 1680363874
transform 1 0 1716 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1680363874
transform 1 0 1748 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1777
timestamp 1680363874
transform 1 0 1716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1680363874
transform 1 0 1732 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1556
timestamp 1680363874
transform 1 0 1732 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1674
timestamp 1680363874
transform 1 0 1756 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1680363874
transform 1 0 1756 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1779
timestamp 1680363874
transform 1 0 1772 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1634
timestamp 1680363874
transform 1 0 1764 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1680363874
transform 1 0 1804 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1780
timestamp 1680363874
transform 1 0 1796 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1423
timestamp 1680363874
transform 1 0 1828 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1675
timestamp 1680363874
transform 1 0 1820 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1680363874
transform 1 0 1828 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1486
timestamp 1680363874
transform 1 0 1852 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1677
timestamp 1680363874
transform 1 0 1860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1680363874
transform 1 0 1820 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1518
timestamp 1680363874
transform 1 0 1828 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1782
timestamp 1680363874
transform 1 0 1836 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1519
timestamp 1680363874
transform 1 0 1844 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1783
timestamp 1680363874
transform 1 0 1852 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1557
timestamp 1680363874
transform 1 0 1820 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1680363874
transform 1 0 1876 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1784
timestamp 1680363874
transform 1 0 1900 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1680363874
transform 1 0 1932 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1680363874
transform 1 0 1964 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1678
timestamp 1680363874
transform 1 0 1940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1680363874
transform 1 0 1948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1680363874
transform 1 0 1964 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1680363874
transform 1 0 1932 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1680363874
transform 1 0 1956 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1520
timestamp 1680363874
transform 1 0 1964 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1787
timestamp 1680363874
transform 1 0 1996 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1680363874
transform 1 0 2004 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1488
timestamp 1680363874
transform 1 0 2028 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1789
timestamp 1680363874
transform 1 0 2028 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1449
timestamp 1680363874
transform 1 0 2076 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1681
timestamp 1680363874
transform 1 0 2044 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1680363874
transform 1 0 2052 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1680363874
transform 1 0 2076 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1521
timestamp 1680363874
transform 1 0 2044 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1680363874
transform 1 0 2036 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1680363874
transform 1 0 2060 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1790
timestamp 1680363874
transform 1 0 2068 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1560
timestamp 1680363874
transform 1 0 2060 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1680363874
transform 1 0 2100 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1680363874
transform 1 0 2108 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1791
timestamp 1680363874
transform 1 0 2100 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1680363874
transform 1 0 2108 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1490
timestamp 1680363874
transform 1 0 2164 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1680363874
transform 1 0 2188 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1680363874
transform 1 0 2204 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1680363874
transform 1 0 2204 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1680363874
transform 1 0 2220 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1680363874
transform 1 0 2212 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1621
timestamp 1680363874
transform 1 0 2252 0 1 3955
box -2 -2 2 2
use M3_M2  M3_M2_1451
timestamp 1680363874
transform 1 0 2252 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1863
timestamp 1680363874
transform 1 0 2252 0 1 3905
box -2 -2 2 2
use M3_M2  M3_M2_1452
timestamp 1680363874
transform 1 0 2268 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1684
timestamp 1680363874
transform 1 0 2276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1680363874
transform 1 0 2292 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1405
timestamp 1680363874
transform 1 0 2308 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1685
timestamp 1680363874
transform 1 0 2308 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1523
timestamp 1680363874
transform 1 0 2308 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1794
timestamp 1680363874
transform 1 0 2316 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1680363874
transform 1 0 2348 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1686
timestamp 1680363874
transform 1 0 2340 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1425
timestamp 1680363874
transform 1 0 2380 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1795
timestamp 1680363874
transform 1 0 2348 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1524
timestamp 1680363874
transform 1 0 2356 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1796
timestamp 1680363874
transform 1 0 2364 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1562
timestamp 1680363874
transform 1 0 2348 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1680363874
transform 1 0 2396 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1687
timestamp 1680363874
transform 1 0 2404 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1680363874
transform 1 0 2396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1525
timestamp 1680363874
transform 1 0 2404 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1680363874
transform 1 0 2436 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1680363874
transform 1 0 2420 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1688
timestamp 1680363874
transform 1 0 2428 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1680363874
transform 1 0 2444 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1680363874
transform 1 0 2452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1680363874
transform 1 0 2412 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1563
timestamp 1680363874
transform 1 0 2412 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1799
timestamp 1680363874
transform 1 0 2436 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1526
timestamp 1680363874
transform 1 0 2444 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1680363874
transform 1 0 2428 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1680363874
transform 1 0 2468 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1800
timestamp 1680363874
transform 1 0 2468 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1680363874
transform 1 0 2492 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1599
timestamp 1680363874
transform 1 0 2484 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1680363874
transform 1 0 2516 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1680363874
transform 1 0 2516 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1680363874
transform 1 0 2532 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1680363874
transform 1 0 2524 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1680363874
transform 1 0 2564 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1691
timestamp 1680363874
transform 1 0 2548 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1528
timestamp 1680363874
transform 1 0 2548 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1802
timestamp 1680363874
transform 1 0 2572 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1680363874
transform 1 0 2628 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1565
timestamp 1680363874
transform 1 0 2548 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1680363874
transform 1 0 2612 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1680363874
transform 1 0 2660 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1680363874
transform 1 0 2684 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1680363874
transform 1 0 2684 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1680363874
transform 1 0 2716 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1680363874
transform 1 0 2748 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1692
timestamp 1680363874
transform 1 0 2684 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1680363874
transform 1 0 2732 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1566
timestamp 1680363874
transform 1 0 2732 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1805
timestamp 1680363874
transform 1 0 2788 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1567
timestamp 1680363874
transform 1 0 2780 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1680363874
transform 1 0 2788 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1806
timestamp 1680363874
transform 1 0 2804 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1680363874
transform 1 0 2820 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1680363874
transform 1 0 2844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1680363874
transform 1 0 2852 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1568
timestamp 1680363874
transform 1 0 2852 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1858
timestamp 1680363874
transform 1 0 2868 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1459
timestamp 1680363874
transform 1 0 2876 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1695
timestamp 1680363874
transform 1 0 2876 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1569
timestamp 1680363874
transform 1 0 2884 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1680363874
transform 1 0 2924 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1808
timestamp 1680363874
transform 1 0 2924 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1680363874
transform 1 0 2940 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1680363874
transform 1 0 2948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1680363874
transform 1 0 2956 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1529
timestamp 1680363874
transform 1 0 2980 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1859
timestamp 1680363874
transform 1 0 2980 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1680363874
transform 1 0 2996 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1530
timestamp 1680363874
transform 1 0 3012 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1680363874
transform 1 0 2996 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1860
timestamp 1680363874
transform 1 0 3012 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1621
timestamp 1680363874
transform 1 0 3012 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1811
timestamp 1680363874
transform 1 0 3028 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1571
timestamp 1680363874
transform 1 0 3028 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1680363874
transform 1 0 3060 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1698
timestamp 1680363874
transform 1 0 3052 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1680363874
transform 1 0 3060 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1531
timestamp 1680363874
transform 1 0 3052 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1680363874
transform 1 0 3044 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1680363874
transform 1 0 3060 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1861
timestamp 1680363874
transform 1 0 3084 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1623
timestamp 1680363874
transform 1 0 3084 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1700
timestamp 1680363874
transform 1 0 3108 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1460
timestamp 1680363874
transform 1 0 3164 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1680363874
transform 1 0 3196 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1680363874
transform 1 0 3132 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1701
timestamp 1680363874
transform 1 0 3196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1680363874
transform 1 0 3116 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1680363874
transform 1 0 3172 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1572
timestamp 1680363874
transform 1 0 3172 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1680363874
transform 1 0 3116 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1680363874
transform 1 0 3196 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1680363874
transform 1 0 3180 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1680363874
transform 1 0 3212 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1814
timestamp 1680363874
transform 1 0 3212 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1573
timestamp 1680363874
transform 1 0 3212 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1680363874
transform 1 0 3228 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1680363874
transform 1 0 3220 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1680363874
transform 1 0 3252 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1680363874
transform 1 0 3308 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1702
timestamp 1680363874
transform 1 0 3284 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1680363874
transform 1 0 3292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1680363874
transform 1 0 3308 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1680363874
transform 1 0 3284 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1680363874
transform 1 0 3300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1680363874
transform 1 0 3316 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1574
timestamp 1680363874
transform 1 0 3284 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1680363874
transform 1 0 3292 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1680363874
transform 1 0 3316 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1680363874
transform 1 0 3316 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1680363874
transform 1 0 3356 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1680363874
transform 1 0 3372 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1705
timestamp 1680363874
transform 1 0 3380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1680363874
transform 1 0 3388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1680363874
transform 1 0 3356 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1680363874
transform 1 0 3372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1680363874
transform 1 0 3388 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1575
timestamp 1680363874
transform 1 0 3388 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1680363874
transform 1 0 3380 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1680363874
transform 1 0 3412 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1680363874
transform 1 0 3428 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1680363874
transform 1 0 3436 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1680363874
transform 1 0 3452 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1680363874
transform 1 0 3540 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1707
timestamp 1680363874
transform 1 0 3540 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1680363874
transform 1 0 3452 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1680363874
transform 1 0 3460 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1680363874
transform 1 0 3492 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1680363874
transform 1 0 3444 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1576
timestamp 1680363874
transform 1 0 3452 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1680363874
transform 1 0 3444 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1680363874
transform 1 0 3492 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1864
timestamp 1680363874
transform 1 0 3452 0 1 3905
box -2 -2 2 2
use M3_M2  M3_M2_1608
timestamp 1680363874
transform 1 0 3460 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1680363874
transform 1 0 3524 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1708
timestamp 1680363874
transform 1 0 3588 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1533
timestamp 1680363874
transform 1 0 3588 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1680363874
transform 1 0 3596 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1680363874
transform 1 0 3604 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1637
timestamp 1680363874
transform 1 0 3604 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1709
timestamp 1680363874
transform 1 0 3620 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1680363874
transform 1 0 3652 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1534
timestamp 1680363874
transform 1 0 3636 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1826
timestamp 1680363874
transform 1 0 3644 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1578
timestamp 1680363874
transform 1 0 3636 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1827
timestamp 1680363874
transform 1 0 3684 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1464
timestamp 1680363874
transform 1 0 3724 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1711
timestamp 1680363874
transform 1 0 3708 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1680363874
transform 1 0 3724 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1500
timestamp 1680363874
transform 1 0 3732 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1680363874
transform 1 0 3748 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1828
timestamp 1680363874
transform 1 0 3716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1680363874
transform 1 0 3732 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1680363874
transform 1 0 3740 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1579
timestamp 1680363874
transform 1 0 3708 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1680363874
transform 1 0 3732 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1680363874
transform 1 0 3716 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1680363874
transform 1 0 3804 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1680363874
transform 1 0 3828 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1680363874
transform 1 0 3860 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1680363874
transform 1 0 3852 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1680363874
transform 1 0 3820 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1680363874
transform 1 0 3844 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1713
timestamp 1680363874
transform 1 0 3820 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1680363874
transform 1 0 3828 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1680363874
transform 1 0 3844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1680363874
transform 1 0 3852 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1680363874
transform 1 0 3860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1680363874
transform 1 0 3836 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1680363874
transform 1 0 3860 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1680363874
transform 1 0 3868 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1638
timestamp 1680363874
transform 1 0 3868 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1680363874
transform 1 0 3916 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1680363874
transform 1 0 3948 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1718
timestamp 1680363874
transform 1 0 3924 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1680363874
transform 1 0 3940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1680363874
transform 1 0 3948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1680363874
transform 1 0 3956 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1535
timestamp 1680363874
transform 1 0 3924 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1834
timestamp 1680363874
transform 1 0 3932 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1611
timestamp 1680363874
transform 1 0 3948 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1835
timestamp 1680363874
transform 1 0 3988 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1581
timestamp 1680363874
transform 1 0 3988 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1680363874
transform 1 0 4004 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1722
timestamp 1680363874
transform 1 0 4004 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1680363874
transform 1 0 4020 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1680363874
transform 1 0 4028 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1680363874
transform 1 0 4012 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1536
timestamp 1680363874
transform 1 0 4020 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1837
timestamp 1680363874
transform 1 0 4028 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1468
timestamp 1680363874
transform 1 0 4044 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1838
timestamp 1680363874
transform 1 0 4116 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1537
timestamp 1680363874
transform 1 0 4132 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1680363874
transform 1 0 4156 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1680363874
transform 1 0 4196 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1725
timestamp 1680363874
transform 1 0 4156 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1680363874
transform 1 0 4172 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1680363874
transform 1 0 4188 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1680363874
transform 1 0 4196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1680363874
transform 1 0 4164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1680363874
transform 1 0 4180 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1612
timestamp 1680363874
transform 1 0 4180 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1680363874
transform 1 0 4164 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1841
timestamp 1680363874
transform 1 0 4196 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1582
timestamp 1680363874
transform 1 0 4196 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1680363874
transform 1 0 4212 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1729
timestamp 1680363874
transform 1 0 4236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1680363874
transform 1 0 4244 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1680363874
transform 1 0 4212 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1680363874
transform 1 0 4228 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1538
timestamp 1680363874
transform 1 0 4236 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1844
timestamp 1680363874
transform 1 0 4244 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1627
timestamp 1680363874
transform 1 0 4244 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1680363874
transform 1 0 4268 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1845
timestamp 1680363874
transform 1 0 4284 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1471
timestamp 1680363874
transform 1 0 4316 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1680363874
transform 1 0 4356 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1731
timestamp 1680363874
transform 1 0 4340 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1505
timestamp 1680363874
transform 1 0 4364 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1680363874
transform 1 0 4340 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1846
timestamp 1680363874
transform 1 0 4388 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1583
timestamp 1680363874
transform 1 0 4388 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1732
timestamp 1680363874
transform 1 0 4476 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1506
timestamp 1680363874
transform 1 0 4484 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1733
timestamp 1680363874
transform 1 0 4492 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1680363874
transform 1 0 4468 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1680363874
transform 1 0 4484 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1540
timestamp 1680363874
transform 1 0 4492 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1849
timestamp 1680363874
transform 1 0 4508 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1613
timestamp 1680363874
transform 1 0 4500 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1680363874
transform 1 0 4492 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1680363874
transform 1 0 4620 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1734
timestamp 1680363874
transform 1 0 4532 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1507
timestamp 1680363874
transform 1 0 4540 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1735
timestamp 1680363874
transform 1 0 4620 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1541
timestamp 1680363874
transform 1 0 4532 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1680363874
transform 1 0 4524 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1850
timestamp 1680363874
transform 1 0 4588 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1628
timestamp 1680363874
transform 1 0 4604 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1851
timestamp 1680363874
transform 1 0 4636 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1542
timestamp 1680363874
transform 1 0 4652 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1680363874
transform 1 0 4644 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1852
timestamp 1680363874
transform 1 0 4676 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1474
timestamp 1680363874
transform 1 0 4764 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1736
timestamp 1680363874
transform 1 0 4764 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1543
timestamp 1680363874
transform 1 0 4700 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1853
timestamp 1680363874
transform 1 0 4724 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1585
timestamp 1680363874
transform 1 0 4724 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1680363874
transform 1 0 4684 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1680363874
transform 1 0 4724 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1680363874
transform 1 0 4780 0 1 3945
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_16
timestamp 1680363874
transform 1 0 24 0 1 3870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_118
timestamp 1680363874
transform 1 0 72 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_108
timestamp 1680363874
transform 1 0 168 0 -1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1680363874
transform 1 0 184 0 -1 3970
box -8 -3 104 105
use M3_M2  M3_M2_1641
timestamp 1680363874
transform 1 0 324 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_91
timestamp 1680363874
transform 1 0 280 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1070
timestamp 1680363874
transform 1 0 320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1680363874
transform 1 0 328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1680363874
transform 1 0 336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1680363874
transform 1 0 344 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_92
timestamp 1680363874
transform 1 0 352 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1074
timestamp 1680363874
transform 1 0 392 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_110
timestamp 1680363874
transform 1 0 400 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1075
timestamp 1680363874
transform 1 0 416 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1680363874
transform 1 0 424 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1680363874
transform 1 0 432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1680363874
transform 1 0 440 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1642
timestamp 1680363874
transform 1 0 460 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_93
timestamp 1680363874
transform -1 0 488 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1079
timestamp 1680363874
transform 1 0 488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1680363874
transform 1 0 496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1680363874
transform 1 0 504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1680363874
transform 1 0 512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1680363874
transform 1 0 520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1680363874
transform 1 0 528 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1643
timestamp 1680363874
transform 1 0 548 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_95
timestamp 1680363874
transform 1 0 536 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1090
timestamp 1680363874
transform 1 0 576 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1680363874
transform 1 0 584 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1680363874
transform 1 0 592 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1680363874
transform 1 0 600 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_97
timestamp 1680363874
transform 1 0 608 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1099
timestamp 1680363874
transform 1 0 648 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1680363874
transform 1 0 656 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1644
timestamp 1680363874
transform 1 0 676 0 1 3875
box -3 -3 3 3
use FILL  FILL_1102
timestamp 1680363874
transform 1 0 664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1680363874
transform 1 0 672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1680363874
transform 1 0 680 0 -1 3970
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1680363874
transform 1 0 688 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1107
timestamp 1680363874
transform 1 0 712 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1680363874
transform 1 0 720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1680363874
transform 1 0 728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1680363874
transform 1 0 736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1680363874
transform 1 0 744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1680363874
transform 1 0 752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1680363874
transform 1 0 760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1680363874
transform 1 0 768 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_15
timestamp 1680363874
transform -1 0 808 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1123
timestamp 1680363874
transform 1 0 808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1680363874
transform 1 0 816 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1680363874
transform 1 0 824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1680363874
transform 1 0 832 0 -1 3970
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1680363874
transform -1 0 864 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1131
timestamp 1680363874
transform 1 0 864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1680363874
transform 1 0 872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1680363874
transform 1 0 880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1680363874
transform 1 0 888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1680363874
transform 1 0 896 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1680363874
transform 1 0 904 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1680363874
transform -1 0 944 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1153
timestamp 1680363874
transform 1 0 944 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1680363874
transform 1 0 952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1680363874
transform 1 0 960 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1680363874
transform 1 0 968 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_101
timestamp 1680363874
transform 1 0 976 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1157
timestamp 1680363874
transform 1 0 1016 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1680363874
transform 1 0 1024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1680363874
transform 1 0 1032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1680363874
transform 1 0 1040 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_102
timestamp 1680363874
transform 1 0 1048 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1161
timestamp 1680363874
transform 1 0 1088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1680363874
transform 1 0 1096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1680363874
transform 1 0 1104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1680363874
transform 1 0 1112 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_103
timestamp 1680363874
transform 1 0 1120 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1165
timestamp 1680363874
transform 1 0 1160 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1680363874
transform 1 0 1168 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_104
timestamp 1680363874
transform 1 0 1176 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_111
timestamp 1680363874
transform -1 0 1232 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1167
timestamp 1680363874
transform 1 0 1232 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1680363874
transform 1 0 1240 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1680363874
transform 1 0 1248 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1680363874
transform 1 0 1256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1680363874
transform 1 0 1264 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_106
timestamp 1680363874
transform 1 0 1272 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1184
timestamp 1680363874
transform 1 0 1312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1680363874
transform 1 0 1320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1680363874
transform 1 0 1328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1680363874
transform 1 0 1336 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_107
timestamp 1680363874
transform -1 0 1384 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1188
timestamp 1680363874
transform 1 0 1384 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1680363874
transform 1 0 1392 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_108
timestamp 1680363874
transform 1 0 1400 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1680363874
transform 1 0 1440 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1190
timestamp 1680363874
transform 1 0 1536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1680363874
transform 1 0 1544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1680363874
transform 1 0 1552 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_114
timestamp 1680363874
transform -1 0 1576 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1680363874
transform -1 0 1592 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1193
timestamp 1680363874
transform 1 0 1592 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1680363874
transform 1 0 1600 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1680363874
transform 1 0 1608 0 -1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1680363874
transform 1 0 1616 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1198
timestamp 1680363874
transform 1 0 1640 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1680363874
transform 1 0 1648 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1680363874
transform 1 0 1656 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1680363874
transform 1 0 1664 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_117
timestamp 1680363874
transform 1 0 1672 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1207
timestamp 1680363874
transform 1 0 1688 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1680363874
transform 1 0 1696 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1680363874
transform 1 0 1704 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_68
timestamp 1680363874
transform -1 0 1752 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1214
timestamp 1680363874
transform 1 0 1752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1680363874
transform 1 0 1760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1680363874
transform 1 0 1768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1680363874
transform 1 0 1776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1680363874
transform 1 0 1784 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_118
timestamp 1680363874
transform -1 0 1808 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1225
timestamp 1680363874
transform 1 0 1808 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_69
timestamp 1680363874
transform 1 0 1816 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1226
timestamp 1680363874
transform 1 0 1856 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1680363874
transform 1 0 1864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1680363874
transform 1 0 1872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1680363874
transform 1 0 1880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1680363874
transform 1 0 1888 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_119
timestamp 1680363874
transform -1 0 1912 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1238
timestamp 1680363874
transform 1 0 1912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1680363874
transform 1 0 1920 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1680363874
transform 1 0 1928 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_70
timestamp 1680363874
transform -1 0 1976 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1249
timestamp 1680363874
transform 1 0 1976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1680363874
transform 1 0 1984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1680363874
transform 1 0 1992 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_120
timestamp 1680363874
transform -1 0 2016 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1257
timestamp 1680363874
transform 1 0 2016 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1680363874
transform 1 0 2024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1680363874
transform 1 0 2032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1680363874
transform 1 0 2040 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_71
timestamp 1680363874
transform -1 0 2088 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1270
timestamp 1680363874
transform 1 0 2088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1680363874
transform 1 0 2096 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_121
timestamp 1680363874
transform 1 0 2104 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1276
timestamp 1680363874
transform 1 0 2120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1680363874
transform 1 0 2128 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1680363874
transform 1 0 2136 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1680363874
transform 1 0 2144 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1680363874
transform 1 0 2152 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1680363874
transform 1 0 2160 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1680363874
transform 1 0 2168 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1680363874
transform 1 0 2176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1680363874
transform 1 0 2184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1680363874
transform 1 0 2192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1680363874
transform 1 0 2200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1680363874
transform 1 0 2208 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1680363874
transform 1 0 2216 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1680363874
transform 1 0 2224 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1680363874
transform 1 0 2232 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1680363874
transform 1 0 2240 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1680363874
transform 1 0 2248 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1680363874
transform 1 0 2256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1680363874
transform 1 0 2264 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_124
timestamp 1680363874
transform 1 0 2272 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1311
timestamp 1680363874
transform 1 0 2288 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1680363874
transform 1 0 2296 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_125
timestamp 1680363874
transform 1 0 2304 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1313
timestamp 1680363874
transform 1 0 2320 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1645
timestamp 1680363874
transform 1 0 2340 0 1 3875
box -3 -3 3 3
use FILL  FILL_1314
timestamp 1680363874
transform 1 0 2328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1680363874
transform 1 0 2336 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1646
timestamp 1680363874
transform 1 0 2372 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_74
timestamp 1680363874
transform -1 0 2384 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1316
timestamp 1680363874
transform 1 0 2384 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1680363874
transform 1 0 2392 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1680363874
transform 1 0 2400 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1680363874
transform 1 0 2408 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_75
timestamp 1680363874
transform -1 0 2456 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1320
timestamp 1680363874
transform 1 0 2456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1680363874
transform 1 0 2464 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1680363874
transform 1 0 2472 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_129
timestamp 1680363874
transform 1 0 2480 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1337
timestamp 1680363874
transform 1 0 2496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1680363874
transform 1 0 2504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1680363874
transform 1 0 2512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1680363874
transform 1 0 2520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1680363874
transform 1 0 2528 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1680363874
transform 1 0 2536 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1342
timestamp 1680363874
transform 1 0 2632 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1680363874
transform 1 0 2640 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1680363874
transform 1 0 2648 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1647
timestamp 1680363874
transform 1 0 2668 0 1 3875
box -3 -3 3 3
use FILL  FILL_1345
timestamp 1680363874
transform 1 0 2656 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1680363874
transform 1 0 2664 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1648
timestamp 1680363874
transform 1 0 2740 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_130
timestamp 1680363874
transform 1 0 2672 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_130
timestamp 1680363874
transform 1 0 2768 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1347
timestamp 1680363874
transform 1 0 2784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1680363874
transform 1 0 2792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1680363874
transform 1 0 2800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1680363874
transform 1 0 2808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1680363874
transform 1 0 2816 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_110
timestamp 1680363874
transform 1 0 2824 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1352
timestamp 1680363874
transform 1 0 2864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1680363874
transform 1 0 2872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1680363874
transform 1 0 2880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1680363874
transform 1 0 2888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1680363874
transform 1 0 2896 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1680363874
transform 1 0 2904 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1680363874
transform 1 0 2912 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1365
timestamp 1680363874
transform 1 0 2944 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1680363874
transform 1 0 2952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1680363874
transform 1 0 2960 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1680363874
transform 1 0 2968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1680363874
transform 1 0 2976 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_22
timestamp 1680363874
transform 1 0 2984 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1375
timestamp 1680363874
transform 1 0 3016 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1680363874
transform 1 0 3024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1680363874
transform 1 0 3032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1680363874
transform 1 0 3040 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1680363874
transform 1 0 3048 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1680363874
transform 1 0 3056 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1392
timestamp 1680363874
transform 1 0 3088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1680363874
transform 1 0 3096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1680363874
transform 1 0 3104 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1649
timestamp 1680363874
transform 1 0 3156 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1680363874
transform 1 0 3188 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_131
timestamp 1680363874
transform -1 0 3208 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1395
timestamp 1680363874
transform 1 0 3208 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1680363874
transform 1 0 3216 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1651
timestamp 1680363874
transform 1 0 3236 0 1 3875
box -3 -3 3 3
use FILL  FILL_1399
timestamp 1680363874
transform 1 0 3224 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1680363874
transform 1 0 3232 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_132
timestamp 1680363874
transform -1 0 3256 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1415
timestamp 1680363874
transform 1 0 3256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1680363874
transform 1 0 3264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1680363874
transform 1 0 3272 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_79
timestamp 1680363874
transform -1 0 3320 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1418
timestamp 1680363874
transform 1 0 3320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1680363874
transform 1 0 3328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1680363874
transform 1 0 3336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1680363874
transform 1 0 3344 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1652
timestamp 1680363874
transform 1 0 3372 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_80
timestamp 1680363874
transform 1 0 3352 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1422
timestamp 1680363874
transform 1 0 3392 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1680363874
transform 1 0 3400 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1680363874
transform 1 0 3408 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1680363874
transform 1 0 3416 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1680363874
transform 1 0 3424 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1426
timestamp 1680363874
transform 1 0 3440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1680363874
transform 1 0 3448 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1653
timestamp 1680363874
transform 1 0 3484 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_133
timestamp 1680363874
transform -1 0 3552 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1428
timestamp 1680363874
transform 1 0 3552 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1680363874
transform 1 0 3560 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1654
timestamp 1680363874
transform 1 0 3580 0 1 3875
box -3 -3 3 3
use FILL  FILL_1432
timestamp 1680363874
transform 1 0 3568 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1680363874
transform 1 0 3576 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_134
timestamp 1680363874
transform 1 0 3584 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1438
timestamp 1680363874
transform 1 0 3600 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1680363874
transform 1 0 3608 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1680363874
transform 1 0 3616 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_81
timestamp 1680363874
transform -1 0 3664 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1447
timestamp 1680363874
transform 1 0 3664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1680363874
transform 1 0 3672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1680363874
transform 1 0 3680 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1680363874
transform 1 0 3688 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1655
timestamp 1680363874
transform 1 0 3708 0 1 3875
box -3 -3 3 3
use FILL  FILL_1456
timestamp 1680363874
transform 1 0 3696 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1656
timestamp 1680363874
transform 1 0 3740 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_111
timestamp 1680363874
transform -1 0 3744 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1457
timestamp 1680363874
transform 1 0 3744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1680363874
transform 1 0 3752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1680363874
transform 1 0 3760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1680363874
transform 1 0 3768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1680363874
transform 1 0 3776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1680363874
transform 1 0 3784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1680363874
transform 1 0 3792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1680363874
transform 1 0 3800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1680363874
transform 1 0 3808 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_83
timestamp 1680363874
transform 1 0 3816 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1478
timestamp 1680363874
transform 1 0 3856 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1680363874
transform 1 0 3864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1680363874
transform 1 0 3872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1680363874
transform 1 0 3880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1680363874
transform 1 0 3888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1680363874
transform 1 0 3896 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1680363874
transform 1 0 3904 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_84
timestamp 1680363874
transform 1 0 3912 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1485
timestamp 1680363874
transform 1 0 3952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1680363874
transform 1 0 3960 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1680363874
transform 1 0 3968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1680363874
transform 1 0 3976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1680363874
transform 1 0 3984 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_85
timestamp 1680363874
transform -1 0 4032 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1498
timestamp 1680363874
transform 1 0 4032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1680363874
transform 1 0 4040 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1680363874
transform 1 0 4048 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_137
timestamp 1680363874
transform 1 0 4056 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1505
timestamp 1680363874
transform 1 0 4072 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1680363874
transform 1 0 4080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1680363874
transform 1 0 4088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1680363874
transform 1 0 4096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1680363874
transform 1 0 4104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1680363874
transform 1 0 4112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1680363874
transform 1 0 4120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1680363874
transform 1 0 4128 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1680363874
transform 1 0 4136 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1680363874
transform 1 0 4144 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_112
timestamp 1680363874
transform 1 0 4152 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1515
timestamp 1680363874
transform 1 0 4192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1680363874
transform 1 0 4200 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_86
timestamp 1680363874
transform -1 0 4248 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1521
timestamp 1680363874
transform 1 0 4248 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1680363874
transform 1 0 4256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1680363874
transform 1 0 4264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1680363874
transform 1 0 4272 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_138
timestamp 1680363874
transform 1 0 4280 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1525
timestamp 1680363874
transform 1 0 4296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1680363874
transform 1 0 4304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1680363874
transform 1 0 4312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1680363874
transform 1 0 4320 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_138
timestamp 1680363874
transform 1 0 4328 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1541
timestamp 1680363874
transform 1 0 4424 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1680363874
transform 1 0 4432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1680363874
transform 1 0 4440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1680363874
transform 1 0 4448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1680363874
transform 1 0 4456 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_87
timestamp 1680363874
transform -1 0 4504 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1546
timestamp 1680363874
transform 1 0 4504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1680363874
transform 1 0 4512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1680363874
transform 1 0 4520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1680363874
transform 1 0 4528 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1680363874
transform -1 0 4632 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1550
timestamp 1680363874
transform 1 0 4632 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1680363874
transform 1 0 4640 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1680363874
transform 1 0 4648 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1680363874
transform 1 0 4656 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1680363874
transform 1 0 4664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1680363874
transform 1 0 4672 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1680363874
transform -1 0 4776 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1574
timestamp 1680363874
transform 1 0 4776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1680363874
transform 1 0 4784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1680363874
transform 1 0 4792 0 -1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_17
timestamp 1680363874
transform 1 0 4851 0 1 3870
box -10 -3 10 3
use M3_M2  M3_M2_1683
timestamp 1680363874
transform 1 0 172 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1872
timestamp 1680363874
transform 1 0 84 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1680363874
transform 1 0 140 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1755
timestamp 1680363874
transform 1 0 140 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1987
timestamp 1680363874
transform 1 0 164 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1772
timestamp 1680363874
transform 1 0 164 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1680363874
transform 1 0 188 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1874
timestamp 1680363874
transform 1 0 180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1680363874
transform 1 0 196 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1703
timestamp 1680363874
transform 1 0 228 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1875
timestamp 1680363874
transform 1 0 228 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1756
timestamp 1680363874
transform 1 0 212 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1989
timestamp 1680363874
transform 1 0 220 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1757
timestamp 1680363874
transform 1 0 228 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1990
timestamp 1680363874
transform 1 0 236 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1704
timestamp 1680363874
transform 1 0 252 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1680363874
transform 1 0 332 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1680363874
transform 1 0 380 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1876
timestamp 1680363874
transform 1 0 332 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1680363874
transform 1 0 380 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1680363874
transform 1 0 300 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1773
timestamp 1680363874
transform 1 0 300 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1680363874
transform 1 0 492 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1680363874
transform 1 0 460 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1878
timestamp 1680363874
transform 1 0 460 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1680363874
transform 1 0 420 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1680363874
transform 1 0 508 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1680363874
transform 1 0 524 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1685
timestamp 1680363874
transform 1 0 540 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1680363874
transform 1 0 572 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1680363874
transform 1 0 548 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1880
timestamp 1680363874
transform 1 0 540 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1680363874
transform 1 0 556 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1680363874
transform 1 0 572 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1680363874
transform 1 0 532 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1680363874
transform 1 0 548 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1774
timestamp 1680363874
transform 1 0 524 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1680363874
transform 1 0 556 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1996
timestamp 1680363874
transform 1 0 564 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1680363874
transform 1 0 572 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1775
timestamp 1680363874
transform 1 0 572 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1883
timestamp 1680363874
transform 1 0 628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1680363874
transform 1 0 644 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1687
timestamp 1680363874
transform 1 0 660 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1998
timestamp 1680363874
transform 1 0 636 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1680363874
transform 1 0 652 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1680363874
transform 1 0 660 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1819
timestamp 1680363874
transform 1 0 636 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1885
timestamp 1680363874
transform 1 0 676 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1709
timestamp 1680363874
transform 1 0 716 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1680363874
transform 1 0 692 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1886
timestamp 1680363874
transform 1 0 716 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1734
timestamp 1680363874
transform 1 0 732 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2001
timestamp 1680363874
transform 1 0 708 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1680363874
transform 1 0 724 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1680363874
transform 1 0 732 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1776
timestamp 1680363874
transform 1 0 708 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1680363874
transform 1 0 780 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1865
timestamp 1680363874
transform 1 0 764 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1710
timestamp 1680363874
transform 1 0 772 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1680363874
transform 1 0 764 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2004
timestamp 1680363874
transform 1 0 788 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1680363874
transform 1 0 796 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1777
timestamp 1680363874
transform 1 0 796 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1680363874
transform 1 0 820 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1887
timestamp 1680363874
transform 1 0 820 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1680363874
transform 1 0 836 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1759
timestamp 1680363874
transform 1 0 836 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1866
timestamp 1680363874
transform 1 0 860 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1680363874
transform 1 0 924 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1680363874
transform 1 0 924 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1820
timestamp 1680363874
transform 1 0 924 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1868
timestamp 1680363874
transform 1 0 972 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1680363874
transform 1 0 948 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1680363874
transform 1 0 956 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1736
timestamp 1680363874
transform 1 0 972 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1680363874
transform 1 0 956 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1680363874
transform 1 0 988 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1891
timestamp 1680363874
transform 1 0 996 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1680363874
transform 1 0 1020 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1712
timestamp 1680363874
transform 1 0 1068 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1680363874
transform 1 0 1044 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1892
timestamp 1680363874
transform 1 0 1052 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1680363874
transform 1 0 1068 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1680363874
transform 1 0 1076 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1680363874
transform 1 0 1084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1680363874
transform 1 0 1044 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1680363874
transform 1 0 1060 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1779
timestamp 1680363874
transform 1 0 1060 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1680363874
transform 1 0 1108 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1680363874
transform 1 0 1140 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1680363874
transform 1 0 1148 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1896
timestamp 1680363874
transform 1 0 1132 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1738
timestamp 1680363874
transform 1 0 1140 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1897
timestamp 1680363874
transform 1 0 1148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1680363874
transform 1 0 1108 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1760
timestamp 1680363874
transform 1 0 1116 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2010
timestamp 1680363874
transform 1 0 1124 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1680363874
transform 1 0 1140 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1680363874
transform 1 0 1188 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1680363874
transform 1 0 1164 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1680363874
transform 1 0 1180 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1780
timestamp 1680363874
transform 1 0 1180 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2014
timestamp 1680363874
transform 1 0 1204 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1680363874
transform 1 0 1244 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1680363874
transform 1 0 1220 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1781
timestamp 1680363874
transform 1 0 1244 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1680363874
transform 1 0 1220 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1680363874
transform 1 0 1268 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1680363874
transform 1 0 1300 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1680363874
transform 1 0 1316 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1680363874
transform 1 0 1332 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1900
timestamp 1680363874
transform 1 0 1324 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1680363874
transform 1 0 1332 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1680363874
transform 1 0 1348 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1680363874
transform 1 0 1340 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1680363874
transform 1 0 1348 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1761
timestamp 1680363874
transform 1 0 1364 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1903
timestamp 1680363874
transform 1 0 1380 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1680363874
transform 1 0 1372 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1716
timestamp 1680363874
transform 1 0 1420 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1904
timestamp 1680363874
transform 1 0 1420 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1740
timestamp 1680363874
transform 1 0 1428 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1680363874
transform 1 0 1468 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1762
timestamp 1680363874
transform 1 0 1468 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2019
timestamp 1680363874
transform 1 0 1516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1782
timestamp 1680363874
transform 1 0 1452 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1680363874
transform 1 0 1516 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1680363874
transform 1 0 1564 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1906
timestamp 1680363874
transform 1 0 1564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1680363874
transform 1 0 1620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1680363874
transform 1 0 1540 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1763
timestamp 1680363874
transform 1 0 1564 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1680363874
transform 1 0 1540 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1680363874
transform 1 0 1572 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1680363874
transform 1 0 1636 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1680363874
transform 1 0 1700 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1764
timestamp 1680363874
transform 1 0 1668 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2021
timestamp 1680363874
transform 1 0 1732 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1786
timestamp 1680363874
transform 1 0 1732 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1680363874
transform 1 0 1756 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1680363874
transform 1 0 1772 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1910
timestamp 1680363874
transform 1 0 1796 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1680363874
transform 1 0 1772 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1788
timestamp 1680363874
transform 1 0 1772 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1911
timestamp 1680363874
transform 1 0 1860 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1676
timestamp 1680363874
transform 1 0 1916 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1680363874
transform 1 0 1876 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1912
timestamp 1680363874
transform 1 0 1900 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1680363874
transform 1 0 1956 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1680363874
transform 1 0 1876 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1789
timestamp 1680363874
transform 1 0 1876 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1680363874
transform 1 0 1908 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1680363874
transform 1 0 1964 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1680363874
transform 1 0 1980 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1914
timestamp 1680363874
transform 1 0 2004 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1744
timestamp 1680363874
transform 1 0 2012 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1915
timestamp 1680363874
transform 1 0 2060 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1680363874
transform 1 0 1980 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1792
timestamp 1680363874
transform 1 0 1980 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1680363874
transform 1 0 2124 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1680363874
transform 1 0 2172 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1680363874
transform 1 0 2164 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1680363874
transform 1 0 2132 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1680363874
transform 1 0 2172 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1916
timestamp 1680363874
transform 1 0 2132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1680363874
transform 1 0 2164 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1680363874
transform 1 0 2172 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1680363874
transform 1 0 2084 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1793
timestamp 1680363874
transform 1 0 2084 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1919
timestamp 1680363874
transform 1 0 2204 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1691
timestamp 1680363874
transform 1 0 2228 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1920
timestamp 1680363874
transform 1 0 2236 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1745
timestamp 1680363874
transform 1 0 2244 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1921
timestamp 1680363874
transform 1 0 2252 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1680363874
transform 1 0 2220 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1680363874
transform 1 0 2228 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1794
timestamp 1680363874
transform 1 0 2244 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1680363874
transform 1 0 2228 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_2028
timestamp 1680363874
transform 1 0 2260 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1657
timestamp 1680363874
transform 1 0 2340 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1680363874
transform 1 0 2300 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1680363874
transform 1 0 2364 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1680363874
transform 1 0 2356 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1680363874
transform 1 0 2380 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1922
timestamp 1680363874
transform 1 0 2316 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1680363874
transform 1 0 2372 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1680363874
transform 1 0 2292 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1795
timestamp 1680363874
transform 1 0 2292 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1680363874
transform 1 0 2332 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1924
timestamp 1680363874
transform 1 0 2388 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1680363874
transform 1 0 2396 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1826
timestamp 1680363874
transform 1 0 2404 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1925
timestamp 1680363874
transform 1 0 2420 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1680363874
transform 1 0 2428 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1827
timestamp 1680363874
transform 1 0 2420 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1680363874
transform 1 0 2476 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1680363874
transform 1 0 2500 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1926
timestamp 1680363874
transform 1 0 2492 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1680363874
transform 1 0 2516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1796
timestamp 1680363874
transform 1 0 2500 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1680363874
transform 1 0 2532 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1680363874
transform 1 0 2540 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_2032
timestamp 1680363874
transform 1 0 2540 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1680363874
transform 1 0 2564 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1680363874
transform 1 0 2572 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1680363874
transform 1 0 2580 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1927
timestamp 1680363874
transform 1 0 2556 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1680363874
transform 1 0 2564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1680363874
transform 1 0 2580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1680363874
transform 1 0 2596 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1680363874
transform 1 0 2572 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1680363874
transform 1 0 2588 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1680363874
transform 1 0 2596 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1693
timestamp 1680363874
transform 1 0 2628 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1680363874
transform 1 0 2676 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1931
timestamp 1680363874
transform 1 0 2628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1680363874
transform 1 0 2684 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1746
timestamp 1680363874
transform 1 0 2708 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1680363874
transform 1 0 2732 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1680363874
transform 1 0 2764 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1680363874
transform 1 0 2804 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1933
timestamp 1680363874
transform 1 0 2732 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1680363874
transform 1 0 2748 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1680363874
transform 1 0 2764 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1680363874
transform 1 0 2788 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1680363874
transform 1 0 2804 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1680363874
transform 1 0 2708 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1680363874
transform 1 0 2724 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1680363874
transform 1 0 2740 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1680363874
transform 1 0 2756 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1680363874
transform 1 0 2764 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1680363874
transform 1 0 2780 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1680363874
transform 1 0 2796 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1798
timestamp 1680363874
transform 1 0 2708 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1680363874
transform 1 0 2756 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1680363874
transform 1 0 2804 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1680363874
transform 1 0 2796 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1938
timestamp 1680363874
transform 1 0 2852 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1726
timestamp 1680363874
transform 1 0 2868 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1939
timestamp 1680363874
transform 1 0 2868 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1680363874
transform 1 0 2828 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1680363874
transform 1 0 2844 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1680363874
transform 1 0 2860 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1801
timestamp 1680363874
transform 1 0 2860 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2046
timestamp 1680363874
transform 1 0 2876 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1680363874
transform 1 0 2916 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1680363874
transform 1 0 2932 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1680363874
transform 1 0 2908 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1680363874
transform 1 0 2924 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1802
timestamp 1680363874
transform 1 0 2924 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1942
timestamp 1680363874
transform 1 0 2956 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1680363874
transform 1 0 2980 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1680363874
transform 1 0 2996 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1680363874
transform 1 0 3020 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1680363874
transform 1 0 3036 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1680363874
transform 1 0 3012 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1766
timestamp 1680363874
transform 1 0 3020 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2051
timestamp 1680363874
transform 1 0 3028 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1694
timestamp 1680363874
transform 1 0 3140 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1946
timestamp 1680363874
transform 1 0 3084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1680363874
transform 1 0 3140 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1680363874
transform 1 0 3076 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1747
timestamp 1680363874
transform 1 0 3164 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2053
timestamp 1680363874
transform 1 0 3164 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1803
timestamp 1680363874
transform 1 0 3124 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1680363874
transform 1 0 3164 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1680363874
transform 1 0 3092 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1948
timestamp 1680363874
transform 1 0 3188 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1748
timestamp 1680363874
transform 1 0 3204 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2054
timestamp 1680363874
transform 1 0 3196 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1680363874
transform 1 0 3228 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1727
timestamp 1680363874
transform 1 0 3244 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1680363874
transform 1 0 3292 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1949
timestamp 1680363874
transform 1 0 3268 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1680363874
transform 1 0 3284 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1680363874
transform 1 0 3292 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1680363874
transform 1 0 3244 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1680363874
transform 1 0 3252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1680363874
transform 1 0 3260 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1680363874
transform 1 0 3276 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1805
timestamp 1680363874
transform 1 0 3268 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1680363874
transform 1 0 3276 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1680363874
transform 1 0 3332 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1871
timestamp 1680363874
transform 1 0 3348 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1680363874
transform 1 0 3340 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1806
timestamp 1680363874
transform 1 0 3340 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1952
timestamp 1680363874
transform 1 0 3436 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1680363874
transform 1 0 3420 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1830
timestamp 1680363874
transform 1 0 3420 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_2061
timestamp 1680363874
transform 1 0 3444 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1749
timestamp 1680363874
transform 1 0 3460 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1953
timestamp 1680363874
transform 1 0 3468 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1680363874
transform 1 0 3484 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1680363874
transform 1 0 3500 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1750
timestamp 1680363874
transform 1 0 3508 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1956
timestamp 1680363874
transform 1 0 3524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1680363874
transform 1 0 3484 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1680363874
transform 1 0 3508 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1680363874
transform 1 0 3516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1668
timestamp 1680363874
transform 1 0 3532 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1680363874
transform 1 0 3540 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1680363874
transform 1 0 3628 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1680363874
transform 1 0 3620 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1680363874
transform 1 0 3652 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1957
timestamp 1680363874
transform 1 0 3556 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1752
timestamp 1680363874
transform 1 0 3572 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1958
timestamp 1680363874
transform 1 0 3604 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1680363874
transform 1 0 3652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1680363874
transform 1 0 3660 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1680363874
transform 1 0 3572 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1696
timestamp 1680363874
transform 1 0 3684 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1680363874
transform 1 0 3700 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1680363874
transform 1 0 3732 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1680363874
transform 1 0 3724 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1961
timestamp 1680363874
transform 1 0 3708 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1680363874
transform 1 0 3724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1680363874
transform 1 0 3716 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1680363874
transform 1 0 3732 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1807
timestamp 1680363874
transform 1 0 3724 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2068
timestamp 1680363874
transform 1 0 3748 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1680363874
transform 1 0 3756 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1808
timestamp 1680363874
transform 1 0 3748 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1680363874
transform 1 0 3812 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1680363874
transform 1 0 3852 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1680363874
transform 1 0 3900 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1680363874
transform 1 0 3804 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1680363874
transform 1 0 3844 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1964
timestamp 1680363874
transform 1 0 3804 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1680363874
transform 1 0 3812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1680363874
transform 1 0 3844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1680363874
transform 1 0 3892 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1809
timestamp 1680363874
transform 1 0 3844 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1680363874
transform 1 0 3868 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1680363874
transform 1 0 3892 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1967
timestamp 1680363874
transform 1 0 3916 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1680363874
transform 1 0 3948 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1680363874
transform 1 0 3924 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1680363874
transform 1 0 3940 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1767
timestamp 1680363874
transform 1 0 3956 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1680363874
transform 1 0 3964 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1660
timestamp 1680363874
transform 1 0 4028 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1969
timestamp 1680363874
transform 1 0 4044 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1680363874
transform 1 0 4076 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1812
timestamp 1680363874
transform 1 0 4076 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2074
timestamp 1680363874
transform 1 0 4092 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1813
timestamp 1680363874
transform 1 0 4108 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1680363874
transform 1 0 4156 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1970
timestamp 1680363874
transform 1 0 4148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1680363874
transform 1 0 4156 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1680363874
transform 1 0 4140 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1768
timestamp 1680363874
transform 1 0 4148 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1972
timestamp 1680363874
transform 1 0 4172 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1729
timestamp 1680363874
transform 1 0 4188 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1680363874
transform 1 0 4204 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2088
timestamp 1680363874
transform 1 0 4220 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1701
timestamp 1680363874
transform 1 0 4244 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1973
timestamp 1680363874
transform 1 0 4292 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1680363874
transform 1 0 4284 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1831
timestamp 1680363874
transform 1 0 4292 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_2089
timestamp 1680363874
transform 1 0 4308 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1730
timestamp 1680363874
transform 1 0 4332 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1680363874
transform 1 0 4324 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1974
timestamp 1680363874
transform 1 0 4332 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1680363874
transform 1 0 4324 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1680363874
transform 1 0 4340 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1681
timestamp 1680363874
transform 1 0 4380 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1680363874
transform 1 0 4404 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1680363874
transform 1 0 4404 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1975
timestamp 1680363874
transform 1 0 4364 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1680363874
transform 1 0 4420 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1680363874
transform 1 0 4444 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1814
timestamp 1680363874
transform 1 0 4412 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1680363874
transform 1 0 4428 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1680363874
transform 1 0 4508 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1680363874
transform 1 0 4484 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1977
timestamp 1680363874
transform 1 0 4484 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1680363874
transform 1 0 4500 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1732
timestamp 1680363874
transform 1 0 4516 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_2079
timestamp 1680363874
transform 1 0 4476 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1680363874
transform 1 0 4492 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1680363874
transform 1 0 4508 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1680363874
transform 1 0 4516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1816
timestamp 1680363874
transform 1 0 4508 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1979
timestamp 1680363874
transform 1 0 4524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1680363874
transform 1 0 4548 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1680363874
transform 1 0 4596 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1754
timestamp 1680363874
transform 1 0 4628 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2083
timestamp 1680363874
transform 1 0 4628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1680363874
transform 1 0 4652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1680363874
transform 1 0 4644 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1817
timestamp 1680363874
transform 1 0 4644 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1983
timestamp 1680363874
transform 1 0 4684 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1680363874
transform 1 0 4700 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1680363874
transform 1 0 4708 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1680363874
transform 1 0 4764 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1770
timestamp 1680363874
transform 1 0 4668 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2085
timestamp 1680363874
transform 1 0 4692 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1771
timestamp 1680363874
transform 1 0 4700 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2086
timestamp 1680363874
transform 1 0 4788 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1818
timestamp 1680363874
transform 1 0 4708 0 1 3795
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_18
timestamp 1680363874
transform 1 0 48 0 1 3770
box -10 -3 10 3
use FILL  FILL_1579
timestamp 1680363874
transform 1 0 72 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1680363874
transform -1 0 176 0 1 3770
box -8 -3 104 105
use FILL  FILL_1580
timestamp 1680363874
transform 1 0 176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1680363874
transform 1 0 184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1680363874
transform 1 0 192 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_114
timestamp 1680363874
transform 1 0 200 0 1 3770
box -8 -3 46 105
use FILL  FILL_1596
timestamp 1680363874
transform 1 0 240 0 1 3770
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1680363874
transform 1 0 248 0 1 3770
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1680363874
transform 1 0 256 0 1 3770
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1680363874
transform 1 0 264 0 1 3770
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1680363874
transform 1 0 272 0 1 3770
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1680363874
transform 1 0 280 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1680363874
transform 1 0 288 0 1 3770
box -8 -3 104 105
use FILL  FILL_1602
timestamp 1680363874
transform 1 0 384 0 1 3770
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1680363874
transform 1 0 392 0 1 3770
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1680363874
transform 1 0 400 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_143
timestamp 1680363874
transform 1 0 408 0 1 3770
box -8 -3 104 105
use FILL  FILL_1613
timestamp 1680363874
transform 1 0 504 0 1 3770
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1680363874
transform 1 0 512 0 1 3770
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1680363874
transform 1 0 520 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_118
timestamp 1680363874
transform 1 0 528 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_145
timestamp 1680363874
transform 1 0 568 0 1 3770
box -9 -3 26 105
use FILL  FILL_1617
timestamp 1680363874
transform 1 0 584 0 1 3770
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1680363874
transform 1 0 592 0 1 3770
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1680363874
transform 1 0 600 0 1 3770
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1680363874
transform 1 0 608 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1832
timestamp 1680363874
transform 1 0 652 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_120
timestamp 1680363874
transform 1 0 616 0 1 3770
box -8 -3 46 105
use FILL  FILL_1624
timestamp 1680363874
transform 1 0 656 0 1 3770
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1680363874
transform 1 0 664 0 1 3770
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1680363874
transform 1 0 672 0 1 3770
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1680363874
transform 1 0 680 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1833
timestamp 1680363874
transform 1 0 716 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_122
timestamp 1680363874
transform 1 0 688 0 1 3770
box -8 -3 46 105
use FILL  FILL_1634
timestamp 1680363874
transform 1 0 728 0 1 3770
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1680363874
transform 1 0 736 0 1 3770
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1680363874
transform 1 0 744 0 1 3770
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1680363874
transform 1 0 752 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_29
timestamp 1680363874
transform -1 0 792 0 1 3770
box -8 -3 34 105
use FILL  FILL_1642
timestamp 1680363874
transform 1 0 792 0 1 3770
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1680363874
transform 1 0 800 0 1 3770
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1680363874
transform 1 0 808 0 1 3770
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1680363874
transform 1 0 816 0 1 3770
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1680363874
transform 1 0 824 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_30
timestamp 1680363874
transform 1 0 832 0 1 3770
box -8 -3 34 105
use FILL  FILL_1652
timestamp 1680363874
transform 1 0 864 0 1 3770
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1680363874
transform 1 0 872 0 1 3770
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1680363874
transform 1 0 880 0 1 3770
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1680363874
transform 1 0 888 0 1 3770
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1680363874
transform 1 0 896 0 1 3770
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1680363874
transform 1 0 904 0 1 3770
box -8 -3 32 105
use FILL  FILL_1660
timestamp 1680363874
transform 1 0 928 0 1 3770
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1680363874
transform 1 0 936 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1680363874
transform 1 0 944 0 1 3770
box -8 -3 34 105
use FILL  FILL_1666
timestamp 1680363874
transform 1 0 976 0 1 3770
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1680363874
transform 1 0 984 0 1 3770
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1680363874
transform 1 0 992 0 1 3770
box -8 -3 32 105
use FILL  FILL_1670
timestamp 1680363874
transform 1 0 1016 0 1 3770
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1680363874
transform 1 0 1024 0 1 3770
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1680363874
transform 1 0 1032 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_125
timestamp 1680363874
transform -1 0 1080 0 1 3770
box -8 -3 46 105
use FILL  FILL_1675
timestamp 1680363874
transform 1 0 1080 0 1 3770
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1680363874
transform 1 0 1088 0 1 3770
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1680363874
transform 1 0 1096 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_127
timestamp 1680363874
transform 1 0 1104 0 1 3770
box -8 -3 46 105
use FILL  FILL_1682
timestamp 1680363874
transform 1 0 1144 0 1 3770
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1680363874
transform 1 0 1152 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1834
timestamp 1680363874
transform 1 0 1188 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_128
timestamp 1680363874
transform 1 0 1160 0 1 3770
box -8 -3 46 105
use FILL  FILL_1684
timestamp 1680363874
transform 1 0 1200 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1680363874
transform 1 0 1208 0 1 3770
box -8 -3 104 105
use FILL  FILL_1691
timestamp 1680363874
transform 1 0 1304 0 1 3770
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1680363874
transform 1 0 1312 0 1 3770
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1680363874
transform 1 0 1320 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_147
timestamp 1680363874
transform -1 0 1344 0 1 3770
box -9 -3 26 105
use FILL  FILL_1696
timestamp 1680363874
transform 1 0 1344 0 1 3770
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1680363874
transform 1 0 1352 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1835
timestamp 1680363874
transform 1 0 1372 0 1 3775
box -3 -3 3 3
use FILL  FILL_1698
timestamp 1680363874
transform 1 0 1360 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_148
timestamp 1680363874
transform 1 0 1368 0 1 3770
box -9 -3 26 105
use FILL  FILL_1699
timestamp 1680363874
transform 1 0 1384 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1836
timestamp 1680363874
transform 1 0 1404 0 1 3775
box -3 -3 3 3
use FILL  FILL_1700
timestamp 1680363874
transform 1 0 1392 0 1 3770
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1680363874
transform 1 0 1400 0 1 3770
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1680363874
transform 1 0 1408 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_149
timestamp 1680363874
transform -1 0 1432 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1680363874
transform -1 0 1528 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1680363874
transform 1 0 1528 0 1 3770
box -8 -3 104 105
use FILL  FILL_1703
timestamp 1680363874
transform 1 0 1624 0 1 3770
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1680363874
transform 1 0 1632 0 1 3770
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1680363874
transform 1 0 1640 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1837
timestamp 1680363874
transform 1 0 1748 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_149
timestamp 1680363874
transform -1 0 1744 0 1 3770
box -8 -3 104 105
use FILL  FILL_1706
timestamp 1680363874
transform 1 0 1744 0 1 3770
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1680363874
transform 1 0 1752 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1838
timestamp 1680363874
transform 1 0 1780 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_150
timestamp 1680363874
transform 1 0 1760 0 1 3770
box -8 -3 104 105
use FILL  FILL_1708
timestamp 1680363874
transform 1 0 1856 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1839
timestamp 1680363874
transform 1 0 1884 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1680363874
transform 1 0 1916 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_151
timestamp 1680363874
transform 1 0 1864 0 1 3770
box -8 -3 104 105
use FILL  FILL_1709
timestamp 1680363874
transform 1 0 1960 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1841
timestamp 1680363874
transform 1 0 2060 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_152
timestamp 1680363874
transform 1 0 1968 0 1 3770
box -8 -3 104 105
use FILL  FILL_1710
timestamp 1680363874
transform 1 0 2064 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1842
timestamp 1680363874
transform 1 0 2092 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_153
timestamp 1680363874
transform 1 0 2072 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_150
timestamp 1680363874
transform -1 0 2184 0 1 3770
box -9 -3 26 105
use FILL  FILL_1711
timestamp 1680363874
transform 1 0 2184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1680363874
transform 1 0 2192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1680363874
transform 1 0 2200 0 1 3770
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1680363874
transform 1 0 2208 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_88
timestamp 1680363874
transform -1 0 2256 0 1 3770
box -8 -3 46 105
use FILL  FILL_1715
timestamp 1680363874
transform 1 0 2256 0 1 3770
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1680363874
transform 1 0 2264 0 1 3770
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1680363874
transform 1 0 2272 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1680363874
transform 1 0 2280 0 1 3770
box -8 -3 104 105
use FILL  FILL_1761
timestamp 1680363874
transform 1 0 2376 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1680363874
transform -1 0 2408 0 1 3770
box -8 -3 32 105
use FILL  FILL_1762
timestamp 1680363874
transform 1 0 2408 0 1 3770
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1680363874
transform 1 0 2416 0 1 3770
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1680363874
transform 1 0 2424 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1680363874
transform -1 0 2528 0 1 3770
box -8 -3 104 105
use FILL  FILL_1765
timestamp 1680363874
transform 1 0 2528 0 1 3770
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1680363874
transform 1 0 2536 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_154
timestamp 1680363874
transform 1 0 2544 0 1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_91
timestamp 1680363874
transform -1 0 2600 0 1 3770
box -8 -3 46 105
use FILL  FILL_1767
timestamp 1680363874
transform 1 0 2600 0 1 3770
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1680363874
transform 1 0 2608 0 1 3770
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1680363874
transform 1 0 2616 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1680363874
transform -1 0 2720 0 1 3770
box -8 -3 104 105
use OAI22X1  OAI22X1_131
timestamp 1680363874
transform 1 0 2720 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_132
timestamp 1680363874
transform 1 0 2760 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_155
timestamp 1680363874
transform 1 0 2800 0 1 3770
box -9 -3 26 105
use FILL  FILL_1770
timestamp 1680363874
transform 1 0 2816 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_133
timestamp 1680363874
transform 1 0 2824 0 1 3770
box -8 -3 46 105
use FILL  FILL_1771
timestamp 1680363874
transform 1 0 2864 0 1 3770
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1680363874
transform 1 0 2872 0 1 3770
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1680363874
transform 1 0 2880 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_134
timestamp 1680363874
transform 1 0 2888 0 1 3770
box -8 -3 46 105
use FILL  FILL_1774
timestamp 1680363874
transform 1 0 2928 0 1 3770
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1680363874
transform 1 0 2936 0 1 3770
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1680363874
transform 1 0 2944 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_156
timestamp 1680363874
transform -1 0 2968 0 1 3770
box -9 -3 26 105
use FILL  FILL_1777
timestamp 1680363874
transform 1 0 2968 0 1 3770
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1680363874
transform 1 0 2976 0 1 3770
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1680363874
transform 1 0 2984 0 1 3770
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1680363874
transform 1 0 2992 0 1 3770
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1680363874
transform 1 0 3000 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_135
timestamp 1680363874
transform 1 0 3008 0 1 3770
box -8 -3 46 105
use FILL  FILL_1817
timestamp 1680363874
transform 1 0 3048 0 1 3770
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1680363874
transform 1 0 3056 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1843
timestamp 1680363874
transform 1 0 3076 0 1 3775
box -3 -3 3 3
use FILL  FILL_1822
timestamp 1680363874
transform 1 0 3064 0 1 3770
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1680363874
transform 1 0 3072 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_162
timestamp 1680363874
transform -1 0 3176 0 1 3770
box -8 -3 104 105
use FILL  FILL_1824
timestamp 1680363874
transform 1 0 3176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1680363874
transform 1 0 3184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1680363874
transform 1 0 3192 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_42
timestamp 1680363874
transform 1 0 3200 0 1 3770
box -8 -3 34 105
use FILL  FILL_1827
timestamp 1680363874
transform 1 0 3232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1680363874
transform 1 0 3240 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_93
timestamp 1680363874
transform 1 0 3248 0 1 3770
box -8 -3 46 105
use FILL  FILL_1829
timestamp 1680363874
transform 1 0 3288 0 1 3770
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1680363874
transform 1 0 3296 0 1 3770
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1680363874
transform 1 0 3304 0 1 3770
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1680363874
transform 1 0 3312 0 1 3770
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1680363874
transform 1 0 3320 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_157
timestamp 1680363874
transform -1 0 3344 0 1 3770
box -9 -3 26 105
use FILL  FILL_1848
timestamp 1680363874
transform 1 0 3344 0 1 3770
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1680363874
transform 1 0 3352 0 1 3770
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1680363874
transform 1 0 3360 0 1 3770
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1680363874
transform 1 0 3368 0 1 3770
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1680363874
transform 1 0 3376 0 1 3770
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1680363874
transform 1 0 3384 0 1 3770
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1680363874
transform 1 0 3392 0 1 3770
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1680363874
transform 1 0 3400 0 1 3770
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1680363874
transform 1 0 3408 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_44
timestamp 1680363874
transform -1 0 3448 0 1 3770
box -8 -3 34 105
use FILL  FILL_1863
timestamp 1680363874
transform 1 0 3448 0 1 3770
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1680363874
transform 1 0 3456 0 1 3770
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1680363874
transform 1 0 3464 0 1 3770
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1680363874
transform 1 0 3472 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_94
timestamp 1680363874
transform 1 0 3480 0 1 3770
box -8 -3 46 105
use FILL  FILL_1867
timestamp 1680363874
transform 1 0 3520 0 1 3770
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1680363874
transform 1 0 3528 0 1 3770
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1680363874
transform 1 0 3536 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_158
timestamp 1680363874
transform 1 0 3544 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1680363874
transform 1 0 3560 0 1 3770
box -8 -3 104 105
use FILL  FILL_1870
timestamp 1680363874
transform 1 0 3656 0 1 3770
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1680363874
transform 1 0 3664 0 1 3770
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1680363874
transform 1 0 3672 0 1 3770
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1680363874
transform 1 0 3680 0 1 3770
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1680363874
transform 1 0 3688 0 1 3770
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1680363874
transform 1 0 3696 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_95
timestamp 1680363874
transform 1 0 3704 0 1 3770
box -8 -3 46 105
use FILL  FILL_1895
timestamp 1680363874
transform 1 0 3744 0 1 3770
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1680363874
transform 1 0 3752 0 1 3770
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1680363874
transform 1 0 3760 0 1 3770
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1680363874
transform 1 0 3768 0 1 3770
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1680363874
transform 1 0 3776 0 1 3770
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1680363874
transform 1 0 3784 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_159
timestamp 1680363874
transform 1 0 3792 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1680363874
transform -1 0 3904 0 1 3770
box -8 -3 104 105
use FILL  FILL_1907
timestamp 1680363874
transform 1 0 3904 0 1 3770
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1680363874
transform 1 0 3912 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_136
timestamp 1680363874
transform 1 0 3920 0 1 3770
box -8 -3 46 105
use FILL  FILL_1913
timestamp 1680363874
transform 1 0 3960 0 1 3770
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1680363874
transform 1 0 3968 0 1 3770
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1680363874
transform 1 0 3976 0 1 3770
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1680363874
transform 1 0 3984 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1844
timestamp 1680363874
transform 1 0 4004 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1680363874
transform 1 0 4068 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1680363874
transform 1 0 4092 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_168
timestamp 1680363874
transform -1 0 4088 0 1 3770
box -8 -3 104 105
use FILL  FILL_1920
timestamp 1680363874
transform 1 0 4088 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_161
timestamp 1680363874
transform 1 0 4096 0 1 3770
box -9 -3 26 105
use FILL  FILL_1928
timestamp 1680363874
transform 1 0 4112 0 1 3770
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1680363874
transform 1 0 4120 0 1 3770
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1680363874
transform 1 0 4128 0 1 3770
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1680363874
transform 1 0 4136 0 1 3770
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1680363874
transform 1 0 4144 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1680363874
transform -1 0 4176 0 1 3770
box -8 -3 32 105
use FILL  FILL_1936
timestamp 1680363874
transform 1 0 4176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1680363874
transform 1 0 4184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1680363874
transform 1 0 4192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1680363874
transform 1 0 4200 0 1 3770
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1680363874
transform 1 0 4208 0 1 3770
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1680363874
transform 1 0 4216 0 1 3770
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1680363874
transform 1 0 4224 0 1 3770
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1680363874
transform 1 0 4232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1680363874
transform 1 0 4240 0 1 3770
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1680363874
transform 1 0 4248 0 1 3770
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1680363874
transform 1 0 4256 0 1 3770
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1680363874
transform 1 0 4264 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1680363874
transform -1 0 4296 0 1 3770
box -8 -3 32 105
use FILL  FILL_1948
timestamp 1680363874
transform 1 0 4296 0 1 3770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1680363874
transform 1 0 4304 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1680363874
transform -1 0 4336 0 1 3770
box -8 -3 32 105
use FILL  FILL_1959
timestamp 1680363874
transform 1 0 4336 0 1 3770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1680363874
transform 1 0 4344 0 1 3770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1680363874
transform 1 0 4352 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1680363874
transform -1 0 4456 0 1 3770
box -8 -3 104 105
use FILL  FILL_1966
timestamp 1680363874
transform 1 0 4456 0 1 3770
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1680363874
transform 1 0 4464 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_137
timestamp 1680363874
transform 1 0 4472 0 1 3770
box -8 -3 46 105
use FILL  FILL_1976
timestamp 1680363874
transform 1 0 4512 0 1 3770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1680363874
transform 1 0 4520 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_165
timestamp 1680363874
transform 1 0 4528 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1680363874
transform -1 0 4640 0 1 3770
box -8 -3 104 105
use FILL  FILL_1978
timestamp 1680363874
transform 1 0 4640 0 1 3770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1680363874
transform 1 0 4648 0 1 3770
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1680363874
transform 1 0 4656 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_101
timestamp 1680363874
transform -1 0 4704 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1680363874
transform -1 0 4800 0 1 3770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_19
timestamp 1680363874
transform 1 0 4827 0 1 3770
box -10 -3 10 3
use M2_M1  M2_M1_2099
timestamp 1680363874
transform 1 0 84 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1863
timestamp 1680363874
transform 1 0 196 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1680363874
transform 1 0 244 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1680363874
transform 1 0 236 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2100
timestamp 1680363874
transform 1 0 196 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1921
timestamp 1680363874
transform 1 0 204 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2101
timestamp 1680363874
transform 1 0 212 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1680363874
transform 1 0 228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1680363874
transform 1 0 204 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1680363874
transform 1 0 220 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1942
timestamp 1680363874
transform 1 0 228 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2210
timestamp 1680363874
transform 1 0 236 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1865
timestamp 1680363874
transform 1 0 284 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1680363874
transform 1 0 284 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2103
timestamp 1680363874
transform 1 0 244 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1680363874
transform 1 0 268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1680363874
transform 1 0 284 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1680363874
transform 1 0 292 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1680363874
transform 1 0 244 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1680363874
transform 1 0 252 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2212
timestamp 1680363874
transform 1 0 276 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2010
timestamp 1680363874
transform 1 0 244 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1680363874
transform 1 0 276 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1680363874
transform 1 0 348 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2107
timestamp 1680363874
transform 1 0 332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1680363874
transform 1 0 348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1680363874
transform 1 0 324 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1680363874
transform 1 0 340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1974
timestamp 1680363874
transform 1 0 324 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1680363874
transform 1 0 340 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2215
timestamp 1680363874
transform 1 0 356 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1975
timestamp 1680363874
transform 1 0 356 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2109
timestamp 1680363874
transform 1 0 380 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1944
timestamp 1680363874
transform 1 0 396 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1680363874
transform 1 0 468 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2110
timestamp 1680363874
transform 1 0 420 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1945
timestamp 1680363874
transform 1 0 420 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2216
timestamp 1680363874
transform 1 0 468 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1847
timestamp 1680363874
transform 1 0 556 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1680363874
transform 1 0 548 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2111
timestamp 1680363874
transform 1 0 532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1680363874
transform 1 0 548 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1680363874
transform 1 0 564 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1680363874
transform 1 0 572 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_2035
timestamp 1680363874
transform 1 0 516 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2217
timestamp 1680363874
transform 1 0 540 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1946
timestamp 1680363874
transform 1 0 548 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2218
timestamp 1680363874
transform 1 0 556 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2026
timestamp 1680363874
transform 1 0 556 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1680363874
transform 1 0 548 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1680363874
transform 1 0 572 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1680363874
transform 1 0 612 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1680363874
transform 1 0 644 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2115
timestamp 1680363874
transform 1 0 620 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1680363874
transform 1 0 636 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1680363874
transform 1 0 612 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1680363874
transform 1 0 628 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1922
timestamp 1680363874
transform 1 0 652 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1680363874
transform 1 0 676 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1680363874
transform 1 0 700 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1680363874
transform 1 0 708 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1680363874
transform 1 0 724 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2117
timestamp 1680363874
transform 1 0 684 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1680363874
transform 1 0 700 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1680363874
transform 1 0 716 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1947
timestamp 1680363874
transform 1 0 684 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2221
timestamp 1680363874
transform 1 0 708 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1976
timestamp 1680363874
transform 1 0 716 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1680363874
transform 1 0 692 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1680363874
transform 1 0 780 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2120
timestamp 1680363874
transform 1 0 780 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1924
timestamp 1680363874
transform 1 0 788 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1680363874
transform 1 0 804 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2121
timestamp 1680363874
transform 1 0 796 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1680363874
transform 1 0 804 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1680363874
transform 1 0 772 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1680363874
transform 1 0 788 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2027
timestamp 1680363874
transform 1 0 764 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1680363874
transform 1 0 796 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1680363874
transform 1 0 836 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2224
timestamp 1680363874
transform 1 0 836 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1680363874
transform 1 0 860 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1849
timestamp 1680363874
transform 1 0 892 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1680363874
transform 1 0 884 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1680363874
transform 1 0 908 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1680363874
transform 1 0 908 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1680363874
transform 1 0 908 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1950
timestamp 1680363874
transform 1 0 908 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2225
timestamp 1680363874
transform 1 0 916 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1680363874
transform 1 0 908 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1895
timestamp 1680363874
transform 1 0 956 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2226
timestamp 1680363874
transform 1 0 956 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1680363874
transform 1 0 972 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1680363874
transform 1 0 1028 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1868
timestamp 1680363874
transform 1 0 1052 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1680363874
transform 1 0 1068 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2124
timestamp 1680363874
transform 1 0 1052 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1680363874
transform 1 0 1068 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1680363874
transform 1 0 1044 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1680363874
transform 1 0 1060 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1680363874
transform 1 0 1076 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1680363874
transform 1 0 1084 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1869
timestamp 1680363874
transform 1 0 1156 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2126
timestamp 1680363874
transform 1 0 1124 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1926
timestamp 1680363874
transform 1 0 1132 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2127
timestamp 1680363874
transform 1 0 1140 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1680363874
transform 1 0 1156 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1680363874
transform 1 0 1148 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1977
timestamp 1680363874
transform 1 0 1124 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1680363874
transform 1 0 1156 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2232
timestamp 1680363874
transform 1 0 1164 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1952
timestamp 1680363874
transform 1 0 1172 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1680363874
transform 1 0 1164 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1680363874
transform 1 0 1172 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2129
timestamp 1680363874
transform 1 0 1300 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1680363874
transform 1 0 1252 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2014
timestamp 1680363874
transform 1 0 1252 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1680363874
transform 1 0 1276 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2234
timestamp 1680363874
transform 1 0 1316 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1870
timestamp 1680363874
transform 1 0 1388 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2130
timestamp 1680363874
transform 1 0 1348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1680363874
transform 1 0 1364 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1680363874
transform 1 0 1380 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1680363874
transform 1 0 1372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1680363874
transform 1 0 1388 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1979
timestamp 1680363874
transform 1 0 1404 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1680363874
transform 1 0 1492 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2133
timestamp 1680363874
transform 1 0 1516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1680363874
transform 1 0 1468 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1980
timestamp 1680363874
transform 1 0 1468 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2134
timestamp 1680363874
transform 1 0 1548 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1680363874
transform 1 0 1564 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1897
timestamp 1680363874
transform 1 0 1580 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2092
timestamp 1680363874
transform 1 0 1588 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1898
timestamp 1680363874
transform 1 0 1604 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2135
timestamp 1680363874
transform 1 0 1588 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1680363874
transform 1 0 1604 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1680363874
transform 1 0 1580 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1928
timestamp 1680363874
transform 1 0 1628 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2137
timestamp 1680363874
transform 1 0 1636 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1680363874
transform 1 0 1644 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1680363874
transform 1 0 1612 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1953
timestamp 1680363874
transform 1 0 1620 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2240
timestamp 1680363874
transform 1 0 1636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1954
timestamp 1680363874
transform 1 0 1644 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1680363874
transform 1 0 1668 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2139
timestamp 1680363874
transform 1 0 1668 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1680363874
transform 1 0 1756 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1680363874
transform 1 0 1660 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1680363874
transform 1 0 1676 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1680363874
transform 1 0 1612 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1981
timestamp 1680363874
transform 1 0 1636 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2316
timestamp 1680363874
transform 1 0 1644 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1982
timestamp 1680363874
transform 1 0 1660 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1680363874
transform 1 0 1684 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2243
timestamp 1680363874
transform 1 0 1732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1680363874
transform 1 0 1772 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1983
timestamp 1680363874
transform 1 0 1732 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1680363874
transform 1 0 1772 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1680363874
transform 1 0 1788 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2245
timestamp 1680363874
transform 1 0 1804 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1680363874
transform 1 0 1828 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1680363874
transform 1 0 1836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1680363874
transform 1 0 1852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1680363874
transform 1 0 1828 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1957
timestamp 1680363874
transform 1 0 1836 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2247
timestamp 1680363874
transform 1 0 1844 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1958
timestamp 1680363874
transform 1 0 1852 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1680363874
transform 1 0 1828 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2144
timestamp 1680363874
transform 1 0 1884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1680363874
transform 1 0 1892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1680363874
transform 1 0 1908 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1680363874
transform 1 0 1916 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1680363874
transform 1 0 1884 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1680363874
transform 1 0 1900 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1959
timestamp 1680363874
transform 1 0 1908 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1680363874
transform 1 0 1884 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2250
timestamp 1680363874
transform 1 0 1924 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1852
timestamp 1680363874
transform 1 0 1956 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2251
timestamp 1680363874
transform 1 0 1972 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1680363874
transform 1 0 1996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1680363874
transform 1 0 2020 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1680363874
transform 1 0 2052 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1680363874
transform 1 0 2092 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1680363874
transform 1 0 2116 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1680363874
transform 1 0 2108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1680363874
transform 1 0 2100 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1987
timestamp 1680363874
transform 1 0 2108 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2151
timestamp 1680363874
transform 1 0 2148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1680363874
transform 1 0 2140 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1988
timestamp 1680363874
transform 1 0 2140 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2152
timestamp 1680363874
transform 1 0 2180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1680363874
transform 1 0 2196 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1680363874
transform 1 0 2212 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1680363874
transform 1 0 2212 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1680363874
transform 1 0 2236 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1680363874
transform 1 0 2268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1680363874
transform 1 0 2276 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1680363874
transform 1 0 2260 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1929
timestamp 1680363874
transform 1 0 2324 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2095
timestamp 1680363874
transform 1 0 2340 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1680363874
transform 1 0 2332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1680363874
transform 1 0 2316 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1989
timestamp 1680363874
transform 1 0 2316 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1680363874
transform 1 0 2332 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2320
timestamp 1680363874
transform 1 0 2348 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1930
timestamp 1680363874
transform 1 0 2396 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2157
timestamp 1680363874
transform 1 0 2404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1680363874
transform 1 0 2412 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1680363874
transform 1 0 2412 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1899
timestamp 1680363874
transform 1 0 2428 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2257
timestamp 1680363874
transform 1 0 2420 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1680363874
transform 1 0 2436 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1991
timestamp 1680363874
transform 1 0 2420 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1680363874
transform 1 0 2436 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2159
timestamp 1680363874
transform 1 0 2452 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1900
timestamp 1680363874
transform 1 0 2476 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1680363874
transform 1 0 2516 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2160
timestamp 1680363874
transform 1 0 2476 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1680363874
transform 1 0 2524 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1680363874
transform 1 0 2556 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2037
timestamp 1680363874
transform 1 0 2516 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2161
timestamp 1680363874
transform 1 0 2596 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1871
timestamp 1680363874
transform 1 0 2628 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2162
timestamp 1680363874
transform 1 0 2620 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1680363874
transform 1 0 2572 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1680363874
transform 1 0 2588 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1680363874
transform 1 0 2604 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1680363874
transform 1 0 2612 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1993
timestamp 1680363874
transform 1 0 2604 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2096
timestamp 1680363874
transform 1 0 2636 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1872
timestamp 1680363874
transform 1 0 2716 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1680363874
transform 1 0 2724 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1680363874
transform 1 0 2772 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1680363874
transform 1 0 2804 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1680363874
transform 1 0 2820 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2163
timestamp 1680363874
transform 1 0 2804 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1874
timestamp 1680363874
transform 1 0 2900 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2164
timestamp 1680363874
transform 1 0 2900 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1931
timestamp 1680363874
transform 1 0 2948 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2265
timestamp 1680363874
transform 1 0 2836 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1680363874
transform 1 0 2884 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1680363874
transform 1 0 2924 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2016
timestamp 1680363874
transform 1 0 2964 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2165
timestamp 1680363874
transform 1 0 2988 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1680363874
transform 1 0 2996 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1680363874
transform 1 0 3012 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1994
timestamp 1680363874
transform 1 0 3004 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1680363874
transform 1 0 3036 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1680363874
transform 1 0 3028 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2270
timestamp 1680363874
transform 1 0 3044 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1680363874
transform 1 0 3036 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1680363874
transform 1 0 3060 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1904
timestamp 1680363874
transform 1 0 3068 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2167
timestamp 1680363874
transform 1 0 3068 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1996
timestamp 1680363874
transform 1 0 3060 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1680363874
transform 1 0 3076 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1680363874
transform 1 0 3100 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2168
timestamp 1680363874
transform 1 0 3092 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1934
timestamp 1680363874
transform 1 0 3100 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2169
timestamp 1680363874
transform 1 0 3108 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1680363874
transform 1 0 3092 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1680363874
transform 1 0 3100 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2028
timestamp 1680363874
transform 1 0 3084 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1680363874
transform 1 0 3124 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1680363874
transform 1 0 3156 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2273
timestamp 1680363874
transform 1 0 3148 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1680363874
transform 1 0 3180 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1855
timestamp 1680363874
transform 1 0 3260 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1680363874
transform 1 0 3252 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1680363874
transform 1 0 3204 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1680363874
transform 1 0 3268 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2170
timestamp 1680363874
transform 1 0 3268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1680363874
transform 1 0 3244 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1680363874
transform 1 0 3284 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_2029
timestamp 1680363874
transform 1 0 3284 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1680363874
transform 1 0 3300 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1680363874
transform 1 0 3308 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1680363874
transform 1 0 3308 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1680363874
transform 1 0 3324 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2171
timestamp 1680363874
transform 1 0 3380 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1935
timestamp 1680363874
transform 1 0 3388 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2275
timestamp 1680363874
transform 1 0 3396 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1936
timestamp 1680363874
transform 1 0 3412 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2276
timestamp 1680363874
transform 1 0 3412 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2018
timestamp 1680363874
transform 1 0 3428 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1680363874
transform 1 0 3444 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1680363874
transform 1 0 3468 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2098
timestamp 1680363874
transform 1 0 3476 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1680363874
transform 1 0 3460 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1680363874
transform 1 0 3476 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1876
timestamp 1680363874
transform 1 0 3492 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2173
timestamp 1680363874
transform 1 0 3500 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1911
timestamp 1680363874
transform 1 0 3572 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1680363874
transform 1 0 3596 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1680363874
transform 1 0 3596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1680363874
transform 1 0 3556 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1961
timestamp 1680363874
transform 1 0 3596 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1680363874
transform 1 0 3556 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1680363874
transform 1 0 3612 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1680363874
transform 1 0 3660 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2175
timestamp 1680363874
transform 1 0 3644 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1680363874
transform 1 0 3644 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1962
timestamp 1680363874
transform 1 0 3660 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2280
timestamp 1680363874
transform 1 0 3668 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1997
timestamp 1680363874
transform 1 0 3660 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2324
timestamp 1680363874
transform 1 0 3668 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_2039
timestamp 1680363874
transform 1 0 3644 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1680363874
transform 1 0 3684 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1680363874
transform 1 0 3724 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1680363874
transform 1 0 3716 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2176
timestamp 1680363874
transform 1 0 3716 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1680363874
transform 1 0 3724 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1680363874
transform 1 0 3756 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1680363874
transform 1 0 3732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1680363874
transform 1 0 3748 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2020
timestamp 1680363874
transform 1 0 3748 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2283
timestamp 1680363874
transform 1 0 3764 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1680363874
transform 1 0 3884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1680363874
transform 1 0 3836 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1998
timestamp 1680363874
transform 1 0 3844 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1680363874
transform 1 0 3844 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1680363874
transform 1 0 3900 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2180
timestamp 1680363874
transform 1 0 3900 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1680363874
transform 1 0 3900 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1999
timestamp 1680363874
transform 1 0 3900 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1680363874
transform 1 0 3916 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1680363874
transform 1 0 3940 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1680363874
transform 1 0 3956 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1680363874
transform 1 0 3932 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2181
timestamp 1680363874
transform 1 0 3932 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1680363874
transform 1 0 3948 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1680363874
transform 1 0 3956 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1680363874
transform 1 0 3940 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1963
timestamp 1680363874
transform 1 0 3948 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2287
timestamp 1680363874
transform 1 0 3956 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1964
timestamp 1680363874
transform 1 0 3964 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1680363874
transform 1 0 3956 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1680363874
transform 1 0 3980 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2184
timestamp 1680363874
transform 1 0 4004 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1861
timestamp 1680363874
transform 1 0 4028 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1680363874
transform 1 0 4084 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1680363874
transform 1 0 4076 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2185
timestamp 1680363874
transform 1 0 4060 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1680363874
transform 1 0 4076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1680363874
transform 1 0 4084 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1680363874
transform 1 0 4044 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1680363874
transform 1 0 4052 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1680363874
transform 1 0 4068 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2000
timestamp 1680363874
transform 1 0 4060 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1680363874
transform 1 0 4052 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1680363874
transform 1 0 4100 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2291
timestamp 1680363874
transform 1 0 4092 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1914
timestamp 1680363874
transform 1 0 4172 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1680363874
transform 1 0 4252 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2188
timestamp 1680363874
transform 1 0 4164 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1938
timestamp 1680363874
transform 1 0 4172 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2189
timestamp 1680363874
transform 1 0 4252 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1680363874
transform 1 0 4156 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1965
timestamp 1680363874
transform 1 0 4164 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1680363874
transform 1 0 4156 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1680363874
transform 1 0 4188 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2293
timestamp 1680363874
transform 1 0 4204 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1967
timestamp 1680363874
transform 1 0 4220 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1680363874
transform 1 0 4252 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1680363874
transform 1 0 4252 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2190
timestamp 1680363874
transform 1 0 4276 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1680363874
transform 1 0 4276 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2003
timestamp 1680363874
transform 1 0 4276 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2191
timestamp 1680363874
transform 1 0 4308 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1680363874
transform 1 0 4332 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2040
timestamp 1680363874
transform 1 0 4332 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2192
timestamp 1680363874
transform 1 0 4348 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1939
timestamp 1680363874
transform 1 0 4356 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2193
timestamp 1680363874
transform 1 0 4364 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_2032
timestamp 1680363874
transform 1 0 4364 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1680363874
transform 1 0 4388 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2194
timestamp 1680363874
transform 1 0 4396 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1680363874
transform 1 0 4404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1680363874
transform 1 0 4412 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1680363874
transform 1 0 4388 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1969
timestamp 1680363874
transform 1 0 4396 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1680363874
transform 1 0 4380 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1680363874
transform 1 0 4412 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2297
timestamp 1680363874
transform 1 0 4420 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1680363874
transform 1 0 4444 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2298
timestamp 1680363874
transform 1 0 4476 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2004
timestamp 1680363874
transform 1 0 4468 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1680363874
transform 1 0 4492 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1680363874
transform 1 0 4532 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2197
timestamp 1680363874
transform 1 0 4492 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1680363874
transform 1 0 4508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1680363874
transform 1 0 4524 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1680363874
transform 1 0 4532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1680363874
transform 1 0 4500 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1680363874
transform 1 0 4516 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1971
timestamp 1680363874
transform 1 0 4524 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2301
timestamp 1680363874
transform 1 0 4532 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2005
timestamp 1680363874
transform 1 0 4532 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2201
timestamp 1680363874
transform 1 0 4548 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1680363874
transform 1 0 4572 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1680363874
transform 1 0 4580 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1941
timestamp 1680363874
transform 1 0 4588 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2302
timestamp 1680363874
transform 1 0 4564 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1680363874
transform 1 0 4588 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1680363874
transform 1 0 4596 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2006
timestamp 1680363874
transform 1 0 4588 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1680363874
transform 1 0 4548 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1680363874
transform 1 0 4572 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1680363874
transform 1 0 4604 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2305
timestamp 1680363874
transform 1 0 4620 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_2041
timestamp 1680363874
transform 1 0 4620 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2204
timestamp 1680363874
transform 1 0 4660 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1680363874
transform 1 0 4652 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1972
timestamp 1680363874
transform 1 0 4660 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1680363874
transform 1 0 4684 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1680363874
transform 1 0 4684 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1680363874
transform 1 0 4700 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2205
timestamp 1680363874
transform 1 0 4692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1680363874
transform 1 0 4700 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1680363874
transform 1 0 4684 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1680363874
transform 1 0 4700 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1973
timestamp 1680363874
transform 1 0 4708 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1680363874
transform 1 0 4700 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1680363874
transform 1 0 4684 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1680363874
transform 1 0 4716 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1680363874
transform 1 0 4748 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2207
timestamp 1680363874
transform 1 0 4748 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1680363874
transform 1 0 4748 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1680363874
transform 1 0 4764 0 1 3725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_20
timestamp 1680363874
transform 1 0 24 0 1 3670
box -10 -3 10 3
use FILL  FILL_1581
timestamp 1680363874
transform 1 0 72 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1680363874
transform 1 0 80 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1680363874
transform 1 0 88 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1680363874
transform 1 0 96 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1680363874
transform 1 0 104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1680363874
transform 1 0 112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1680363874
transform 1 0 120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1680363874
transform 1 0 128 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1680363874
transform 1 0 136 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_141
timestamp 1680363874
transform 1 0 144 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1590
timestamp 1680363874
transform 1 0 160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1680363874
transform 1 0 168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1680363874
transform 1 0 176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1680363874
transform 1 0 184 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_115
timestamp 1680363874
transform 1 0 192 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_142
timestamp 1680363874
transform -1 0 248 0 -1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_116
timestamp 1680363874
transform 1 0 248 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1603
timestamp 1680363874
transform 1 0 288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1680363874
transform 1 0 296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1680363874
transform 1 0 304 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_117
timestamp 1680363874
transform 1 0 312 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1606
timestamp 1680363874
transform 1 0 352 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_143
timestamp 1680363874
transform -1 0 376 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1607
timestamp 1680363874
transform 1 0 376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1680363874
transform 1 0 384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1680363874
transform 1 0 392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1680363874
transform 1 0 400 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_144
timestamp 1680363874
transform 1 0 408 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1614
timestamp 1680363874
transform 1 0 504 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_144
timestamp 1680363874
transform 1 0 512 0 -1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_119
timestamp 1680363874
transform 1 0 528 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1618
timestamp 1680363874
transform 1 0 568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1680363874
transform 1 0 576 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1680363874
transform 1 0 584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1680363874
transform 1 0 592 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_121
timestamp 1680363874
transform -1 0 640 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1626
timestamp 1680363874
transform 1 0 640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1680363874
transform 1 0 648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1680363874
transform 1 0 656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1680363874
transform 1 0 664 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1680363874
transform 1 0 672 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_123
timestamp 1680363874
transform 1 0 680 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1635
timestamp 1680363874
transform 1 0 720 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1680363874
transform 1 0 728 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1680363874
transform 1 0 736 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1680363874
transform 1 0 744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1680363874
transform 1 0 752 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_124
timestamp 1680363874
transform -1 0 800 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1645
timestamp 1680363874
transform 1 0 800 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1680363874
transform 1 0 808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1680363874
transform 1 0 816 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1680363874
transform 1 0 824 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1680363874
transform 1 0 832 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1653
timestamp 1680363874
transform 1 0 864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1680363874
transform 1 0 872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1680363874
transform 1 0 880 0 -1 3770
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1680363874
transform 1 0 888 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1661
timestamp 1680363874
transform 1 0 912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1680363874
transform 1 0 920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1680363874
transform 1 0 928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1680363874
transform 1 0 936 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_33
timestamp 1680363874
transform 1 0 944 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1667
timestamp 1680363874
transform 1 0 976 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1680363874
transform 1 0 984 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1680363874
transform 1 0 992 0 -1 3770
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1680363874
transform 1 0 1000 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1673
timestamp 1680363874
transform 1 0 1024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1680363874
transform 1 0 1032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1680363874
transform 1 0 1040 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_126
timestamp 1680363874
transform -1 0 1088 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1679
timestamp 1680363874
transform 1 0 1088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1680363874
transform 1 0 1096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1680363874
transform 1 0 1104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1680363874
transform 1 0 1112 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_129
timestamp 1680363874
transform 1 0 1120 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1687
timestamp 1680363874
transform 1 0 1160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1680363874
transform 1 0 1168 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_146
timestamp 1680363874
transform -1 0 1192 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1689
timestamp 1680363874
transform 1 0 1192 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1680363874
transform 1 0 1200 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1680363874
transform 1 0 1208 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_146
timestamp 1680363874
transform -1 0 1312 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1694
timestamp 1680363874
transform 1 0 1312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1680363874
transform 1 0 1320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1680363874
transform 1 0 1328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1680363874
transform 1 0 1336 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_130
timestamp 1680363874
transform 1 0 1344 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1721
timestamp 1680363874
transform 1 0 1384 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_151
timestamp 1680363874
transform -1 0 1408 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1722
timestamp 1680363874
transform 1 0 1408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1680363874
transform 1 0 1416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1680363874
transform 1 0 1424 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_154
timestamp 1680363874
transform -1 0 1528 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1725
timestamp 1680363874
transform 1 0 1528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1680363874
transform 1 0 1536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1680363874
transform 1 0 1544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1680363874
transform 1 0 1552 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1680363874
transform 1 0 1560 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1680363874
transform 1 0 1584 0 -1 3770
box -8 -3 32 105
use OAI21X1  OAI21X1_34
timestamp 1680363874
transform -1 0 1640 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1680363874
transform -1 0 1672 0 -1 3770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1680363874
transform -1 0 1768 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_152
timestamp 1680363874
transform -1 0 1784 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1729
timestamp 1680363874
transform 1 0 1784 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1680363874
transform 1 0 1792 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1680363874
transform 1 0 1800 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1680363874
transform 1 0 1808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1680363874
transform 1 0 1816 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_89
timestamp 1680363874
transform -1 0 1864 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1734
timestamp 1680363874
transform 1 0 1864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1680363874
transform 1 0 1872 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_90
timestamp 1680363874
transform -1 0 1920 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1736
timestamp 1680363874
transform 1 0 1920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1680363874
transform 1 0 1928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1680363874
transform 1 0 1936 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1680363874
transform 1 0 1944 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1680363874
transform 1 0 1952 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_153
timestamp 1680363874
transform 1 0 1960 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1741
timestamp 1680363874
transform 1 0 1976 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1680363874
transform 1 0 1984 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1680363874
transform 1 0 1992 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1680363874
transform 1 0 2000 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1680363874
transform 1 0 2008 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1680363874
transform 1 0 2016 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1746
timestamp 1680363874
transform 1 0 2040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1680363874
transform 1 0 2048 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1680363874
transform 1 0 2056 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_36
timestamp 1680363874
transform -1 0 2096 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1749
timestamp 1680363874
transform 1 0 2096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1680363874
transform 1 0 2104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1680363874
transform 1 0 2112 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_2043
timestamp 1680363874
transform 1 0 2140 0 1 3675
box -3 -3 3 3
use OAI21X1  OAI21X1_37
timestamp 1680363874
transform -1 0 2152 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1752
timestamp 1680363874
transform 1 0 2152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1680363874
transform 1 0 2160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1680363874
transform 1 0 2168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1680363874
transform 1 0 2176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1680363874
transform 1 0 2184 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1680363874
transform -1 0 2216 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1757
timestamp 1680363874
transform 1 0 2216 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1680363874
transform 1 0 2224 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1680363874
transform 1 0 2232 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_38
timestamp 1680363874
transform -1 0 2272 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1760
timestamp 1680363874
transform 1 0 2272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1680363874
transform 1 0 2280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1680363874
transform 1 0 2288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1680363874
transform 1 0 2296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1680363874
transform 1 0 2304 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1680363874
transform -1 0 2336 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1784
timestamp 1680363874
transform 1 0 2336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1680363874
transform 1 0 2344 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_39
timestamp 1680363874
transform -1 0 2384 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1786
timestamp 1680363874
transform 1 0 2384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1680363874
transform 1 0 2392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1680363874
transform 1 0 2400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1680363874
transform 1 0 2408 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1680363874
transform -1 0 2448 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1790
timestamp 1680363874
transform 1 0 2448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1680363874
transform 1 0 2456 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_159
timestamp 1680363874
transform 1 0 2464 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1792
timestamp 1680363874
transform 1 0 2560 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_92
timestamp 1680363874
transform -1 0 2608 0 -1 3770
box -8 -3 46 105
use NOR2X1  NOR2X1_11
timestamp 1680363874
transform -1 0 2632 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1793
timestamp 1680363874
transform 1 0 2632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1680363874
transform 1 0 2640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1680363874
transform 1 0 2648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1680363874
transform 1 0 2656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1680363874
transform 1 0 2664 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1680363874
transform 1 0 2672 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1680363874
transform 1 0 2680 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1680363874
transform 1 0 2688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1680363874
transform 1 0 2696 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1680363874
transform 1 0 2704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1680363874
transform 1 0 2712 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1680363874
transform 1 0 2720 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1680363874
transform 1 0 2728 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1680363874
transform 1 0 2736 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1680363874
transform 1 0 2744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1680363874
transform 1 0 2752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1680363874
transform 1 0 2760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1680363874
transform 1 0 2768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1680363874
transform 1 0 2776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1680363874
transform 1 0 2784 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1680363874
transform 1 0 2792 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_161
timestamp 1680363874
transform 1 0 2888 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1813
timestamp 1680363874
transform 1 0 2984 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1680363874
transform 1 0 2992 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_41
timestamp 1680363874
transform 1 0 3000 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1818
timestamp 1680363874
transform 1 0 3032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1680363874
transform 1 0 3040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1680363874
transform 1 0 3048 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1680363874
transform 1 0 3056 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_2044
timestamp 1680363874
transform 1 0 3092 0 1 3675
box -3 -3 3 3
use OAI21X1  OAI21X1_43
timestamp 1680363874
transform -1 0 3096 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1831
timestamp 1680363874
transform 1 0 3096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1680363874
transform 1 0 3104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1680363874
transform 1 0 3112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1680363874
transform 1 0 3120 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1680363874
transform -1 0 3152 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1835
timestamp 1680363874
transform 1 0 3152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1680363874
transform 1 0 3160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1680363874
transform 1 0 3168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1680363874
transform 1 0 3176 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1680363874
transform -1 0 3280 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1839
timestamp 1680363874
transform 1 0 3280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1680363874
transform 1 0 3288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1680363874
transform 1 0 3296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1680363874
transform 1 0 3304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1680363874
transform 1 0 3312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1680363874
transform 1 0 3320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1680363874
transform 1 0 3328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1680363874
transform 1 0 3336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1680363874
transform 1 0 3344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1680363874
transform 1 0 3352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1680363874
transform 1 0 3360 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_2045
timestamp 1680363874
transform 1 0 3380 0 1 3675
box -3 -3 3 3
use FILL  FILL_1873
timestamp 1680363874
transform 1 0 3368 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_2046
timestamp 1680363874
transform 1 0 3396 0 1 3675
box -3 -3 3 3
use OAI21X1  OAI21X1_45
timestamp 1680363874
transform -1 0 3408 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1874
timestamp 1680363874
transform 1 0 3408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1680363874
transform 1 0 3416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1680363874
transform 1 0 3424 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1680363874
transform 1 0 3432 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1680363874
transform 1 0 3440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1680363874
transform 1 0 3448 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1680363874
transform -1 0 3480 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1880
timestamp 1680363874
transform 1 0 3480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1680363874
transform 1 0 3488 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1680363874
transform 1 0 3496 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1680363874
transform 1 0 3504 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1680363874
transform -1 0 3608 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1884
timestamp 1680363874
transform 1 0 3608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1680363874
transform 1 0 3616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1680363874
transform 1 0 3624 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1680363874
transform 1 0 3632 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_46
timestamp 1680363874
transform 1 0 3640 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1888
timestamp 1680363874
transform 1 0 3672 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1680363874
transform 1 0 3680 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1680363874
transform 1 0 3688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1680363874
transform 1 0 3696 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1680363874
transform 1 0 3704 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_96
timestamp 1680363874
transform 1 0 3712 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1898
timestamp 1680363874
transform 1 0 3752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1680363874
transform 1 0 3760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1680363874
transform 1 0 3768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1680363874
transform 1 0 3776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1680363874
transform 1 0 3784 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1680363874
transform 1 0 3792 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_167
timestamp 1680363874
transform -1 0 3896 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1909
timestamp 1680363874
transform 1 0 3896 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1680363874
transform 1 0 3904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1680363874
transform 1 0 3912 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_97
timestamp 1680363874
transform 1 0 3920 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1914
timestamp 1680363874
transform 1 0 3960 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1680363874
transform 1 0 3968 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1680363874
transform 1 0 3976 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_160
timestamp 1680363874
transform 1 0 3984 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1921
timestamp 1680363874
transform 1 0 4000 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1680363874
transform 1 0 4008 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1680363874
transform 1 0 4016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1680363874
transform 1 0 4024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1680363874
transform 1 0 4032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1680363874
transform 1 0 4040 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_98
timestamp 1680363874
transform -1 0 4088 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1927
timestamp 1680363874
transform 1 0 4088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1680363874
transform 1 0 4096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1680363874
transform 1 0 4104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1680363874
transform 1 0 4112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1680363874
transform 1 0 4120 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_162
timestamp 1680363874
transform -1 0 4144 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1950
timestamp 1680363874
transform 1 0 4144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1680363874
transform 1 0 4152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1680363874
transform 1 0 4160 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1680363874
transform -1 0 4264 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1953
timestamp 1680363874
transform 1 0 4264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1680363874
transform 1 0 4272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1680363874
transform 1 0 4280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1680363874
transform 1 0 4288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1680363874
transform 1 0 4296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1680363874
transform 1 0 4304 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_163
timestamp 1680363874
transform -1 0 4328 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1961
timestamp 1680363874
transform 1 0 4328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1680363874
transform 1 0 4336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1680363874
transform 1 0 4344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1680363874
transform 1 0 4352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1680363874
transform 1 0 4360 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_99
timestamp 1680363874
transform -1 0 4408 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1969
timestamp 1680363874
transform 1 0 4408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1680363874
transform 1 0 4416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1680363874
transform 1 0 4424 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_164
timestamp 1680363874
transform 1 0 4432 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1972
timestamp 1680363874
transform 1 0 4448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1680363874
transform 1 0 4456 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1680363874
transform 1 0 4464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1680363874
transform 1 0 4472 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1680363874
transform 1 0 4480 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_138
timestamp 1680363874
transform 1 0 4488 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1981
timestamp 1680363874
transform 1 0 4528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1680363874
transform 1 0 4536 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_100
timestamp 1680363874
transform -1 0 4584 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_166
timestamp 1680363874
transform 1 0 4584 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1983
timestamp 1680363874
transform 1 0 4600 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1680363874
transform 1 0 4608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1680363874
transform 1 0 4616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1680363874
transform 1 0 4624 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1680363874
transform 1 0 4632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1680363874
transform 1 0 4640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1680363874
transform 1 0 4648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1680363874
transform 1 0 4656 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_102
timestamp 1680363874
transform -1 0 4704 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1993
timestamp 1680363874
transform 1 0 4704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1680363874
transform 1 0 4712 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1680363874
transform 1 0 4720 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_167
timestamp 1680363874
transform 1 0 4728 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1996
timestamp 1680363874
transform 1 0 4744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1680363874
transform 1 0 4752 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_168
timestamp 1680363874
transform 1 0 4760 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1998
timestamp 1680363874
transform 1 0 4776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1680363874
transform 1 0 4784 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1680363874
transform 1 0 4792 0 -1 3770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_21
timestamp 1680363874
transform 1 0 4851 0 1 3670
box -10 -3 10 3
use M3_M2  M3_M2_2088
timestamp 1680363874
transform 1 0 132 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2343
timestamp 1680363874
transform 1 0 132 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1680363874
transform 1 0 84 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2072
timestamp 1680363874
transform 1 0 204 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2344
timestamp 1680363874
transform 1 0 204 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1680363874
transform 1 0 204 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1680363874
transform 1 0 220 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1680363874
transform 1 0 228 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2056
timestamp 1680363874
transform 1 0 260 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1680363874
transform 1 0 276 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1680363874
transform 1 0 244 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1680363874
transform 1 0 268 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2346
timestamp 1680363874
transform 1 0 292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1680363874
transform 1 0 244 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2180
timestamp 1680363874
transform 1 0 292 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1680363874
transform 1 0 244 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1680363874
transform 1 0 380 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2347
timestamp 1680363874
transform 1 0 380 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1680363874
transform 1 0 444 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1680363874
transform 1 0 396 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2157
timestamp 1680363874
transform 1 0 444 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1680363874
transform 1 0 396 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1680363874
transform 1 0 484 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1680363874
transform 1 0 524 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1680363874
transform 1 0 516 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2349
timestamp 1680363874
transform 1 0 508 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1680363874
transform 1 0 516 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1680363874
transform 1 0 500 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1680363874
transform 1 0 548 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1680363874
transform 1 0 540 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2159
timestamp 1680363874
transform 1 0 548 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2452
timestamp 1680363874
transform 1 0 556 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2181
timestamp 1680363874
transform 1 0 540 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1680363874
transform 1 0 620 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1680363874
transform 1 0 636 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2453
timestamp 1680363874
transform 1 0 636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2219
timestamp 1680363874
transform 1 0 636 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1680363874
transform 1 0 684 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2352
timestamp 1680363874
transform 1 0 668 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1680363874
transform 1 0 684 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1680363874
transform 1 0 676 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1680363874
transform 1 0 692 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1680363874
transform 1 0 700 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2182
timestamp 1680363874
transform 1 0 676 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1680363874
transform 1 0 684 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1680363874
transform 1 0 716 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1680363874
transform 1 0 708 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2354
timestamp 1680363874
transform 1 0 724 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2059
timestamp 1680363874
transform 1 0 748 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1680363874
transform 1 0 740 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2326
timestamp 1680363874
transform 1 0 748 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2060
timestamp 1680363874
transform 1 0 764 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1680363874
transform 1 0 772 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2355
timestamp 1680363874
transform 1 0 764 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2076
timestamp 1680363874
transform 1 0 788 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2457
timestamp 1680363874
transform 1 0 796 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2183
timestamp 1680363874
transform 1 0 820 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2458
timestamp 1680363874
transform 1 0 836 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2184
timestamp 1680363874
transform 1 0 836 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1680363874
transform 1 0 860 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2327
timestamp 1680363874
transform 1 0 868 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1680363874
transform 1 0 852 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1680363874
transform 1 0 860 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2185
timestamp 1680363874
transform 1 0 860 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1680363874
transform 1 0 892 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2328
timestamp 1680363874
transform 1 0 892 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2096
timestamp 1680363874
transform 1 0 900 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1680363874
transform 1 0 924 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2460
timestamp 1680363874
transform 1 0 924 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2078
timestamp 1680363874
transform 1 0 972 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2357
timestamp 1680363874
transform 1 0 956 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1680363874
transform 1 0 964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1680363874
transform 1 0 972 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1680363874
transform 1 0 964 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2186
timestamp 1680363874
transform 1 0 956 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1680363874
transform 1 0 964 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1680363874
transform 1 0 980 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2360
timestamp 1680363874
transform 1 0 988 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2097
timestamp 1680363874
transform 1 0 1028 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1680363874
transform 1 0 1004 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2361
timestamp 1680363874
transform 1 0 1028 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2131
timestamp 1680363874
transform 1 0 1044 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2462
timestamp 1680363874
transform 1 0 1004 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1680363874
transform 1 0 1020 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1680363874
transform 1 0 1036 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1680363874
transform 1 0 1044 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2223
timestamp 1680363874
transform 1 0 996 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1680363874
transform 1 0 1020 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1680363874
transform 1 0 1036 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1680363874
transform 1 0 1060 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2362
timestamp 1680363874
transform 1 0 1060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1680363874
transform 1 0 1084 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1680363874
transform 1 0 1100 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2161
timestamp 1680363874
transform 1 0 1076 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2466
timestamp 1680363874
transform 1 0 1092 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2162
timestamp 1680363874
transform 1 0 1100 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2467
timestamp 1680363874
transform 1 0 1108 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2189
timestamp 1680363874
transform 1 0 1108 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1680363874
transform 1 0 1108 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1680363874
transform 1 0 1132 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2365
timestamp 1680363874
transform 1 0 1124 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2163
timestamp 1680363874
transform 1 0 1148 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1680363874
transform 1 0 1180 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2366
timestamp 1680363874
transform 1 0 1180 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2132
timestamp 1680363874
transform 1 0 1188 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2367
timestamp 1680363874
transform 1 0 1196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1680363874
transform 1 0 1156 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1680363874
transform 1 0 1172 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1680363874
transform 1 0 1204 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2133
timestamp 1680363874
transform 1 0 1228 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1680363874
transform 1 0 1260 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2368
timestamp 1680363874
transform 1 0 1244 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1680363874
transform 1 0 1260 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2134
timestamp 1680363874
transform 1 0 1268 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2471
timestamp 1680363874
transform 1 0 1228 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1680363874
transform 1 0 1236 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1680363874
transform 1 0 1252 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1680363874
transform 1 0 1268 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2225
timestamp 1680363874
transform 1 0 1244 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1680363874
transform 1 0 1324 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2370
timestamp 1680363874
transform 1 0 1324 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1680363874
transform 1 0 1340 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1680363874
transform 1 0 1316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1680363874
transform 1 0 1332 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2164
timestamp 1680363874
transform 1 0 1340 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2477
timestamp 1680363874
transform 1 0 1348 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2190
timestamp 1680363874
transform 1 0 1332 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1680363874
transform 1 0 1356 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1680363874
transform 1 0 1372 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1680363874
transform 1 0 1412 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1680363874
transform 1 0 1412 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2372
timestamp 1680363874
transform 1 0 1388 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1680363874
transform 1 0 1412 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1680363874
transform 1 0 1428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1680363874
transform 1 0 1388 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1680363874
transform 1 0 1404 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1680363874
transform 1 0 1420 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1680363874
transform 1 0 1388 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1680363874
transform 1 0 1412 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1680363874
transform 1 0 1428 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2375
timestamp 1680363874
transform 1 0 1524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1680363874
transform 1 0 1572 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2191
timestamp 1680363874
transform 1 0 1524 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1680363874
transform 1 0 1588 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2482
timestamp 1680363874
transform 1 0 1588 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2137
timestamp 1680363874
transform 1 0 1612 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2376
timestamp 1680363874
transform 1 0 1620 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2138
timestamp 1680363874
transform 1 0 1636 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2483
timestamp 1680363874
transform 1 0 1636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2192
timestamp 1680363874
transform 1 0 1636 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2329
timestamp 1680363874
transform 1 0 1660 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2193
timestamp 1680363874
transform 1 0 1652 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2484
timestamp 1680363874
transform 1 0 1700 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1680363874
transform 1 0 1708 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_2079
timestamp 1680363874
transform 1 0 1740 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2330
timestamp 1680363874
transform 1 0 1748 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1680363874
transform 1 0 1788 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1680363874
transform 1 0 1804 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2101
timestamp 1680363874
transform 1 0 1820 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2377
timestamp 1680363874
transform 1 0 1820 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1680363874
transform 1 0 1828 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1680363874
transform 1 0 1852 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1680363874
transform 1 0 1844 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1680363874
transform 1 0 1844 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_2229
timestamp 1680363874
transform 1 0 1844 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1680363874
transform 1 0 1884 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2379
timestamp 1680363874
transform 1 0 1884 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1680363874
transform 1 0 1892 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2230
timestamp 1680363874
transform 1 0 1876 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1680363874
transform 1 0 1996 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1680363874
transform 1 0 1964 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2381
timestamp 1680363874
transform 1 0 1972 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2140
timestamp 1680363874
transform 1 0 1996 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2488
timestamp 1680363874
transform 1 0 1996 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2194
timestamp 1680363874
transform 1 0 1932 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2489
timestamp 1680363874
transform 1 0 2020 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1680363874
transform 1 0 2012 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1680363874
transform 1 0 2044 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2195
timestamp 1680363874
transform 1 0 2044 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1680363874
transform 1 0 2100 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2382
timestamp 1680363874
transform 1 0 2108 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1680363874
transform 1 0 2116 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2103
timestamp 1680363874
transform 1 0 2132 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2490
timestamp 1680363874
transform 1 0 2132 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1680363874
transform 1 0 2140 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1680363874
transform 1 0 2148 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2104
timestamp 1680363874
transform 1 0 2164 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1680363874
transform 1 0 2164 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2384
timestamp 1680363874
transform 1 0 2196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1680363874
transform 1 0 2188 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1680363874
transform 1 0 2220 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2142
timestamp 1680363874
transform 1 0 2220 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2493
timestamp 1680363874
transform 1 0 2212 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1680363874
transform 1 0 2228 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1680363874
transform 1 0 2260 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2231
timestamp 1680363874
transform 1 0 2260 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2386
timestamp 1680363874
transform 1 0 2292 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2166
timestamp 1680363874
transform 1 0 2292 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1680363874
transform 1 0 2308 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2494
timestamp 1680363874
transform 1 0 2308 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1680363874
transform 1 0 2316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1680363874
transform 1 0 2340 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2196
timestamp 1680363874
transform 1 0 2340 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1680363874
transform 1 0 2356 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2387
timestamp 1680363874
transform 1 0 2356 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2167
timestamp 1680363874
transform 1 0 2356 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1680363874
transform 1 0 2380 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1680363874
transform 1 0 2372 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2496
timestamp 1680363874
transform 1 0 2380 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2106
timestamp 1680363874
transform 1 0 2404 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2335
timestamp 1680363874
transform 1 0 2420 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1680363874
transform 1 0 2396 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2197
timestamp 1680363874
transform 1 0 2420 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1680363874
transform 1 0 2436 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1680363874
transform 1 0 2460 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2388
timestamp 1680363874
transform 1 0 2468 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1680363874
transform 1 0 2460 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1680363874
transform 1 0 2492 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2146
timestamp 1680363874
transform 1 0 2492 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2499
timestamp 1680363874
transform 1 0 2476 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1680363874
transform 1 0 2484 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2168
timestamp 1680363874
transform 1 0 2492 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2549
timestamp 1680363874
transform 1 0 2500 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_2048
timestamp 1680363874
transform 1 0 2532 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2389
timestamp 1680363874
transform 1 0 2532 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1680363874
transform 1 0 2540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1680363874
transform 1 0 2540 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2064
timestamp 1680363874
transform 1 0 2564 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2337
timestamp 1680363874
transform 1 0 2564 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2198
timestamp 1680363874
transform 1 0 2540 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1680363874
transform 1 0 2556 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1680363874
transform 1 0 2588 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2502
timestamp 1680363874
transform 1 0 2580 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1680363874
transform 1 0 2588 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2108
timestamp 1680363874
transform 1 0 2612 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2391
timestamp 1680363874
transform 1 0 2612 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2232
timestamp 1680363874
transform 1 0 2612 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2392
timestamp 1680363874
transform 1 0 2644 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1680363874
transform 1 0 2652 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1680363874
transform 1 0 2636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2169
timestamp 1680363874
transform 1 0 2660 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1680363874
transform 1 0 2700 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2394
timestamp 1680363874
transform 1 0 2676 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1680363874
transform 1 0 2700 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1680363874
transform 1 0 2692 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1680363874
transform 1 0 2708 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1680363874
transform 1 0 2716 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2110
timestamp 1680363874
transform 1 0 2724 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2396
timestamp 1680363874
transform 1 0 2724 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2053
timestamp 1680363874
transform 1 0 2820 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2338
timestamp 1680363874
transform 1 0 2844 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2111
timestamp 1680363874
transform 1 0 2868 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2397
timestamp 1680363874
transform 1 0 2868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1680363874
transform 1 0 2884 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1680363874
transform 1 0 2908 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1680363874
transform 1 0 2940 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1680363874
transform 1 0 2956 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2398
timestamp 1680363874
transform 1 0 2940 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2055
timestamp 1680363874
transform 1 0 2972 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1680363874
transform 1 0 2972 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2339
timestamp 1680363874
transform 1 0 2964 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2147
timestamp 1680363874
transform 1 0 2964 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2399
timestamp 1680363874
transform 1 0 2972 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1680363874
transform 1 0 2964 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2112
timestamp 1680363874
transform 1 0 2988 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1680363874
transform 1 0 3012 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2400
timestamp 1680363874
transform 1 0 2996 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2170
timestamp 1680363874
transform 1 0 2996 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1680363874
transform 1 0 3020 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2148
timestamp 1680363874
transform 1 0 3020 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1680363874
transform 1 0 3044 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2401
timestamp 1680363874
transform 1 0 3052 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1680363874
transform 1 0 3036 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1680363874
transform 1 0 3044 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2171
timestamp 1680363874
transform 1 0 3052 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2341
timestamp 1680363874
transform 1 0 3076 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2150
timestamp 1680363874
transform 1 0 3076 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1680363874
transform 1 0 3100 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1680363874
transform 1 0 3092 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1680363874
transform 1 0 3132 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2402
timestamp 1680363874
transform 1 0 3132 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1680363874
transform 1 0 3116 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2172
timestamp 1680363874
transform 1 0 3132 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1680363874
transform 1 0 3116 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1680363874
transform 1 0 3148 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2513
timestamp 1680363874
transform 1 0 3148 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1680363874
transform 1 0 3164 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1680363874
transform 1 0 3188 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1680363874
transform 1 0 3196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1680363874
transform 1 0 3188 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1680363874
transform 1 0 3204 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1680363874
transform 1 0 3236 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2404
timestamp 1680363874
transform 1 0 3244 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1680363874
transform 1 0 3228 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1680363874
transform 1 0 3260 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1680363874
transform 1 0 3284 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1680363874
transform 1 0 3316 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2405
timestamp 1680363874
transform 1 0 3268 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1680363874
transform 1 0 3276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1680363874
transform 1 0 3292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1680363874
transform 1 0 3308 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1680363874
transform 1 0 3316 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2174
timestamp 1680363874
transform 1 0 3268 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2515
timestamp 1680363874
transform 1 0 3276 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1680363874
transform 1 0 3284 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1680363874
transform 1 0 3300 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2235
timestamp 1680363874
transform 1 0 3276 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1680363874
transform 1 0 3348 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2518
timestamp 1680363874
transform 1 0 3340 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2202
timestamp 1680363874
transform 1 0 3340 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1680363874
transform 1 0 3332 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2410
timestamp 1680363874
transform 1 0 3364 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2175
timestamp 1680363874
transform 1 0 3364 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1680363874
transform 1 0 3364 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1680363874
transform 1 0 3396 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2411
timestamp 1680363874
transform 1 0 3404 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1680363874
transform 1 0 3428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1680363874
transform 1 0 3388 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1680363874
transform 1 0 3396 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1680363874
transform 1 0 3412 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1680363874
transform 1 0 3420 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2238
timestamp 1680363874
transform 1 0 3380 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1680363874
transform 1 0 3412 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1680363874
transform 1 0 3412 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1680363874
transform 1 0 3428 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2523
timestamp 1680363874
transform 1 0 3476 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2204
timestamp 1680363874
transform 1 0 3476 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2413
timestamp 1680363874
transform 1 0 3492 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1680363874
transform 1 0 3516 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2205
timestamp 1680363874
transform 1 0 3516 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2415
timestamp 1680363874
transform 1 0 3620 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2177
timestamp 1680363874
transform 1 0 3620 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2416
timestamp 1680363874
transform 1 0 3660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1680363874
transform 1 0 3636 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1680363874
transform 1 0 3652 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2240
timestamp 1680363874
transform 1 0 3660 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1680363874
transform 1 0 3676 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1680363874
transform 1 0 3716 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2417
timestamp 1680363874
transform 1 0 3732 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1680363874
transform 1 0 3740 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2342
timestamp 1680363874
transform 1 0 3756 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2115
timestamp 1680363874
transform 1 0 3844 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2418
timestamp 1680363874
transform 1 0 3820 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1680363874
transform 1 0 3828 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1680363874
transform 1 0 3844 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1680363874
transform 1 0 3812 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1680363874
transform 1 0 3868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1680363874
transform 1 0 3860 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2207
timestamp 1680363874
transform 1 0 3860 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1680363874
transform 1 0 3884 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1680363874
transform 1 0 3892 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2528
timestamp 1680363874
transform 1 0 3892 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2070
timestamp 1680363874
transform 1 0 3964 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1680363874
transform 1 0 3980 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1680363874
transform 1 0 3924 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1680363874
transform 1 0 3908 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1680363874
transform 1 0 3948 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2422
timestamp 1680363874
transform 1 0 3908 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1680363874
transform 1 0 3916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1680363874
transform 1 0 3948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1680363874
transform 1 0 3996 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2208
timestamp 1680363874
transform 1 0 3916 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1680363874
transform 1 0 3972 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1680363874
transform 1 0 3996 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2425
timestamp 1680363874
transform 1 0 4092 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1680363874
transform 1 0 4044 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2211
timestamp 1680363874
transform 1 0 4044 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1680363874
transform 1 0 4060 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2531
timestamp 1680363874
transform 1 0 4132 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2119
timestamp 1680363874
transform 1 0 4204 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1680363874
transform 1 0 4292 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2426
timestamp 1680363874
transform 1 0 4164 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1680363874
transform 1 0 4172 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1680363874
transform 1 0 4188 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1680363874
transform 1 0 4204 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1680363874
transform 1 0 4252 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2212
timestamp 1680363874
transform 1 0 4164 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2532
timestamp 1680363874
transform 1 0 4196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2213
timestamp 1680363874
transform 1 0 4196 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2533
timestamp 1680363874
transform 1 0 4220 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2085
timestamp 1680363874
transform 1 0 4372 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1680363874
transform 1 0 4372 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2431
timestamp 1680363874
transform 1 0 4332 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1680363874
transform 1 0 4348 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1680363874
transform 1 0 4364 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1680363874
transform 1 0 4372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1680363874
transform 1 0 4340 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1680363874
transform 1 0 4356 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2214
timestamp 1680363874
transform 1 0 4396 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1680363874
transform 1 0 4436 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2435
timestamp 1680363874
transform 1 0 4436 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1680363874
transform 1 0 4428 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1680363874
transform 1 0 4444 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2123
timestamp 1680363874
transform 1 0 4468 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1680363874
transform 1 0 4492 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2436
timestamp 1680363874
transform 1 0 4460 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2154
timestamp 1680363874
transform 1 0 4468 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2437
timestamp 1680363874
transform 1 0 4476 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1680363874
transform 1 0 4492 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1680363874
transform 1 0 4492 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2243
timestamp 1680363874
transform 1 0 4484 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1680363874
transform 1 0 4516 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1680363874
transform 1 0 4596 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1680363874
transform 1 0 4556 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1680363874
transform 1 0 4652 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2439
timestamp 1680363874
transform 1 0 4572 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1680363874
transform 1 0 4636 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2156
timestamp 1680363874
transform 1 0 4644 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2441
timestamp 1680363874
transform 1 0 4652 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1680363874
transform 1 0 4620 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1680363874
transform 1 0 4636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2179
timestamp 1680363874
transform 1 0 4652 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2541
timestamp 1680363874
transform 1 0 4660 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2215
timestamp 1680363874
transform 1 0 4636 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1680363874
transform 1 0 4628 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1680363874
transform 1 0 4676 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1680363874
transform 1 0 4676 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2542
timestamp 1680363874
transform 1 0 4676 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2245
timestamp 1680363874
transform 1 0 4668 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2442
timestamp 1680363874
transform 1 0 4684 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1680363874
transform 1 0 4700 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1680363874
transform 1 0 4708 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1680363874
transform 1 0 4748 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2216
timestamp 1680363874
transform 1 0 4692 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2543
timestamp 1680363874
transform 1 0 4788 0 1 3605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_22
timestamp 1680363874
transform 1 0 48 0 1 3570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_173
timestamp 1680363874
transform 1 0 72 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_169
timestamp 1680363874
transform 1 0 168 0 1 3570
box -9 -3 26 105
use FILL  FILL_2001
timestamp 1680363874
transform 1 0 184 0 1 3570
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1680363874
transform 1 0 192 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1680363874
transform 1 0 200 0 1 3570
box -8 -3 32 105
use FILL  FILL_2007
timestamp 1680363874
transform 1 0 224 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1680363874
transform 1 0 232 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_2246
timestamp 1680363874
transform 1 0 348 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_170
timestamp 1680363874
transform 1 0 328 0 1 3570
box -9 -3 26 105
use FILL  FILL_2008
timestamp 1680363874
transform 1 0 344 0 1 3570
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1680363874
transform 1 0 352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1680363874
transform 1 0 360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1680363874
transform 1 0 368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1680363874
transform 1 0 376 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2247
timestamp 1680363874
transform 1 0 404 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_177
timestamp 1680363874
transform 1 0 384 0 1 3570
box -8 -3 104 105
use FILL  FILL_2022
timestamp 1680363874
transform 1 0 480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1680363874
transform 1 0 488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1680363874
transform 1 0 496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1680363874
transform 1 0 504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1680363874
transform 1 0 512 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_141
timestamp 1680363874
transform 1 0 520 0 1 3570
box -8 -3 46 105
use FILL  FILL_2036
timestamp 1680363874
transform 1 0 560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1680363874
transform 1 0 568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1680363874
transform 1 0 576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1680363874
transform 1 0 584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1680363874
transform 1 0 592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1680363874
transform 1 0 600 0 1 3570
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1680363874
transform 1 0 608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1680363874
transform 1 0 616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1680363874
transform 1 0 624 0 1 3570
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1680363874
transform 1 0 632 0 1 3570
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1680363874
transform 1 0 640 0 1 3570
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1680363874
transform 1 0 648 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_143
timestamp 1680363874
transform 1 0 656 0 1 3570
box -8 -3 46 105
use FILL  FILL_2058
timestamp 1680363874
transform 1 0 696 0 1 3570
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1680363874
transform 1 0 704 0 1 3570
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1680363874
transform 1 0 712 0 1 3570
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1680363874
transform 1 0 720 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_9
timestamp 1680363874
transform 1 0 728 0 1 3570
box -8 -3 32 105
use FILL  FILL_2070
timestamp 1680363874
transform 1 0 752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1680363874
transform 1 0 760 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_11
timestamp 1680363874
transform -1 0 792 0 1 3570
box -8 -3 32 105
use FILL  FILL_2074
timestamp 1680363874
transform 1 0 792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1680363874
transform 1 0 800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1680363874
transform 1 0 808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1680363874
transform 1 0 816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1680363874
transform 1 0 824 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_12
timestamp 1680363874
transform 1 0 832 0 1 3570
box -8 -3 32 105
use FILL  FILL_2084
timestamp 1680363874
transform 1 0 856 0 1 3570
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1680363874
transform 1 0 864 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2248
timestamp 1680363874
transform 1 0 884 0 1 3575
box -3 -3 3 3
use FILL  FILL_2091
timestamp 1680363874
transform 1 0 872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1680363874
transform 1 0 880 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_48
timestamp 1680363874
transform -1 0 920 0 1 3570
box -8 -3 34 105
use FILL  FILL_2093
timestamp 1680363874
transform 1 0 920 0 1 3570
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1680363874
transform 1 0 928 0 1 3570
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1680363874
transform 1 0 936 0 1 3570
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1680363874
transform 1 0 944 0 1 3570
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1680363874
transform 1 0 952 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_172
timestamp 1680363874
transform 1 0 960 0 1 3570
box -9 -3 26 105
use FILL  FILL_2102
timestamp 1680363874
transform 1 0 976 0 1 3570
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1680363874
transform 1 0 984 0 1 3570
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1680363874
transform 1 0 992 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_144
timestamp 1680363874
transform 1 0 1000 0 1 3570
box -8 -3 46 105
use FILL  FILL_2105
timestamp 1680363874
transform 1 0 1040 0 1 3570
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1680363874
transform 1 0 1048 0 1 3570
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1680363874
transform 1 0 1056 0 1 3570
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1680363874
transform 1 0 1064 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2249
timestamp 1680363874
transform 1 0 1092 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_146
timestamp 1680363874
transform 1 0 1072 0 1 3570
box -8 -3 46 105
use FILL  FILL_2115
timestamp 1680363874
transform 1 0 1112 0 1 3570
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1680363874
transform 1 0 1120 0 1 3570
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1680363874
transform 1 0 1128 0 1 3570
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1680363874
transform 1 0 1136 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2250
timestamp 1680363874
transform 1 0 1156 0 1 3575
box -3 -3 3 3
use FILL  FILL_2126
timestamp 1680363874
transform 1 0 1144 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2251
timestamp 1680363874
transform 1 0 1180 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_148
timestamp 1680363874
transform 1 0 1152 0 1 3570
box -8 -3 46 105
use FILL  FILL_2128
timestamp 1680363874
transform 1 0 1192 0 1 3570
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1680363874
transform 1 0 1200 0 1 3570
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1680363874
transform 1 0 1208 0 1 3570
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1680363874
transform 1 0 1216 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2252
timestamp 1680363874
transform 1 0 1236 0 1 3575
box -3 -3 3 3
use FILL  FILL_2140
timestamp 1680363874
transform 1 0 1224 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_149
timestamp 1680363874
transform 1 0 1232 0 1 3570
box -8 -3 46 105
use FILL  FILL_2141
timestamp 1680363874
transform 1 0 1272 0 1 3570
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1680363874
transform 1 0 1280 0 1 3570
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1680363874
transform 1 0 1288 0 1 3570
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1680363874
transform 1 0 1296 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2253
timestamp 1680363874
transform 1 0 1316 0 1 3575
box -3 -3 3 3
use FILL  FILL_2145
timestamp 1680363874
transform 1 0 1304 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_150
timestamp 1680363874
transform -1 0 1352 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_2254
timestamp 1680363874
transform 1 0 1364 0 1 3575
box -3 -3 3 3
use FILL  FILL_2146
timestamp 1680363874
transform 1 0 1352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1680363874
transform 1 0 1360 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2255
timestamp 1680363874
transform 1 0 1380 0 1 3575
box -3 -3 3 3
use FILL  FILL_2153
timestamp 1680363874
transform 1 0 1368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1680363874
transform 1 0 1376 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2256
timestamp 1680363874
transform 1 0 1420 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_151
timestamp 1680363874
transform 1 0 1384 0 1 3570
box -8 -3 46 105
use FILL  FILL_2155
timestamp 1680363874
transform 1 0 1424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1680363874
transform 1 0 1432 0 1 3570
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1680363874
transform 1 0 1440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1680363874
transform 1 0 1448 0 1 3570
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1680363874
transform 1 0 1456 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_174
timestamp 1680363874
transform -1 0 1480 0 1 3570
box -9 -3 26 105
use FILL  FILL_2164
timestamp 1680363874
transform 1 0 1480 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1680363874
transform -1 0 1584 0 1 3570
box -8 -3 104 105
use FILL  FILL_2165
timestamp 1680363874
transform 1 0 1584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1680363874
transform 1 0 1592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1680363874
transform 1 0 1600 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_50
timestamp 1680363874
transform 1 0 1608 0 1 3570
box -8 -3 34 105
use FILL  FILL_2175
timestamp 1680363874
transform 1 0 1640 0 1 3570
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1680363874
transform 1 0 1648 0 1 3570
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1680363874
transform 1 0 1656 0 1 3570
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1680363874
transform 1 0 1664 0 1 3570
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1680363874
transform 1 0 1672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1680363874
transform 1 0 1680 0 1 3570
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1680363874
transform 1 0 1688 0 1 3570
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1680363874
transform 1 0 1696 0 1 3570
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1680363874
transform 1 0 1704 0 1 3570
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1680363874
transform 1 0 1712 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_17
timestamp 1680363874
transform 1 0 1720 0 1 3570
box -8 -3 32 105
use FILL  FILL_2191
timestamp 1680363874
transform 1 0 1744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1680363874
transform 1 0 1752 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_53
timestamp 1680363874
transform -1 0 1792 0 1 3570
box -8 -3 34 105
use FILL  FILL_2193
timestamp 1680363874
transform 1 0 1792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1680363874
transform 1 0 1800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1680363874
transform 1 0 1808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1680363874
transform 1 0 1816 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_18
timestamp 1680363874
transform -1 0 1848 0 1 3570
box -8 -3 32 105
use FILL  FILL_2197
timestamp 1680363874
transform 1 0 1848 0 1 3570
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1680363874
transform 1 0 1856 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_56
timestamp 1680363874
transform -1 0 1896 0 1 3570
box -8 -3 34 105
use FILL  FILL_2208
timestamp 1680363874
transform 1 0 1896 0 1 3570
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1680363874
transform 1 0 1904 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1680363874
transform -1 0 2008 0 1 3570
box -8 -3 104 105
use FILL  FILL_2210
timestamp 1680363874
transform 1 0 2008 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_19
timestamp 1680363874
transform 1 0 2016 0 1 3570
box -8 -3 32 105
use FILL  FILL_2223
timestamp 1680363874
transform 1 0 2040 0 1 3570
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1680363874
transform 1 0 2048 0 1 3570
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1680363874
transform 1 0 2056 0 1 3570
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1680363874
transform 1 0 2064 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_60
timestamp 1680363874
transform -1 0 2104 0 1 3570
box -8 -3 34 105
use FILL  FILL_2229
timestamp 1680363874
transform 1 0 2104 0 1 3570
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1680363874
transform 1 0 2112 0 1 3570
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1680363874
transform 1 0 2120 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_20
timestamp 1680363874
transform -1 0 2152 0 1 3570
box -8 -3 32 105
use FILL  FILL_2232
timestamp 1680363874
transform 1 0 2152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1680363874
transform 1 0 2160 0 1 3570
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1680363874
transform 1 0 2168 0 1 3570
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1680363874
transform 1 0 2176 0 1 3570
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1680363874
transform 1 0 2184 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_21
timestamp 1680363874
transform -1 0 2216 0 1 3570
box -8 -3 32 105
use FILL  FILL_2246
timestamp 1680363874
transform 1 0 2216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1680363874
transform 1 0 2224 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2257
timestamp 1680363874
transform 1 0 2252 0 1 3575
box -3 -3 3 3
use OAI21X1  OAI21X1_63
timestamp 1680363874
transform -1 0 2264 0 1 3570
box -8 -3 34 105
use FILL  FILL_2251
timestamp 1680363874
transform 1 0 2264 0 1 3570
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1680363874
transform 1 0 2272 0 1 3570
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1680363874
transform 1 0 2280 0 1 3570
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1680363874
transform 1 0 2288 0 1 3570
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1680363874
transform 1 0 2296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1680363874
transform 1 0 2304 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1680363874
transform 1 0 2312 0 1 3570
box -8 -3 34 105
use FILL  FILL_2264
timestamp 1680363874
transform 1 0 2344 0 1 3570
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1680363874
transform 1 0 2352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1680363874
transform 1 0 2360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1680363874
transform 1 0 2368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1680363874
transform 1 0 2376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1680363874
transform 1 0 2384 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_67
timestamp 1680363874
transform 1 0 2392 0 1 3570
box -8 -3 34 105
use FILL  FILL_2275
timestamp 1680363874
transform 1 0 2424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1680363874
transform 1 0 2432 0 1 3570
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1680363874
transform 1 0 2440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1680363874
transform 1 0 2448 0 1 3570
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1680363874
transform 1 0 2456 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2258
timestamp 1680363874
transform 1 0 2484 0 1 3575
box -3 -3 3 3
use NOR2X1  NOR2X1_22
timestamp 1680363874
transform -1 0 2488 0 1 3570
box -8 -3 32 105
use FILL  FILL_2285
timestamp 1680363874
transform 1 0 2488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1680363874
transform 1 0 2496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1680363874
transform 1 0 2504 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_68
timestamp 1680363874
transform -1 0 2544 0 1 3570
box -8 -3 34 105
use INVX2  INVX2_177
timestamp 1680363874
transform -1 0 2560 0 1 3570
box -9 -3 26 105
use FILL  FILL_2288
timestamp 1680363874
transform 1 0 2560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1680363874
transform 1 0 2568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1680363874
transform 1 0 2576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1680363874
transform 1 0 2584 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_69
timestamp 1680363874
transform -1 0 2624 0 1 3570
box -8 -3 34 105
use FILL  FILL_2298
timestamp 1680363874
transform 1 0 2624 0 1 3570
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1680363874
transform 1 0 2632 0 1 3570
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1680363874
transform 1 0 2640 0 1 3570
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1680363874
transform 1 0 2648 0 1 3570
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1680363874
transform 1 0 2656 0 1 3570
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1680363874
transform 1 0 2664 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_153
timestamp 1680363874
transform 1 0 2672 0 1 3570
box -8 -3 46 105
use FILL  FILL_2314
timestamp 1680363874
transform 1 0 2712 0 1 3570
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1680363874
transform 1 0 2720 0 1 3570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1680363874
transform 1 0 2728 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_178
timestamp 1680363874
transform 1 0 2736 0 1 3570
box -9 -3 26 105
use FILL  FILL_2317
timestamp 1680363874
transform 1 0 2752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1680363874
transform 1 0 2760 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2259
timestamp 1680363874
transform 1 0 2780 0 1 3575
box -3 -3 3 3
use FILL  FILL_2320
timestamp 1680363874
transform 1 0 2768 0 1 3570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1680363874
transform 1 0 2776 0 1 3570
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1680363874
transform 1 0 2784 0 1 3570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1680363874
transform 1 0 2792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1680363874
transform 1 0 2800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1680363874
transform 1 0 2808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1680363874
transform 1 0 2816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1680363874
transform 1 0 2824 0 1 3570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1680363874
transform 1 0 2832 0 1 3570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1680363874
transform 1 0 2840 0 1 3570
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1680363874
transform 1 0 2848 0 1 3570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1680363874
transform 1 0 2856 0 1 3570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1680363874
transform 1 0 2864 0 1 3570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1680363874
transform 1 0 2872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1680363874
transform 1 0 2880 0 1 3570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1680363874
transform 1 0 2888 0 1 3570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1680363874
transform 1 0 2896 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_180
timestamp 1680363874
transform 1 0 2904 0 1 3570
box -9 -3 26 105
use FILL  FILL_2345
timestamp 1680363874
transform 1 0 2920 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_70
timestamp 1680363874
transform 1 0 2928 0 1 3570
box -8 -3 34 105
use FILL  FILL_2346
timestamp 1680363874
transform 1 0 2960 0 1 3570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1680363874
transform 1 0 2968 0 1 3570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1680363874
transform 1 0 2976 0 1 3570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1680363874
transform 1 0 2984 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_71
timestamp 1680363874
transform 1 0 2992 0 1 3570
box -8 -3 34 105
use FILL  FILL_2350
timestamp 1680363874
transform 1 0 3024 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2260
timestamp 1680363874
transform 1 0 3044 0 1 3575
box -3 -3 3 3
use FILL  FILL_2357
timestamp 1680363874
transform 1 0 3032 0 1 3570
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1680363874
transform 1 0 3040 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_72
timestamp 1680363874
transform 1 0 3048 0 1 3570
box -8 -3 34 105
use FILL  FILL_2361
timestamp 1680363874
transform 1 0 3080 0 1 3570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1680363874
transform 1 0 3088 0 1 3570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1680363874
transform 1 0 3096 0 1 3570
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1680363874
transform 1 0 3104 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1680363874
transform -1 0 3144 0 1 3570
box -8 -3 34 105
use FILL  FILL_2368
timestamp 1680363874
transform 1 0 3144 0 1 3570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1680363874
transform 1 0 3152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1680363874
transform 1 0 3160 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_23
timestamp 1680363874
transform 1 0 3168 0 1 3570
box -8 -3 32 105
use FILL  FILL_2375
timestamp 1680363874
transform 1 0 3192 0 1 3570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1680363874
transform 1 0 3200 0 1 3570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1680363874
transform 1 0 3208 0 1 3570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1680363874
transform 1 0 3216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1680363874
transform 1 0 3224 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_181
timestamp 1680363874
transform -1 0 3248 0 1 3570
box -9 -3 26 105
use FILL  FILL_2383
timestamp 1680363874
transform 1 0 3248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1680363874
transform 1 0 3256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1680363874
transform 1 0 3264 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_103
timestamp 1680363874
transform -1 0 3312 0 1 3570
box -8 -3 46 105
use FILL  FILL_2386
timestamp 1680363874
transform 1 0 3312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1680363874
transform 1 0 3320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1680363874
transform 1 0 3328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1680363874
transform 1 0 3336 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_182
timestamp 1680363874
transform -1 0 3360 0 1 3570
box -9 -3 26 105
use FILL  FILL_2390
timestamp 1680363874
transform 1 0 3360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1680363874
transform 1 0 3368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1680363874
transform 1 0 3376 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2261
timestamp 1680363874
transform 1 0 3420 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_104
timestamp 1680363874
transform -1 0 3424 0 1 3570
box -8 -3 46 105
use FILL  FILL_2393
timestamp 1680363874
transform 1 0 3424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1680363874
transform 1 0 3432 0 1 3570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1680363874
transform 1 0 3440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1680363874
transform 1 0 3448 0 1 3570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1680363874
transform 1 0 3456 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_183
timestamp 1680363874
transform -1 0 3480 0 1 3570
box -9 -3 26 105
use FILL  FILL_2410
timestamp 1680363874
transform 1 0 3480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1680363874
transform 1 0 3488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1680363874
transform 1 0 3496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1680363874
transform 1 0 3504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1680363874
transform 1 0 3512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1680363874
transform 1 0 3520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1680363874
transform 1 0 3528 0 1 3570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1680363874
transform 1 0 3536 0 1 3570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1680363874
transform 1 0 3544 0 1 3570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1680363874
transform 1 0 3552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1680363874
transform 1 0 3560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1680363874
transform 1 0 3568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1680363874
transform 1 0 3576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1680363874
transform 1 0 3584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1680363874
transform 1 0 3592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1680363874
transform 1 0 3600 0 1 3570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1680363874
transform 1 0 3608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1680363874
transform 1 0 3616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1680363874
transform 1 0 3624 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_155
timestamp 1680363874
transform 1 0 3632 0 1 3570
box -8 -3 46 105
use FILL  FILL_2441
timestamp 1680363874
transform 1 0 3672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1680363874
transform 1 0 3680 0 1 3570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1680363874
transform 1 0 3688 0 1 3570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1680363874
transform 1 0 3696 0 1 3570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1680363874
transform 1 0 3704 0 1 3570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1680363874
transform 1 0 3712 0 1 3570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1680363874
transform 1 0 3720 0 1 3570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1680363874
transform 1 0 3728 0 1 3570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1680363874
transform 1 0 3736 0 1 3570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1680363874
transform 1 0 3744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1680363874
transform 1 0 3752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1680363874
transform 1 0 3760 0 1 3570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1680363874
transform 1 0 3768 0 1 3570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1680363874
transform 1 0 3776 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_185
timestamp 1680363874
transform 1 0 3784 0 1 3570
box -9 -3 26 105
use FILL  FILL_2464
timestamp 1680363874
transform 1 0 3800 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2262
timestamp 1680363874
transform 1 0 3820 0 1 3575
box -3 -3 3 3
use FILL  FILL_2465
timestamp 1680363874
transform 1 0 3808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1680363874
transform 1 0 3816 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2263
timestamp 1680363874
transform 1 0 3844 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_107
timestamp 1680363874
transform 1 0 3824 0 1 3570
box -8 -3 46 105
use FILL  FILL_2467
timestamp 1680363874
transform 1 0 3864 0 1 3570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1680363874
transform 1 0 3872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1680363874
transform 1 0 3880 0 1 3570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1680363874
transform 1 0 3888 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_187
timestamp 1680363874
transform 1 0 3896 0 1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1680363874
transform -1 0 4008 0 1 3570
box -8 -3 104 105
use FILL  FILL_2479
timestamp 1680363874
transform 1 0 4008 0 1 3570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1680363874
transform 1 0 4016 0 1 3570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1680363874
transform 1 0 4024 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1680363874
transform 1 0 4032 0 1 3570
box -8 -3 104 105
use FILL  FILL_2482
timestamp 1680363874
transform 1 0 4128 0 1 3570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1680363874
transform 1 0 4136 0 1 3570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1680363874
transform 1 0 4144 0 1 3570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1680363874
transform 1 0 4152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1680363874
transform 1 0 4160 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2264
timestamp 1680363874
transform 1 0 4180 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_110
timestamp 1680363874
transform 1 0 4168 0 1 3570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1680363874
transform 1 0 4208 0 1 3570
box -8 -3 104 105
use FILL  FILL_2502
timestamp 1680363874
transform 1 0 4304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1680363874
transform 1 0 4312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1680363874
transform 1 0 4320 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_112
timestamp 1680363874
transform -1 0 4368 0 1 3570
box -8 -3 46 105
use FILL  FILL_2516
timestamp 1680363874
transform 1 0 4368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1680363874
transform 1 0 4376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1680363874
transform 1 0 4384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1680363874
transform 1 0 4392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1680363874
transform 1 0 4400 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2265
timestamp 1680363874
transform 1 0 4420 0 1 3575
box -3 -3 3 3
use FILL  FILL_2521
timestamp 1680363874
transform 1 0 4408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1680363874
transform 1 0 4416 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2266
timestamp 1680363874
transform 1 0 4436 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_189
timestamp 1680363874
transform 1 0 4424 0 1 3570
box -9 -3 26 105
use FILL  FILL_2531
timestamp 1680363874
transform 1 0 4440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1680363874
transform 1 0 4448 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_114
timestamp 1680363874
transform 1 0 4456 0 1 3570
box -8 -3 46 105
use FILL  FILL_2537
timestamp 1680363874
transform 1 0 4496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1680363874
transform 1 0 4504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1680363874
transform 1 0 4512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1680363874
transform 1 0 4520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1680363874
transform 1 0 4528 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1680363874
transform -1 0 4632 0 1 3570
box -8 -3 104 105
use AOI22X1  AOI22X1_115
timestamp 1680363874
transform 1 0 4632 0 1 3570
box -8 -3 46 105
use FILL  FILL_2542
timestamp 1680363874
transform 1 0 4672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1680363874
transform 1 0 4680 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_190
timestamp 1680363874
transform 1 0 4688 0 1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1680363874
transform -1 0 4800 0 1 3570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_23
timestamp 1680363874
transform 1 0 4827 0 1 3570
box -10 -3 10 3
use M3_M2  M3_M2_2298
timestamp 1680363874
transform 1 0 84 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1680363874
transform 1 0 4 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2553
timestamp 1680363874
transform 1 0 84 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2334
timestamp 1680363874
transform 1 0 164 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2654
timestamp 1680363874
transform 1 0 132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1680363874
transform 1 0 164 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2386
timestamp 1680363874
transform 1 0 132 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1680363874
transform 1 0 180 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1680363874
transform 1 0 196 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1680363874
transform 1 0 220 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1680363874
transform 1 0 236 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1680363874
transform 1 0 284 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2554
timestamp 1680363874
transform 1 0 236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1680363874
transform 1 0 284 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2433
timestamp 1680363874
transform 1 0 252 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2555
timestamp 1680363874
transform 1 0 332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1680363874
transform 1 0 324 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2354
timestamp 1680363874
transform 1 0 332 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2658
timestamp 1680363874
transform 1 0 340 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2301
timestamp 1680363874
transform 1 0 388 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2556
timestamp 1680363874
transform 1 0 388 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2335
timestamp 1680363874
transform 1 0 396 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2557
timestamp 1680363874
transform 1 0 404 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1680363874
transform 1 0 380 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1680363874
transform 1 0 396 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2388
timestamp 1680363874
transform 1 0 380 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2558
timestamp 1680363874
transform 1 0 428 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2336
timestamp 1680363874
transform 1 0 436 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1680363874
transform 1 0 468 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2559
timestamp 1680363874
transform 1 0 468 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2337
timestamp 1680363874
transform 1 0 476 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2560
timestamp 1680363874
transform 1 0 484 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1680363874
transform 1 0 500 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1680363874
transform 1 0 508 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1680363874
transform 1 0 476 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2441
timestamp 1680363874
transform 1 0 476 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1680363874
transform 1 0 556 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1680363874
transform 1 0 604 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1680363874
transform 1 0 596 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2563
timestamp 1680363874
transform 1 0 604 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1680363874
transform 1 0 620 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1680363874
transform 1 0 588 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1680363874
transform 1 0 596 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2355
timestamp 1680363874
transform 1 0 604 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2664
timestamp 1680363874
transform 1 0 612 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2339
timestamp 1680363874
transform 1 0 628 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1680363874
transform 1 0 620 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1680363874
transform 1 0 644 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2749
timestamp 1680363874
transform 1 0 652 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2340
timestamp 1680363874
transform 1 0 676 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1680363874
transform 1 0 684 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1680363874
transform 1 0 708 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2665
timestamp 1680363874
transform 1 0 708 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2356
timestamp 1680363874
transform 1 0 716 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2750
timestamp 1680363874
transform 1 0 732 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1680363874
transform 1 0 764 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1680363874
transform 1 0 772 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1680363874
transform 1 0 788 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2305
timestamp 1680363874
transform 1 0 812 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2567
timestamp 1680363874
transform 1 0 812 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1680363874
transform 1 0 820 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2391
timestamp 1680363874
transform 1 0 836 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1680363874
transform 1 0 868 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2666
timestamp 1680363874
transform 1 0 868 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1680363874
transform 1 0 884 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1680363874
transform 1 0 900 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1680363874
transform 1 0 924 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1680363874
transform 1 0 932 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2307
timestamp 1680363874
transform 1 0 996 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1680363874
transform 1 0 1012 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2569
timestamp 1680363874
transform 1 0 980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1680363874
transform 1 0 996 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2341
timestamp 1680363874
transform 1 0 1004 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2571
timestamp 1680363874
transform 1 0 1012 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1680363874
transform 1 0 1020 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2357
timestamp 1680363874
transform 1 0 980 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2669
timestamp 1680363874
transform 1 0 988 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1680363874
transform 1 0 1004 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2342
timestamp 1680363874
transform 1 0 1028 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1680363874
transform 1 0 1020 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1680363874
transform 1 0 1052 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1680363874
transform 1 0 1084 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2573
timestamp 1680363874
transform 1 0 1068 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1680363874
transform 1 0 1084 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1680363874
transform 1 0 1060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1680363874
transform 1 0 1076 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2359
timestamp 1680363874
transform 1 0 1084 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1680363874
transform 1 0 1100 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1680363874
transform 1 0 1260 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2575
timestamp 1680363874
transform 1 0 1228 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2360
timestamp 1680363874
transform 1 0 1228 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2673
timestamp 1680363874
transform 1 0 1252 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2361
timestamp 1680363874
transform 1 0 1308 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1680363874
transform 1 0 1276 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2674
timestamp 1680363874
transform 1 0 1332 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1680363874
transform 1 0 1348 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1680363874
transform 1 0 1356 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1680363874
transform 1 0 1364 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2310
timestamp 1680363874
transform 1 0 1396 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2578
timestamp 1680363874
transform 1 0 1396 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2343
timestamp 1680363874
transform 1 0 1404 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2579
timestamp 1680363874
transform 1 0 1412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1680363874
transform 1 0 1388 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1680363874
transform 1 0 1404 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1680363874
transform 1 0 1444 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2311
timestamp 1680363874
transform 1 0 1484 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1680363874
transform 1 0 1532 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2580
timestamp 1680363874
transform 1 0 1532 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1680363874
transform 1 0 1484 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2313
timestamp 1680363874
transform 1 0 1572 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2581
timestamp 1680363874
transform 1 0 1572 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2362
timestamp 1680363874
transform 1 0 1572 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2680
timestamp 1680363874
transform 1 0 1588 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1680363874
transform 1 0 1596 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2363
timestamp 1680363874
transform 1 0 1604 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2583
timestamp 1680363874
transform 1 0 1636 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1680363874
transform 1 0 1620 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2393
timestamp 1680363874
transform 1 0 1620 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1680363874
transform 1 0 1652 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2584
timestamp 1680363874
transform 1 0 1644 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2364
timestamp 1680363874
transform 1 0 1660 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2682
timestamp 1680363874
transform 1 0 1676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1680363874
transform 1 0 1660 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2394
timestamp 1680363874
transform 1 0 1676 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2585
timestamp 1680363874
transform 1 0 1692 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1680363874
transform 1 0 1716 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1680363874
transform 1 0 1748 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1680363874
transform 1 0 1732 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2365
timestamp 1680363874
transform 1 0 1748 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1680363874
transform 1 0 1732 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2755
timestamp 1680363874
transform 1 0 1748 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2269
timestamp 1680363874
transform 1 0 1764 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2588
timestamp 1680363874
transform 1 0 1796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1680363874
transform 1 0 1788 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1680363874
transform 1 0 1820 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1680363874
transform 1 0 1828 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2396
timestamp 1680363874
transform 1 0 1828 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2589
timestamp 1680363874
transform 1 0 1860 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1680363874
transform 1 0 1876 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2366
timestamp 1680363874
transform 1 0 1900 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2686
timestamp 1680363874
transform 1 0 1908 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1680363874
transform 1 0 1900 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2397
timestamp 1680363874
transform 1 0 1908 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2591
timestamp 1680363874
transform 1 0 1932 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1680363874
transform 1 0 1948 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2367
timestamp 1680363874
transform 1 0 1972 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2687
timestamp 1680363874
transform 1 0 1980 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1680363874
transform 1 0 1972 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2398
timestamp 1680363874
transform 1 0 1980 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1680363874
transform 1 0 2020 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1680363874
transform 1 0 2020 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2593
timestamp 1680363874
transform 1 0 2020 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1680363874
transform 1 0 2028 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2286
timestamp 1680363874
transform 1 0 2052 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1680363874
transform 1 0 2052 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2688
timestamp 1680363874
transform 1 0 2060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1680363874
transform 1 0 2052 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2399
timestamp 1680363874
transform 1 0 2060 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2595
timestamp 1680363874
transform 1 0 2084 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1680363874
transform 1 0 2092 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2344
timestamp 1680363874
transform 1 0 2116 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1680363874
transform 1 0 2140 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1680363874
transform 1 0 2132 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2689
timestamp 1680363874
transform 1 0 2140 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1680363874
transform 1 0 2132 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2400
timestamp 1680363874
transform 1 0 2140 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2597
timestamp 1680363874
transform 1 0 2164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1680363874
transform 1 0 2172 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1680363874
transform 1 0 2196 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2370
timestamp 1680363874
transform 1 0 2204 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2761
timestamp 1680363874
transform 1 0 2204 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1680363874
transform 1 0 2236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1680363874
transform 1 0 2252 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2371
timestamp 1680363874
transform 1 0 2276 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1680363874
transform 1 0 2252 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1680363874
transform 1 0 2268 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2762
timestamp 1680363874
transform 1 0 2276 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1680363874
transform 1 0 2284 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2403
timestamp 1680363874
transform 1 0 2292 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1680363874
transform 1 0 2308 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2600
timestamp 1680363874
transform 1 0 2308 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2272
timestamp 1680363874
transform 1 0 2348 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2693
timestamp 1680363874
transform 1 0 2332 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2372
timestamp 1680363874
transform 1 0 2348 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1680363874
transform 1 0 2332 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2763
timestamp 1680363874
transform 1 0 2348 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1680363874
transform 1 0 2356 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2287
timestamp 1680363874
transform 1 0 2380 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2601
timestamp 1680363874
transform 1 0 2380 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1680363874
transform 1 0 2396 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2288
timestamp 1680363874
transform 1 0 2412 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2602
timestamp 1680363874
transform 1 0 2436 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2443
timestamp 1680363874
transform 1 0 2436 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2603
timestamp 1680363874
transform 1 0 2452 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1680363874
transform 1 0 2500 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1680363874
transform 1 0 2500 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1680363874
transform 1 0 2460 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2697
timestamp 1680363874
transform 1 0 2540 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2406
timestamp 1680363874
transform 1 0 2628 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2604
timestamp 1680363874
transform 1 0 2676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1680363874
transform 1 0 2724 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2445
timestamp 1680363874
transform 1 0 2732 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1680363874
transform 1 0 2788 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2605
timestamp 1680363874
transform 1 0 2788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1680363874
transform 1 0 2780 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2446
timestamp 1680363874
transform 1 0 2780 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2606
timestamp 1680363874
transform 1 0 2836 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1680363874
transform 1 0 2820 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1680363874
transform 1 0 2844 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2407
timestamp 1680363874
transform 1 0 2844 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1680363874
transform 1 0 2820 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1680363874
transform 1 0 2836 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2607
timestamp 1680363874
transform 1 0 2876 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2316
timestamp 1680363874
transform 1 0 2900 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1680363874
transform 1 0 2980 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2608
timestamp 1680363874
transform 1 0 2980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1680363874
transform 1 0 2900 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1680363874
transform 1 0 2932 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2408
timestamp 1680363874
transform 1 0 2932 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1680363874
transform 1 0 2916 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2609
timestamp 1680363874
transform 1 0 3012 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1680363874
transform 1 0 3084 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1680363874
transform 1 0 3092 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1680363874
transform 1 0 3052 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1680363874
transform 1 0 3060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1680363874
transform 1 0 3076 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2373
timestamp 1680363874
transform 1 0 3084 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2764
timestamp 1680363874
transform 1 0 3076 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1680363874
transform 1 0 3100 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2425
timestamp 1680363874
transform 1 0 3092 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1680363874
transform 1 0 3100 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1680363874
transform 1 0 3148 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2766
timestamp 1680363874
transform 1 0 3140 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2435
timestamp 1680363874
transform 1 0 3140 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2767
timestamp 1680363874
transform 1 0 3148 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1680363874
transform 1 0 3180 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2318
timestamp 1680363874
transform 1 0 3188 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2613
timestamp 1680363874
transform 1 0 3188 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2375
timestamp 1680363874
transform 1 0 3180 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2707
timestamp 1680363874
transform 1 0 3204 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2409
timestamp 1680363874
transform 1 0 3204 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2708
timestamp 1680363874
transform 1 0 3236 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2273
timestamp 1680363874
transform 1 0 3268 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1680363874
transform 1 0 3292 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2614
timestamp 1680363874
transform 1 0 3324 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1680363874
transform 1 0 3300 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2410
timestamp 1680363874
transform 1 0 3252 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2551
timestamp 1680363874
transform 1 0 3356 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1680363874
transform 1 0 3356 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2275
timestamp 1680363874
transform 1 0 3388 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1680363874
transform 1 0 3380 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2710
timestamp 1680363874
transform 1 0 3380 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2320
timestamp 1680363874
transform 1 0 3420 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2616
timestamp 1680363874
transform 1 0 3436 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2411
timestamp 1680363874
transform 1 0 3436 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1680363874
transform 1 0 3452 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2617
timestamp 1680363874
transform 1 0 3460 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2346
timestamp 1680363874
transform 1 0 3492 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2618
timestamp 1680363874
transform 1 0 3516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1680363874
transform 1 0 3484 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1680363874
transform 1 0 3492 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1680363874
transform 1 0 3508 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2412
timestamp 1680363874
transform 1 0 3508 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2714
timestamp 1680363874
transform 1 0 3548 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1680363874
transform 1 0 3548 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2619
timestamp 1680363874
transform 1 0 3572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1680363874
transform 1 0 3564 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1680363874
transform 1 0 3580 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1680363874
transform 1 0 3604 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2347
timestamp 1680363874
transform 1 0 3620 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2717
timestamp 1680363874
transform 1 0 3620 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2321
timestamp 1680363874
transform 1 0 3652 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2718
timestamp 1680363874
transform 1 0 3644 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2376
timestamp 1680363874
transform 1 0 3668 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2768
timestamp 1680363874
transform 1 0 3668 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1680363874
transform 1 0 3676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1680363874
transform 1 0 3708 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1680363874
transform 1 0 3716 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1680363874
transform 1 0 3732 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2377
timestamp 1680363874
transform 1 0 3708 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2720
timestamp 1680363874
transform 1 0 3716 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1680363874
transform 1 0 3740 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2436
timestamp 1680363874
transform 1 0 3748 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1680363874
transform 1 0 3764 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1680363874
transform 1 0 3788 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1680363874
transform 1 0 3780 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1680363874
transform 1 0 3772 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1680363874
transform 1 0 3828 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2624
timestamp 1680363874
transform 1 0 3780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1680363874
transform 1 0 3788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1680363874
transform 1 0 3796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1680363874
transform 1 0 3812 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1680363874
transform 1 0 3820 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1680363874
transform 1 0 3804 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2413
timestamp 1680363874
transform 1 0 3804 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2723
timestamp 1680363874
transform 1 0 3828 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2427
timestamp 1680363874
transform 1 0 3828 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1680363874
transform 1 0 3876 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1680363874
transform 1 0 3868 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2629
timestamp 1680363874
transform 1 0 3868 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1680363874
transform 1 0 3876 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2414
timestamp 1680363874
transform 1 0 3868 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2725
timestamp 1680363874
transform 1 0 3908 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1680363874
transform 1 0 3932 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1680363874
transform 1 0 3932 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1680363874
transform 1 0 3948 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1680363874
transform 1 0 3964 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1680363874
transform 1 0 3964 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2631
timestamp 1680363874
transform 1 0 3964 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1680363874
transform 1 0 3956 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1680363874
transform 1 0 3972 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2416
timestamp 1680363874
transform 1 0 3964 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1680363874
transform 1 0 3940 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1680363874
transform 1 0 3972 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1680363874
transform 1 0 3972 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2632
timestamp 1680363874
transform 1 0 4100 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1680363874
transform 1 0 4068 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2291
timestamp 1680363874
transform 1 0 4116 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2633
timestamp 1680363874
transform 1 0 4116 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2378
timestamp 1680363874
transform 1 0 4116 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2769
timestamp 1680363874
transform 1 0 4116 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2324
timestamp 1680363874
transform 1 0 4164 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2634
timestamp 1680363874
transform 1 0 4164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1680363874
transform 1 0 4180 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1680363874
transform 1 0 4188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1680363874
transform 1 0 4156 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1680363874
transform 1 0 4172 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1680363874
transform 1 0 4188 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1680363874
transform 1 0 4196 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2428
timestamp 1680363874
transform 1 0 4156 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1680363874
transform 1 0 4188 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1680363874
transform 1 0 4196 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1680363874
transform 1 0 4188 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1680363874
transform 1 0 4236 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1680363874
transform 1 0 4260 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2733
timestamp 1680363874
transform 1 0 4260 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1680363874
transform 1 0 4276 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1680363874
transform 1 0 4300 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1680363874
transform 1 0 4300 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2418
timestamp 1680363874
transform 1 0 4300 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1680363874
transform 1 0 4316 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2735
timestamp 1680363874
transform 1 0 4332 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2325
timestamp 1680363874
transform 1 0 4356 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1680363874
transform 1 0 4396 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2638
timestamp 1680363874
transform 1 0 4380 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1680363874
transform 1 0 4396 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1680363874
transform 1 0 4388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2379
timestamp 1680363874
transform 1 0 4396 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1680363874
transform 1 0 4380 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1680363874
transform 1 0 4396 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1680363874
transform 1 0 4420 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2640
timestamp 1680363874
transform 1 0 4412 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2380
timestamp 1680363874
transform 1 0 4412 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2770
timestamp 1680363874
transform 1 0 4412 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2381
timestamp 1680363874
transform 1 0 4428 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2737
timestamp 1680363874
transform 1 0 4436 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1680363874
transform 1 0 4452 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2327
timestamp 1680363874
transform 1 0 4476 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1680363874
transform 1 0 4508 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1680363874
transform 1 0 4524 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2641
timestamp 1680363874
transform 1 0 4492 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2349
timestamp 1680363874
transform 1 0 4500 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1680363874
transform 1 0 4532 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2642
timestamp 1680363874
transform 1 0 4508 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1680363874
transform 1 0 4524 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1680363874
transform 1 0 4532 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1680363874
transform 1 0 4500 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1680363874
transform 1 0 4516 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2420
timestamp 1680363874
transform 1 0 4500 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1680363874
transform 1 0 4516 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1680363874
transform 1 0 4548 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1680363874
transform 1 0 4564 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1680363874
transform 1 0 4580 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1680363874
transform 1 0 4620 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1680363874
transform 1 0 4612 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2645
timestamp 1680363874
transform 1 0 4580 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1680363874
transform 1 0 4596 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1680363874
transform 1 0 4604 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1680363874
transform 1 0 4620 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1680363874
transform 1 0 4572 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1680363874
transform 1 0 4588 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1680363874
transform 1 0 4612 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2383
timestamp 1680363874
transform 1 0 4620 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1680363874
transform 1 0 4644 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2649
timestamp 1680363874
transform 1 0 4636 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2296
timestamp 1680363874
transform 1 0 4660 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1680363874
transform 1 0 4676 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1680363874
transform 1 0 4660 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2650
timestamp 1680363874
transform 1 0 4676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1680363874
transform 1 0 4684 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1680363874
transform 1 0 4692 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2297
timestamp 1680363874
transform 1 0 4708 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1680363874
transform 1 0 4700 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1680363874
transform 1 0 4748 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2653
timestamp 1680363874
transform 1 0 4788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1680363874
transform 1 0 4652 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1680363874
transform 1 0 4668 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2384
timestamp 1680363874
transform 1 0 4676 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1680363874
transform 1 0 4692 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2746
timestamp 1680363874
transform 1 0 4700 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1680363874
transform 1 0 4708 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1680363874
transform 1 0 4748 0 1 3525
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_24
timestamp 1680363874
transform 1 0 24 0 1 3470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_174
timestamp 1680363874
transform 1 0 72 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2002
timestamp 1680363874
transform 1 0 168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1680363874
transform 1 0 176 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1680363874
transform 1 0 184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1680363874
transform 1 0 192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1680363874
transform 1 0 200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1680363874
transform 1 0 208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1680363874
transform 1 0 216 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1680363874
transform 1 0 224 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2012
timestamp 1680363874
transform 1 0 320 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1680363874
transform 1 0 328 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1680363874
transform 1 0 336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1680363874
transform 1 0 344 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1680363874
transform 1 0 352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1680363874
transform 1 0 360 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_139
timestamp 1680363874
transform 1 0 368 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2026
timestamp 1680363874
transform 1 0 408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1680363874
transform 1 0 416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1680363874
transform 1 0 424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1680363874
transform 1 0 432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1680363874
transform 1 0 440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1680363874
transform 1 0 448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1680363874
transform 1 0 456 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_140
timestamp 1680363874
transform -1 0 504 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2033
timestamp 1680363874
transform 1 0 504 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1680363874
transform 1 0 512 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1680363874
transform 1 0 520 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1680363874
transform 1 0 528 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_171
timestamp 1680363874
transform 1 0 536 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2039
timestamp 1680363874
transform 1 0 552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1680363874
transform 1 0 560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1680363874
transform 1 0 568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1680363874
transform 1 0 576 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_142
timestamp 1680363874
transform 1 0 584 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2051
timestamp 1680363874
transform 1 0 624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1680363874
transform 1 0 632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1680363874
transform 1 0 640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1680363874
transform 1 0 648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1680363874
transform 1 0 656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1680363874
transform 1 0 664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1680363874
transform 1 0 672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1680363874
transform 1 0 680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1680363874
transform 1 0 688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1680363874
transform 1 0 696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1680363874
transform 1 0 704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1680363874
transform 1 0 712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1680363874
transform 1 0 720 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_10
timestamp 1680363874
transform -1 0 752 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2072
timestamp 1680363874
transform 1 0 752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1680363874
transform 1 0 760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1680363874
transform 1 0 768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1680363874
transform 1 0 776 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_47
timestamp 1680363874
transform -1 0 816 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2081
timestamp 1680363874
transform 1 0 816 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1680363874
transform 1 0 824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1680363874
transform 1 0 832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1680363874
transform 1 0 840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1680363874
transform 1 0 848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1680363874
transform 1 0 856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1680363874
transform 1 0 864 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_49
timestamp 1680363874
transform 1 0 872 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2096
timestamp 1680363874
transform 1 0 904 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1680363874
transform 1 0 912 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2097
timestamp 1680363874
transform 1 0 936 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1680363874
transform 1 0 944 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1680363874
transform 1 0 952 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1680363874
transform 1 0 960 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1680363874
transform 1 0 968 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_145
timestamp 1680363874
transform 1 0 976 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2108
timestamp 1680363874
transform 1 0 1016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1680363874
transform 1 0 1024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1680363874
transform 1 0 1032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1680363874
transform 1 0 1040 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_147
timestamp 1680363874
transform 1 0 1048 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2116
timestamp 1680363874
transform 1 0 1088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1680363874
transform 1 0 1096 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1680363874
transform 1 0 1104 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1680363874
transform 1 0 1112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1680363874
transform 1 0 1120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1680363874
transform 1 0 1128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1680363874
transform 1 0 1136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1680363874
transform 1 0 1144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1680363874
transform 1 0 1152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1680363874
transform 1 0 1160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1680363874
transform 1 0 1168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1680363874
transform 1 0 1176 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1680363874
transform 1 0 1184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1680363874
transform 1 0 1192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1680363874
transform 1 0 1200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1680363874
transform 1 0 1208 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1680363874
transform 1 0 1216 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2147
timestamp 1680363874
transform 1 0 1312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1680363874
transform 1 0 1320 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1680363874
transform 1 0 1328 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_173
timestamp 1680363874
transform -1 0 1352 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2150
timestamp 1680363874
transform 1 0 1352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1680363874
transform 1 0 1360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1680363874
transform 1 0 1368 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_152
timestamp 1680363874
transform -1 0 1416 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2157
timestamp 1680363874
transform 1 0 1416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1680363874
transform 1 0 1424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1680363874
transform 1 0 1432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1680363874
transform 1 0 1440 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1680363874
transform -1 0 1544 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2167
timestamp 1680363874
transform 1 0 1544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1680363874
transform 1 0 1552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1680363874
transform 1 0 1560 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_175
timestamp 1680363874
transform 1 0 1568 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2170
timestamp 1680363874
transform 1 0 1584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1680363874
transform 1 0 1592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1680363874
transform 1 0 1600 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_51
timestamp 1680363874
transform 1 0 1608 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2176
timestamp 1680363874
transform 1 0 1640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1680363874
transform 1 0 1648 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_52
timestamp 1680363874
transform -1 0 1688 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2184
timestamp 1680363874
transform 1 0 1688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1680363874
transform 1 0 1696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1680363874
transform 1 0 1704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1680363874
transform 1 0 1712 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1680363874
transform 1 0 1720 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2198
timestamp 1680363874
transform 1 0 1752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1680363874
transform 1 0 1760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1680363874
transform 1 0 1768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1680363874
transform 1 0 1776 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1680363874
transform 1 0 1784 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1680363874
transform 1 0 1792 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1680363874
transform -1 0 1832 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2204
timestamp 1680363874
transform 1 0 1832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1680363874
transform 1 0 1840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1680363874
transform 1 0 1848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1680363874
transform 1 0 1856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1680363874
transform 1 0 1864 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1680363874
transform 1 0 1872 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2213
timestamp 1680363874
transform 1 0 1904 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1680363874
transform 1 0 1912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1680363874
transform 1 0 1920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1680363874
transform 1 0 1928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1680363874
transform 1 0 1936 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_58
timestamp 1680363874
transform 1 0 1944 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2218
timestamp 1680363874
transform 1 0 1976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1680363874
transform 1 0 1984 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1680363874
transform 1 0 1992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1680363874
transform 1 0 2000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1680363874
transform 1 0 2008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1680363874
transform 1 0 2016 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_59
timestamp 1680363874
transform 1 0 2024 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2227
timestamp 1680363874
transform 1 0 2056 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1680363874
transform 1 0 2064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1680363874
transform 1 0 2072 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1680363874
transform 1 0 2080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1680363874
transform 1 0 2088 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2449
timestamp 1680363874
transform 1 0 2108 0 1 3475
box -3 -3 3 3
use OAI21X1  OAI21X1_61
timestamp 1680363874
transform 1 0 2096 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2237
timestamp 1680363874
transform 1 0 2128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1680363874
transform 1 0 2136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1680363874
transform 1 0 2144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1680363874
transform 1 0 2152 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2450
timestamp 1680363874
transform 1 0 2172 0 1 3475
box -3 -3 3 3
use FILL  FILL_2242
timestamp 1680363874
transform 1 0 2160 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1680363874
transform 1 0 2168 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2247
timestamp 1680363874
transform 1 0 2200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1680363874
transform 1 0 2208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1680363874
transform 1 0 2216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1680363874
transform 1 0 2224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1680363874
transform 1 0 2232 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1680363874
transform 1 0 2240 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1680363874
transform 1 0 2248 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2257
timestamp 1680363874
transform 1 0 2280 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1680363874
transform 1 0 2288 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1680363874
transform 1 0 2296 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1680363874
transform 1 0 2304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1680363874
transform 1 0 2312 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1680363874
transform 1 0 2320 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2267
timestamp 1680363874
transform 1 0 2352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1680363874
transform 1 0 2360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1680363874
transform 1 0 2368 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2451
timestamp 1680363874
transform 1 0 2388 0 1 3475
box -3 -3 3 3
use FILL  FILL_2273
timestamp 1680363874
transform 1 0 2376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1680363874
transform 1 0 2384 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_176
timestamp 1680363874
transform -1 0 2408 0 -1 3570
box -9 -3 26 105
use M3_M2  M3_M2_2452
timestamp 1680363874
transform 1 0 2420 0 1 3475
box -3 -3 3 3
use FILL  FILL_2277
timestamp 1680363874
transform 1 0 2408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1680363874
transform 1 0 2416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1680363874
transform 1 0 2424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1680363874
transform 1 0 2432 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1680363874
transform 1 0 2440 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2289
timestamp 1680363874
transform 1 0 2536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1680363874
transform 1 0 2544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1680363874
transform 1 0 2552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1680363874
transform 1 0 2560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1680363874
transform 1 0 2568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1680363874
transform 1 0 2576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1680363874
transform 1 0 2584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1680363874
transform 1 0 2592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1680363874
transform 1 0 2600 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1680363874
transform 1 0 2608 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1680363874
transform 1 0 2616 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1680363874
transform 1 0 2624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1680363874
transform 1 0 2632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1680363874
transform 1 0 2640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1680363874
transform 1 0 2648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1680363874
transform 1 0 2656 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1680363874
transform 1 0 2664 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2319
timestamp 1680363874
transform 1 0 2760 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_179
timestamp 1680363874
transform 1 0 2768 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2323
timestamp 1680363874
transform 1 0 2784 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1680363874
transform 1 0 2792 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1680363874
transform 1 0 2800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1680363874
transform 1 0 2808 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_154
timestamp 1680363874
transform 1 0 2816 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2336
timestamp 1680363874
transform 1 0 2856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1680363874
transform 1 0 2864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1680363874
transform 1 0 2872 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1680363874
transform 1 0 2880 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1680363874
transform 1 0 2888 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1680363874
transform -1 0 2992 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2352
timestamp 1680363874
transform 1 0 2992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1680363874
transform 1 0 3000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1680363874
transform 1 0 3008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1680363874
transform 1 0 3016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1680363874
transform 1 0 3024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1680363874
transform 1 0 3032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1680363874
transform 1 0 3040 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_73
timestamp 1680363874
transform 1 0 3048 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2362
timestamp 1680363874
transform 1 0 3080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1680363874
transform 1 0 3088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1680363874
transform 1 0 3096 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1680363874
transform 1 0 3104 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_75
timestamp 1680363874
transform 1 0 3112 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2370
timestamp 1680363874
transform 1 0 3144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1680363874
transform 1 0 3152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1680363874
transform 1 0 3160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1680363874
transform 1 0 3168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1680363874
transform 1 0 3176 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_76
timestamp 1680363874
transform -1 0 3216 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2381
timestamp 1680363874
transform 1 0 3216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1680363874
transform 1 0 3224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1680363874
transform 1 0 3232 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1680363874
transform -1 0 3336 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2396
timestamp 1680363874
transform 1 0 3336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1680363874
transform 1 0 3344 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_24
timestamp 1680363874
transform 1 0 3352 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2398
timestamp 1680363874
transform 1 0 3376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1680363874
transform 1 0 3384 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1680363874
transform 1 0 3392 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1680363874
transform 1 0 3400 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1680363874
transform 1 0 3408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1680363874
transform 1 0 3416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1680363874
transform 1 0 3424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1680363874
transform 1 0 3432 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_184
timestamp 1680363874
transform 1 0 3440 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2417
timestamp 1680363874
transform 1 0 3456 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1680363874
transform 1 0 3464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1680363874
transform 1 0 3472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1680363874
transform 1 0 3480 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_105
timestamp 1680363874
transform -1 0 3528 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2421
timestamp 1680363874
transform 1 0 3528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1680363874
transform 1 0 3536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1680363874
transform 1 0 3544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1680363874
transform 1 0 3552 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_106
timestamp 1680363874
transform 1 0 3560 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2434
timestamp 1680363874
transform 1 0 3600 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1680363874
transform 1 0 3608 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1680363874
transform 1 0 3616 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1680363874
transform 1 0 3624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1680363874
transform 1 0 3632 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2453
timestamp 1680363874
transform 1 0 3660 0 1 3475
box -3 -3 3 3
use OAI21X1  OAI21X1_77
timestamp 1680363874
transform 1 0 3640 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2443
timestamp 1680363874
transform 1 0 3672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1680363874
transform 1 0 3680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1680363874
transform 1 0 3688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1680363874
transform 1 0 3696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1680363874
transform 1 0 3704 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_156
timestamp 1680363874
transform 1 0 3712 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2458
timestamp 1680363874
transform 1 0 3752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1680363874
transform 1 0 3760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1680363874
transform 1 0 3768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1680363874
transform 1 0 3776 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_108
timestamp 1680363874
transform -1 0 3824 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2470
timestamp 1680363874
transform 1 0 3824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1680363874
transform 1 0 3832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1680363874
transform 1 0 3840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1680363874
transform 1 0 3848 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_186
timestamp 1680363874
transform -1 0 3872 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2474
timestamp 1680363874
transform 1 0 3872 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1680363874
transform 1 0 3880 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1680363874
transform 1 0 3888 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1680363874
transform 1 0 3896 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1680363874
transform 1 0 3904 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1680363874
transform 1 0 3912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1680363874
transform 1 0 3920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1680363874
transform 1 0 3928 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_109
timestamp 1680363874
transform 1 0 3936 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2488
timestamp 1680363874
transform 1 0 3976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1680363874
transform 1 0 3984 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1680363874
transform 1 0 3992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1680363874
transform 1 0 4000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1680363874
transform 1 0 4008 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2454
timestamp 1680363874
transform 1 0 4116 0 1 3475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_188
timestamp 1680363874
transform -1 0 4112 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2493
timestamp 1680363874
transform 1 0 4112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1680363874
transform 1 0 4120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1680363874
transform 1 0 4128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1680363874
transform 1 0 4136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1680363874
transform 1 0 4144 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_111
timestamp 1680363874
transform 1 0 4152 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2503
timestamp 1680363874
transform 1 0 4192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1680363874
transform 1 0 4200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1680363874
transform 1 0 4208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1680363874
transform 1 0 4216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1680363874
transform 1 0 4224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1680363874
transform 1 0 4232 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_188
timestamp 1680363874
transform 1 0 4240 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2509
timestamp 1680363874
transform 1 0 4256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1680363874
transform 1 0 4264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1680363874
transform 1 0 4272 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_25
timestamp 1680363874
transform -1 0 4304 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2512
timestamp 1680363874
transform 1 0 4304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1680363874
transform 1 0 4312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1680363874
transform 1 0 4320 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1680363874
transform 1 0 4328 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1680363874
transform 1 0 4336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1680363874
transform 1 0 4344 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1680363874
transform 1 0 4352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1680363874
transform 1 0 4360 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_113
timestamp 1680363874
transform -1 0 4408 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2528
timestamp 1680363874
transform 1 0 4408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1680363874
transform 1 0 4416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1680363874
transform 1 0 4424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1680363874
transform 1 0 4432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1680363874
transform 1 0 4440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1680363874
transform 1 0 4448 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_191
timestamp 1680363874
transform 1 0 4456 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2544
timestamp 1680363874
transform 1 0 4472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1680363874
transform 1 0 4480 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_157
timestamp 1680363874
transform 1 0 4488 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2546
timestamp 1680363874
transform 1 0 4528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1680363874
transform 1 0 4536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1680363874
transform 1 0 4544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1680363874
transform 1 0 4552 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_192
timestamp 1680363874
transform 1 0 4560 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1680363874
transform 1 0 4576 0 -1 3570
box -9 -3 26 105
use AOI22X1  AOI22X1_116
timestamp 1680363874
transform -1 0 4632 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2550
timestamp 1680363874
transform 1 0 4632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1680363874
transform 1 0 4640 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_117
timestamp 1680363874
transform 1 0 4648 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_194
timestamp 1680363874
transform 1 0 4688 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1680363874
transform -1 0 4800 0 -1 3570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_25
timestamp 1680363874
transform 1 0 4851 0 1 3470
box -10 -3 10 3
use M3_M2  M3_M2_2543
timestamp 1680363874
transform 1 0 132 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2881
timestamp 1680363874
transform 1 0 132 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2472
timestamp 1680363874
transform 1 0 188 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1680363874
transform 1 0 164 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2779
timestamp 1680363874
transform 1 0 172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1680363874
transform 1 0 188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1680363874
transform 1 0 164 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2561
timestamp 1680363874
transform 1 0 172 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2883
timestamp 1680363874
transform 1 0 180 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2578
timestamp 1680363874
transform 1 0 164 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1680363874
transform 1 0 196 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2884
timestamp 1680363874
transform 1 0 212 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2482
timestamp 1680363874
transform 1 0 252 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1680363874
transform 1 0 228 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1680363874
transform 1 0 260 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2781
timestamp 1680363874
transform 1 0 276 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1680363874
transform 1 0 228 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2580
timestamp 1680363874
transform 1 0 276 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1680363874
transform 1 0 220 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1680363874
transform 1 0 252 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2782
timestamp 1680363874
transform 1 0 316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1680363874
transform 1 0 324 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1680363874
transform 1 0 340 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2473
timestamp 1680363874
transform 1 0 388 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2784
timestamp 1680363874
transform 1 0 356 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2545
timestamp 1680363874
transform 1 0 364 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2785
timestamp 1680363874
transform 1 0 388 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1680363874
transform 1 0 364 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1680363874
transform 1 0 380 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2581
timestamp 1680363874
transform 1 0 380 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2889
timestamp 1680363874
transform 1 0 412 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2510
timestamp 1680363874
transform 1 0 452 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2786
timestamp 1680363874
transform 1 0 428 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1680363874
transform 1 0 420 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1680363874
transform 1 0 436 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1680363874
transform 1 0 476 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2547
timestamp 1680363874
transform 1 0 500 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2788
timestamp 1680363874
transform 1 0 532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1680363874
transform 1 0 436 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1680363874
transform 1 0 452 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2582
timestamp 1680363874
transform 1 0 436 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1680363874
transform 1 0 476 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1680363874
transform 1 0 444 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2789
timestamp 1680363874
transform 1 0 556 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1680363874
transform 1 0 588 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2511
timestamp 1680363874
transform 1 0 620 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2790
timestamp 1680363874
transform 1 0 620 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1680363874
transform 1 0 636 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2483
timestamp 1680363874
transform 1 0 652 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2771
timestamp 1680363874
transform 1 0 652 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1680363874
transform 1 0 628 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1680363874
transform 1 0 644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1680363874
transform 1 0 628 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1680363874
transform 1 0 652 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1680363874
transform 1 0 668 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1680363874
transform 1 0 684 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2792
timestamp 1680363874
transform 1 0 684 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1680363874
transform 1 0 700 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1680363874
transform 1 0 780 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1680363874
transform 1 0 788 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1680363874
transform 1 0 772 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1680363874
transform 1 0 804 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1680363874
transform 1 0 804 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1680363874
transform 1 0 828 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1680363874
transform 1 0 820 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1680363874
transform 1 0 900 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2548
timestamp 1680363874
transform 1 0 908 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1680363874
transform 1 0 900 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1680363874
transform 1 0 940 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2897
timestamp 1680363874
transform 1 0 932 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1680363874
transform 1 0 940 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1680363874
transform 1 0 932 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2898
timestamp 1680363874
transform 1 0 1028 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1680363874
transform 1 0 1068 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1680363874
transform 1 0 1068 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1680363874
transform 1 0 1084 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2513
timestamp 1680363874
transform 1 0 1172 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1680363874
transform 1 0 1204 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2799
timestamp 1680363874
transform 1 0 1204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1680363874
transform 1 0 1172 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1680363874
transform 1 0 1180 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1680363874
transform 1 0 1196 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2586
timestamp 1680363874
transform 1 0 1196 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1680363874
transform 1 0 1220 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2800
timestamp 1680363874
transform 1 0 1220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1680363874
transform 1 0 1220 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2455
timestamp 1680363874
transform 1 0 1332 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2801
timestamp 1680363874
transform 1 0 1260 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1680363874
transform 1 0 1324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1680363874
transform 1 0 1308 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2587
timestamp 1680363874
transform 1 0 1260 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1680363874
transform 1 0 1308 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2905
timestamp 1680363874
transform 1 0 1340 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1680363874
transform 1 0 1348 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2589
timestamp 1680363874
transform 1 0 1348 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1680363874
transform 1 0 1364 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1680363874
transform 1 0 1396 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1680363874
transform 1 0 1388 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1680363874
transform 1 0 1412 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1680363874
transform 1 0 1404 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2803
timestamp 1680363874
transform 1 0 1404 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1680363874
transform 1 0 1412 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2616
timestamp 1680363874
transform 1 0 1428 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1680363874
transform 1 0 1452 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2805
timestamp 1680363874
transform 1 0 1452 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1680363874
transform 1 0 1444 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2617
timestamp 1680363874
transform 1 0 1444 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1680363874
transform 1 0 1484 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2908
timestamp 1680363874
transform 1 0 1484 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2618
timestamp 1680363874
transform 1 0 1484 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1680363874
transform 1 0 1532 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1680363874
transform 1 0 1588 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2806
timestamp 1680363874
transform 1 0 1572 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1680363874
transform 1 0 1604 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1680363874
transform 1 0 1524 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2590
timestamp 1680363874
transform 1 0 1572 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2910
timestamp 1680363874
transform 1 0 1644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2477
timestamp 1680363874
transform 1 0 1660 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2808
timestamp 1680363874
transform 1 0 1660 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1680363874
transform 1 0 1676 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1680363874
transform 1 0 1668 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2591
timestamp 1680363874
transform 1 0 1668 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1680363874
transform 1 0 1668 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1680363874
transform 1 0 1692 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2912
timestamp 1680363874
transform 1 0 1708 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2621
timestamp 1680363874
transform 1 0 1708 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2775
timestamp 1680363874
transform 1 0 1748 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1680363874
transform 1 0 1732 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1680363874
transform 1 0 1724 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2622
timestamp 1680363874
transform 1 0 1732 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1680363874
transform 1 0 1780 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1680363874
transform 1 0 1780 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2914
timestamp 1680363874
transform 1 0 1780 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1680363874
transform 1 0 1796 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1680363874
transform 1 0 1796 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2550
timestamp 1680363874
transform 1 0 1820 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2975
timestamp 1680363874
transform 1 0 1812 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2488
timestamp 1680363874
transform 1 0 1844 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1680363874
transform 1 0 1852 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1680363874
transform 1 0 1868 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1680363874
transform 1 0 1916 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2812
timestamp 1680363874
transform 1 0 1860 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1680363874
transform 1 0 1916 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1680363874
transform 1 0 1956 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1680363874
transform 1 0 1940 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1680363874
transform 1 0 1956 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2592
timestamp 1680363874
transform 1 0 1860 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1680363874
transform 1 0 1956 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2815
timestamp 1680363874
transform 1 0 2004 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1680363874
transform 1 0 2004 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2478
timestamp 1680363874
transform 1 0 2044 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1680363874
transform 1 0 2028 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1680363874
transform 1 0 2028 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2816
timestamp 1680363874
transform 1 0 2020 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1680363874
transform 1 0 2020 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2919
timestamp 1680363874
transform 1 0 2028 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2566
timestamp 1680363874
transform 1 0 2036 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1680363874
transform 1 0 2052 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2920
timestamp 1680363874
transform 1 0 2044 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1680363874
transform 1 0 2060 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2521
timestamp 1680363874
transform 1 0 2084 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2817
timestamp 1680363874
transform 1 0 2076 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1680363874
transform 1 0 2108 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1680363874
transform 1 0 2100 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1680363874
transform 1 0 2148 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2819
timestamp 1680363874
transform 1 0 2196 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1680363874
transform 1 0 2148 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2567
timestamp 1680363874
transform 1 0 2212 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1680363874
transform 1 0 2196 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1680363874
transform 1 0 2196 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1680363874
transform 1 0 2236 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1680363874
transform 1 0 2236 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1680363874
transform 1 0 2252 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2923
timestamp 1680363874
transform 1 0 2276 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2491
timestamp 1680363874
transform 1 0 2308 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1680363874
transform 1 0 2292 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1680363874
transform 1 0 2316 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2820
timestamp 1680363874
transform 1 0 2292 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1680363874
transform 1 0 2300 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1680363874
transform 1 0 2316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1680363874
transform 1 0 2308 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2595
timestamp 1680363874
transform 1 0 2308 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1680363874
transform 1 0 2332 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2925
timestamp 1680363874
transform 1 0 2340 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2627
timestamp 1680363874
transform 1 0 2340 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2823
timestamp 1680363874
transform 1 0 2404 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1680363874
transform 1 0 2460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1680363874
transform 1 0 2380 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2596
timestamp 1680363874
transform 1 0 2380 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1680363874
transform 1 0 2396 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1680363874
transform 1 0 2484 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2927
timestamp 1680363874
transform 1 0 2508 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2493
timestamp 1680363874
transform 1 0 2524 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2825
timestamp 1680363874
transform 1 0 2532 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2568
timestamp 1680363874
transform 1 0 2532 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2928
timestamp 1680363874
transform 1 0 2540 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1680363874
transform 1 0 2564 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2569
timestamp 1680363874
transform 1 0 2596 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1680363874
transform 1 0 2636 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1680363874
transform 1 0 2620 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1680363874
transform 1 0 2612 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1680363874
transform 1 0 2636 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1680363874
transform 1 0 2612 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1680363874
transform 1 0 2620 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1680363874
transform 1 0 2636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1680363874
transform 1 0 2652 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1680363874
transform 1 0 2628 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1680363874
transform 1 0 2644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2597
timestamp 1680363874
transform 1 0 2620 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1680363874
transform 1 0 2612 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2932
timestamp 1680363874
transform 1 0 2660 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2598
timestamp 1680363874
transform 1 0 2652 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1680363874
transform 1 0 2644 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2830
timestamp 1680363874
transform 1 0 2732 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1680363874
transform 1 0 2724 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1680363874
transform 1 0 2740 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2632
timestamp 1680363874
transform 1 0 2716 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1680363874
transform 1 0 2740 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1680363874
transform 1 0 2756 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1680363874
transform 1 0 2772 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2935
timestamp 1680363874
transform 1 0 2780 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1680363874
transform 1 0 2796 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2527
timestamp 1680363874
transform 1 0 2820 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2832
timestamp 1680363874
transform 1 0 2820 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1680363874
transform 1 0 2812 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1680363874
transform 1 0 2836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1680363874
transform 1 0 2852 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1680363874
transform 1 0 2868 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1680363874
transform 1 0 2844 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1680363874
transform 1 0 2860 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2634
timestamp 1680363874
transform 1 0 2836 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1680363874
transform 1 0 2860 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2939
timestamp 1680363874
transform 1 0 2876 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1680363874
transform 1 0 2900 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1680363874
transform 1 0 2900 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2836
timestamp 1680363874
transform 1 0 2916 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1680363874
transform 1 0 2924 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2636
timestamp 1680363874
transform 1 0 2908 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1680363874
transform 1 0 2924 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1680363874
transform 1 0 2956 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2941
timestamp 1680363874
transform 1 0 2964 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2528
timestamp 1680363874
transform 1 0 2972 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2942
timestamp 1680363874
transform 1 0 2972 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2529
timestamp 1680363874
transform 1 0 2996 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2838
timestamp 1680363874
transform 1 0 2996 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2570
timestamp 1680363874
transform 1 0 3012 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1680363874
transform 1 0 3036 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2839
timestamp 1680363874
transform 1 0 3036 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1680363874
transform 1 0 3052 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2496
timestamp 1680363874
transform 1 0 3076 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2776
timestamp 1680363874
transform 1 0 3076 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2497
timestamp 1680363874
transform 1 0 3116 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2777
timestamp 1680363874
transform 1 0 3116 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1680363874
transform 1 0 3100 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1680363874
transform 1 0 3116 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1680363874
transform 1 0 3084 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1680363874
transform 1 0 3092 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2601
timestamp 1680363874
transform 1 0 3092 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1680363874
transform 1 0 3228 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1680363874
transform 1 0 3148 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1680363874
transform 1 0 3140 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1680363874
transform 1 0 3204 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2843
timestamp 1680363874
transform 1 0 3148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1680363874
transform 1 0 3204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1680363874
transform 1 0 3140 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1680363874
transform 1 0 3228 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2532
timestamp 1680363874
transform 1 0 3244 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2845
timestamp 1680363874
transform 1 0 3244 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1680363874
transform 1 0 3300 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2460
timestamp 1680363874
transform 1 0 3324 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1680363874
transform 1 0 3316 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2847
timestamp 1680363874
transform 1 0 3324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1680363874
transform 1 0 3308 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1680363874
transform 1 0 3316 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1680363874
transform 1 0 3332 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2499
timestamp 1680363874
transform 1 0 3348 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2778
timestamp 1680363874
transform 1 0 3348 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1680363874
transform 1 0 3364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1680363874
transform 1 0 3412 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1680363874
transform 1 0 3396 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2551
timestamp 1680363874
transform 1 0 3428 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1680363874
transform 1 0 3476 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1680363874
transform 1 0 3516 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2850
timestamp 1680363874
transform 1 0 3460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1680363874
transform 1 0 3492 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2552
timestamp 1680363874
transform 1 0 3540 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2951
timestamp 1680363874
transform 1 0 3540 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2602
timestamp 1680363874
transform 1 0 3540 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1680363874
transform 1 0 3564 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1680363874
transform 1 0 3572 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1680363874
transform 1 0 3564 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1680363874
transform 1 0 3564 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1680363874
transform 1 0 3588 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1680363874
transform 1 0 3580 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2852
timestamp 1680363874
transform 1 0 3588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1680363874
transform 1 0 3572 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2471
timestamp 1680363874
transform 1 0 3652 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1680363874
transform 1 0 3692 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1680363874
transform 1 0 3636 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2853
timestamp 1680363874
transform 1 0 3604 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1680363874
transform 1 0 3636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1680363874
transform 1 0 3684 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2603
timestamp 1680363874
transform 1 0 3684 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1680363874
transform 1 0 3708 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1680363874
transform 1 0 3796 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2855
timestamp 1680363874
transform 1 0 3708 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1680363874
transform 1 0 3764 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2554
timestamp 1680363874
transform 1 0 3788 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2954
timestamp 1680363874
transform 1 0 3788 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1680363874
transform 1 0 3804 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1680363874
transform 1 0 3836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1680363874
transform 1 0 3892 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2535
timestamp 1680363874
transform 1 0 3956 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2859
timestamp 1680363874
transform 1 0 3940 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1680363874
transform 1 0 3956 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1680363874
transform 1 0 3972 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1680363874
transform 1 0 3932 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1680363874
transform 1 0 3964 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2571
timestamp 1680363874
transform 1 0 3972 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2862
timestamp 1680363874
transform 1 0 3988 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1680363874
transform 1 0 3980 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2604
timestamp 1680363874
transform 1 0 3956 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1680363874
transform 1 0 3980 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1680363874
transform 1 0 3972 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1680363874
transform 1 0 3996 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1680363874
transform 1 0 4012 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1680363874
transform 1 0 4036 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2959
timestamp 1680363874
transform 1 0 4036 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2572
timestamp 1680363874
transform 1 0 4044 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2863
timestamp 1680363874
transform 1 0 4068 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1680363874
transform 1 0 4156 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1680363874
transform 1 0 4188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1680363874
transform 1 0 4108 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2606
timestamp 1680363874
transform 1 0 4188 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1680363874
transform 1 0 4148 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2961
timestamp 1680363874
transform 1 0 4204 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2556
timestamp 1680363874
transform 1 0 4220 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1680363874
transform 1 0 4236 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2866
timestamp 1680363874
transform 1 0 4236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1680363874
transform 1 0 4252 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1680363874
transform 1 0 4244 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2573
timestamp 1680363874
transform 1 0 4252 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2963
timestamp 1680363874
transform 1 0 4260 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2607
timestamp 1680363874
transform 1 0 4260 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1680363874
transform 1 0 4244 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1680363874
transform 1 0 4300 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2868
timestamp 1680363874
transform 1 0 4300 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1680363874
transform 1 0 4300 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1680363874
transform 1 0 4308 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1680363874
transform 1 0 4308 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1680363874
transform 1 0 4332 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1680363874
transform 1 0 4324 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2869
timestamp 1680363874
transform 1 0 4340 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1680363874
transform 1 0 4332 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2575
timestamp 1680363874
transform 1 0 4340 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2966
timestamp 1680363874
transform 1 0 4348 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1680363874
transform 1 0 4356 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2641
timestamp 1680363874
transform 1 0 4340 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1680363874
transform 1 0 4364 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2870
timestamp 1680363874
transform 1 0 4364 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2609
timestamp 1680363874
transform 1 0 4356 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1680363874
transform 1 0 4388 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2871
timestamp 1680363874
transform 1 0 4396 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2463
timestamp 1680363874
transform 1 0 4412 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1680363874
transform 1 0 4484 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2872
timestamp 1680363874
transform 1 0 4452 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2557
timestamp 1680363874
transform 1 0 4484 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1680363874
transform 1 0 4404 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1680363874
transform 1 0 4452 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2968
timestamp 1680363874
transform 1 0 4484 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2642
timestamp 1680363874
transform 1 0 4420 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1680363874
transform 1 0 4508 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2873
timestamp 1680363874
transform 1 0 4516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1680363874
transform 1 0 4532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1680363874
transform 1 0 4508 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1680363874
transform 1 0 4524 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1680363874
transform 1 0 4556 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2559
timestamp 1680363874
transform 1 0 4604 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2876
timestamp 1680363874
transform 1 0 4612 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2560
timestamp 1680363874
transform 1 0 4652 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2971
timestamp 1680363874
transform 1 0 4644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1680363874
transform 1 0 4636 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1680363874
transform 1 0 4700 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2877
timestamp 1680363874
transform 1 0 4684 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1680363874
transform 1 0 4692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1680363874
transform 1 0 4700 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1680363874
transform 1 0 4676 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1680363874
transform 1 0 4684 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2610
timestamp 1680363874
transform 1 0 4676 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1680363874
transform 1 0 4684 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1680363874
transform 1 0 4700 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1680363874
transform 1 0 4788 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1680363874
transform 1 0 4756 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2880
timestamp 1680363874
transform 1 0 4756 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1680363874
transform 1 0 4788 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2645
timestamp 1680363874
transform 1 0 4708 0 1 3385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_26
timestamp 1680363874
transform 1 0 48 0 1 3370
box -10 -3 10 3
use FILL  FILL_2552
timestamp 1680363874
transform 1 0 72 0 1 3370
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1680363874
transform 1 0 80 0 1 3370
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1680363874
transform 1 0 88 0 1 3370
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1680363874
transform 1 0 96 0 1 3370
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1680363874
transform 1 0 104 0 1 3370
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1680363874
transform 1 0 112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1680363874
transform 1 0 120 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_195
timestamp 1680363874
transform 1 0 128 0 1 3370
box -9 -3 26 105
use FILL  FILL_2560
timestamp 1680363874
transform 1 0 144 0 1 3370
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1680363874
transform 1 0 152 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_158
timestamp 1680363874
transform 1 0 160 0 1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2646
timestamp 1680363874
transform 1 0 212 0 1 3375
box -3 -3 3 3
use FILL  FILL_2562
timestamp 1680363874
transform 1 0 200 0 1 3370
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1680363874
transform 1 0 208 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2647
timestamp 1680363874
transform 1 0 276 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_194
timestamp 1680363874
transform 1 0 216 0 1 3370
box -8 -3 104 105
use FILL  FILL_2566
timestamp 1680363874
transform 1 0 312 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_196
timestamp 1680363874
transform 1 0 320 0 1 3370
box -9 -3 26 105
use FILL  FILL_2575
timestamp 1680363874
transform 1 0 336 0 1 3370
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1680363874
transform 1 0 344 0 1 3370
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1680363874
transform 1 0 352 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2648
timestamp 1680363874
transform 1 0 404 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_160
timestamp 1680363874
transform 1 0 360 0 1 3370
box -8 -3 46 105
use FILL  FILL_2581
timestamp 1680363874
transform 1 0 400 0 1 3370
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1680363874
transform 1 0 408 0 1 3370
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1680363874
transform 1 0 416 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_198
timestamp 1680363874
transform -1 0 440 0 1 3370
box -9 -3 26 105
use M3_M2  M3_M2_2649
timestamp 1680363874
transform 1 0 452 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_195
timestamp 1680363874
transform 1 0 440 0 1 3370
box -8 -3 104 105
use FILL  FILL_2590
timestamp 1680363874
transform 1 0 536 0 1 3370
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1680363874
transform 1 0 544 0 1 3370
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1680363874
transform 1 0 552 0 1 3370
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1680363874
transform 1 0 560 0 1 3370
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1680363874
transform 1 0 568 0 1 3370
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1680363874
transform 1 0 576 0 1 3370
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1680363874
transform 1 0 584 0 1 3370
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1680363874
transform 1 0 592 0 1 3370
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1680363874
transform 1 0 600 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_163
timestamp 1680363874
transform 1 0 608 0 1 3370
box -8 -3 46 105
use FILL  FILL_2612
timestamp 1680363874
transform 1 0 648 0 1 3370
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1680363874
transform 1 0 656 0 1 3370
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1680363874
transform 1 0 664 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1680363874
transform -1 0 696 0 1 3370
box -8 -3 32 105
use FILL  FILL_2617
timestamp 1680363874
transform 1 0 696 0 1 3370
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1680363874
transform 1 0 704 0 1 3370
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1680363874
transform 1 0 712 0 1 3370
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1680363874
transform 1 0 720 0 1 3370
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1680363874
transform 1 0 728 0 1 3370
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1680363874
transform 1 0 736 0 1 3370
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1680363874
transform 1 0 744 0 1 3370
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1680363874
transform 1 0 752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1680363874
transform 1 0 760 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_16
timestamp 1680363874
transform 1 0 768 0 1 3370
box -8 -3 32 105
use FILL  FILL_2634
timestamp 1680363874
transform 1 0 792 0 1 3370
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1680363874
transform 1 0 800 0 1 3370
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1680363874
transform 1 0 808 0 1 3370
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1680363874
transform 1 0 816 0 1 3370
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1680363874
transform 1 0 824 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_17
timestamp 1680363874
transform -1 0 856 0 1 3370
box -8 -3 32 105
use FILL  FILL_2642
timestamp 1680363874
transform 1 0 856 0 1 3370
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1680363874
transform 1 0 864 0 1 3370
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1680363874
transform 1 0 872 0 1 3370
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1680363874
transform 1 0 880 0 1 3370
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1680363874
transform 1 0 888 0 1 3370
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1680363874
transform 1 0 896 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_79
timestamp 1680363874
transform -1 0 936 0 1 3370
box -8 -3 34 105
use FILL  FILL_2654
timestamp 1680363874
transform 1 0 936 0 1 3370
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1680363874
transform 1 0 944 0 1 3370
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1680363874
transform 1 0 952 0 1 3370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1680363874
transform 1 0 960 0 1 3370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1680363874
transform 1 0 968 0 1 3370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1680363874
transform 1 0 976 0 1 3370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1680363874
transform 1 0 984 0 1 3370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1680363874
transform 1 0 992 0 1 3370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1680363874
transform 1 0 1000 0 1 3370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1680363874
transform 1 0 1008 0 1 3370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1680363874
transform 1 0 1016 0 1 3370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1680363874
transform 1 0 1024 0 1 3370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1680363874
transform 1 0 1032 0 1 3370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1680363874
transform 1 0 1040 0 1 3370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1680363874
transform 1 0 1048 0 1 3370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1680363874
transform 1 0 1056 0 1 3370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1680363874
transform 1 0 1064 0 1 3370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1680363874
transform 1 0 1072 0 1 3370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1680363874
transform 1 0 1080 0 1 3370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1680363874
transform 1 0 1088 0 1 3370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1680363874
transform 1 0 1096 0 1 3370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1680363874
transform 1 0 1104 0 1 3370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1680363874
transform 1 0 1112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1680363874
transform 1 0 1120 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_200
timestamp 1680363874
transform -1 0 1144 0 1 3370
box -9 -3 26 105
use FILL  FILL_2694
timestamp 1680363874
transform 1 0 1144 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2650
timestamp 1680363874
transform 1 0 1164 0 1 3375
box -3 -3 3 3
use FILL  FILL_2695
timestamp 1680363874
transform 1 0 1152 0 1 3370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1680363874
transform 1 0 1160 0 1 3370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1680363874
transform 1 0 1168 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_168
timestamp 1680363874
transform 1 0 1176 0 1 3370
box -8 -3 46 105
use FILL  FILL_2700
timestamp 1680363874
transform 1 0 1216 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2651
timestamp 1680363874
transform 1 0 1316 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_196
timestamp 1680363874
transform -1 0 1320 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_201
timestamp 1680363874
transform -1 0 1336 0 1 3370
box -9 -3 26 105
use FILL  FILL_2701
timestamp 1680363874
transform 1 0 1336 0 1 3370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1680363874
transform 1 0 1344 0 1 3370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1680363874
transform 1 0 1352 0 1 3370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1680363874
transform 1 0 1360 0 1 3370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1680363874
transform 1 0 1368 0 1 3370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1680363874
transform 1 0 1376 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_2
timestamp 1680363874
transform -1 0 1408 0 1 3370
box -5 -3 28 105
use FILL  FILL_2707
timestamp 1680363874
transform 1 0 1408 0 1 3370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1680363874
transform 1 0 1416 0 1 3370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1680363874
transform 1 0 1424 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_202
timestamp 1680363874
transform -1 0 1448 0 1 3370
box -9 -3 26 105
use FILL  FILL_2710
timestamp 1680363874
transform 1 0 1448 0 1 3370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1680363874
transform 1 0 1456 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_3
timestamp 1680363874
transform 1 0 1464 0 1 3370
box -5 -3 28 105
use FILL  FILL_2712
timestamp 1680363874
transform 1 0 1488 0 1 3370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1680363874
transform 1 0 1496 0 1 3370
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1680363874
transform 1 0 1504 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2652
timestamp 1680363874
transform 1 0 1548 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_197
timestamp 1680363874
transform 1 0 1512 0 1 3370
box -8 -3 104 105
use FILL  FILL_2715
timestamp 1680363874
transform 1 0 1608 0 1 3370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1680363874
transform 1 0 1616 0 1 3370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1680363874
transform 1 0 1624 0 1 3370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1680363874
transform 1 0 1632 0 1 3370
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1680363874
transform 1 0 1640 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_169
timestamp 1680363874
transform -1 0 1688 0 1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2653
timestamp 1680363874
transform 1 0 1700 0 1 3375
box -3 -3 3 3
use FILL  FILL_2720
timestamp 1680363874
transform 1 0 1688 0 1 3370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1680363874
transform 1 0 1696 0 1 3370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1680363874
transform 1 0 1704 0 1 3370
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1680363874
transform 1 0 1712 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_81
timestamp 1680363874
transform 1 0 1720 0 1 3370
box -8 -3 34 105
use FILL  FILL_2746
timestamp 1680363874
transform 1 0 1752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1680363874
transform 1 0 1760 0 1 3370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1680363874
transform 1 0 1768 0 1 3370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1680363874
transform 1 0 1776 0 1 3370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1680363874
transform 1 0 1784 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_26
timestamp 1680363874
transform -1 0 1816 0 1 3370
box -8 -3 32 105
use FILL  FILL_2757
timestamp 1680363874
transform 1 0 1816 0 1 3370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1680363874
transform 1 0 1824 0 1 3370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1680363874
transform 1 0 1832 0 1 3370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1680363874
transform 1 0 1840 0 1 3370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1680363874
transform 1 0 1848 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_200
timestamp 1680363874
transform -1 0 1952 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_206
timestamp 1680363874
transform 1 0 1952 0 1 3370
box -9 -3 26 105
use FILL  FILL_2766
timestamp 1680363874
transform 1 0 1968 0 1 3370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1680363874
transform 1 0 1976 0 1 3370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1680363874
transform 1 0 1984 0 1 3370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1680363874
transform 1 0 1992 0 1 3370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1680363874
transform 1 0 2000 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2654
timestamp 1680363874
transform 1 0 2052 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_173
timestamp 1680363874
transform -1 0 2048 0 1 3370
box -8 -3 46 105
use FILL  FILL_2771
timestamp 1680363874
transform 1 0 2048 0 1 3370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1680363874
transform 1 0 2056 0 1 3370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1680363874
transform 1 0 2064 0 1 3370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1680363874
transform 1 0 2072 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2655
timestamp 1680363874
transform 1 0 2092 0 1 3375
box -3 -3 3 3
use FILL  FILL_2792
timestamp 1680363874
transform 1 0 2080 0 1 3370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1680363874
transform 1 0 2088 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_209
timestamp 1680363874
transform 1 0 2096 0 1 3370
box -9 -3 26 105
use FILL  FILL_2794
timestamp 1680363874
transform 1 0 2112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1680363874
transform 1 0 2120 0 1 3370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1680363874
transform 1 0 2128 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1680363874
transform 1 0 2136 0 1 3370
box -8 -3 104 105
use FILL  FILL_2797
timestamp 1680363874
transform 1 0 2232 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_210
timestamp 1680363874
transform 1 0 2240 0 1 3370
box -9 -3 26 105
use FILL  FILL_2798
timestamp 1680363874
transform 1 0 2256 0 1 3370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1680363874
transform 1 0 2264 0 1 3370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1680363874
transform 1 0 2272 0 1 3370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1680363874
transform 1 0 2280 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_176
timestamp 1680363874
transform 1 0 2288 0 1 3370
box -8 -3 46 105
use FILL  FILL_2811
timestamp 1680363874
transform 1 0 2328 0 1 3370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1680363874
transform 1 0 2336 0 1 3370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1680363874
transform 1 0 2344 0 1 3370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1680363874
transform 1 0 2352 0 1 3370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1680363874
transform 1 0 2360 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2656
timestamp 1680363874
transform 1 0 2380 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1680363874
transform 1 0 2404 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_203
timestamp 1680363874
transform 1 0 2368 0 1 3370
box -8 -3 104 105
use FILL  FILL_2826
timestamp 1680363874
transform 1 0 2464 0 1 3370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1680363874
transform 1 0 2472 0 1 3370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1680363874
transform 1 0 2480 0 1 3370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1680363874
transform 1 0 2488 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2658
timestamp 1680363874
transform 1 0 2508 0 1 3375
box -3 -3 3 3
use FILL  FILL_2830
timestamp 1680363874
transform 1 0 2496 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2659
timestamp 1680363874
transform 1 0 2532 0 1 3375
box -3 -3 3 3
use INVX2  INVX2_212
timestamp 1680363874
transform 1 0 2504 0 1 3370
box -9 -3 26 105
use FILL  FILL_2831
timestamp 1680363874
transform 1 0 2520 0 1 3370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1680363874
transform 1 0 2528 0 1 3370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1680363874
transform 1 0 2536 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_213
timestamp 1680363874
transform 1 0 2544 0 1 3370
box -9 -3 26 105
use FILL  FILL_2840
timestamp 1680363874
transform 1 0 2560 0 1 3370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1680363874
transform 1 0 2568 0 1 3370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1680363874
transform 1 0 2576 0 1 3370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1680363874
transform 1 0 2584 0 1 3370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1680363874
transform 1 0 2592 0 1 3370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1680363874
transform 1 0 2600 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_178
timestamp 1680363874
transform 1 0 2608 0 1 3370
box -8 -3 46 105
use FILL  FILL_2849
timestamp 1680363874
transform 1 0 2648 0 1 3370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1680363874
transform 1 0 2656 0 1 3370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1680363874
transform 1 0 2664 0 1 3370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1680363874
transform 1 0 2672 0 1 3370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1680363874
transform 1 0 2680 0 1 3370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1680363874
transform 1 0 2688 0 1 3370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1680363874
transform 1 0 2696 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_180
timestamp 1680363874
transform 1 0 2704 0 1 3370
box -8 -3 46 105
use FILL  FILL_2864
timestamp 1680363874
transform 1 0 2744 0 1 3370
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1680363874
transform 1 0 2752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1680363874
transform 1 0 2760 0 1 3370
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1680363874
transform 1 0 2768 0 1 3370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1680363874
transform 1 0 2776 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_214
timestamp 1680363874
transform 1 0 2784 0 1 3370
box -9 -3 26 105
use FILL  FILL_2871
timestamp 1680363874
transform 1 0 2800 0 1 3370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1680363874
transform 1 0 2808 0 1 3370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1680363874
transform 1 0 2816 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_181
timestamp 1680363874
transform 1 0 2824 0 1 3370
box -8 -3 46 105
use FILL  FILL_2874
timestamp 1680363874
transform 1 0 2864 0 1 3370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1680363874
transform 1 0 2872 0 1 3370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1680363874
transform 1 0 2880 0 1 3370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1680363874
transform 1 0 2888 0 1 3370
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1680363874
transform 1 0 2896 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_215
timestamp 1680363874
transform 1 0 2904 0 1 3370
box -9 -3 26 105
use FILL  FILL_2885
timestamp 1680363874
transform 1 0 2920 0 1 3370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1680363874
transform 1 0 2928 0 1 3370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1680363874
transform 1 0 2936 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_216
timestamp 1680363874
transform -1 0 2960 0 1 3370
box -9 -3 26 105
use FILL  FILL_2891
timestamp 1680363874
transform 1 0 2960 0 1 3370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1680363874
transform 1 0 2968 0 1 3370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1680363874
transform 1 0 2976 0 1 3370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1680363874
transform 1 0 2984 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_83
timestamp 1680363874
transform 1 0 2992 0 1 3370
box -8 -3 34 105
use FILL  FILL_2895
timestamp 1680363874
transform 1 0 3024 0 1 3370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1680363874
transform 1 0 3032 0 1 3370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1680363874
transform 1 0 3040 0 1 3370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1680363874
transform 1 0 3048 0 1 3370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1680363874
transform 1 0 3056 0 1 3370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1680363874
transform 1 0 3064 0 1 3370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1680363874
transform 1 0 3072 0 1 3370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1680363874
transform 1 0 3080 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_84
timestamp 1680363874
transform 1 0 3088 0 1 3370
box -8 -3 34 105
use FILL  FILL_2910
timestamp 1680363874
transform 1 0 3120 0 1 3370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1680363874
transform 1 0 3128 0 1 3370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1680363874
transform 1 0 3136 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_207
timestamp 1680363874
transform -1 0 3240 0 1 3370
box -8 -3 104 105
use FILL  FILL_2918
timestamp 1680363874
transform 1 0 3240 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_217
timestamp 1680363874
transform -1 0 3264 0 1 3370
box -9 -3 26 105
use FILL  FILL_2919
timestamp 1680363874
transform 1 0 3264 0 1 3370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1680363874
transform 1 0 3272 0 1 3370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1680363874
transform 1 0 3280 0 1 3370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1680363874
transform 1 0 3288 0 1 3370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1680363874
transform 1 0 3296 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_118
timestamp 1680363874
transform -1 0 3344 0 1 3370
box -8 -3 46 105
use FILL  FILL_2936
timestamp 1680363874
transform 1 0 3344 0 1 3370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1680363874
transform 1 0 3352 0 1 3370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1680363874
transform 1 0 3360 0 1 3370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1680363874
transform 1 0 3368 0 1 3370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1680363874
transform 1 0 3376 0 1 3370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1680363874
transform 1 0 3384 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_87
timestamp 1680363874
transform -1 0 3424 0 1 3370
box -8 -3 34 105
use FILL  FILL_2947
timestamp 1680363874
transform 1 0 3424 0 1 3370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1680363874
transform 1 0 3432 0 1 3370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1680363874
transform 1 0 3440 0 1 3370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1680363874
transform 1 0 3448 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_208
timestamp 1680363874
transform -1 0 3552 0 1 3370
box -8 -3 104 105
use FILL  FILL_2951
timestamp 1680363874
transform 1 0 3552 0 1 3370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1680363874
transform 1 0 3560 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_219
timestamp 1680363874
transform 1 0 3568 0 1 3370
box -9 -3 26 105
use FILL  FILL_2953
timestamp 1680363874
transform 1 0 3584 0 1 3370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1680363874
transform 1 0 3592 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1680363874
transform -1 0 3696 0 1 3370
box -8 -3 104 105
use FILL  FILL_2965
timestamp 1680363874
transform 1 0 3696 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1680363874
transform -1 0 3800 0 1 3370
box -8 -3 104 105
use FILL  FILL_2966
timestamp 1680363874
transform 1 0 3800 0 1 3370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1680363874
transform 1 0 3808 0 1 3370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1680363874
transform 1 0 3816 0 1 3370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1680363874
transform 1 0 3824 0 1 3370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1680363874
transform 1 0 3832 0 1 3370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1680363874
transform 1 0 3840 0 1 3370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1680363874
transform 1 0 3848 0 1 3370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1680363874
transform 1 0 3856 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2660
timestamp 1680363874
transform 1 0 3876 0 1 3375
box -3 -3 3 3
use FILL  FILL_2995
timestamp 1680363874
transform 1 0 3864 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_220
timestamp 1680363874
transform 1 0 3872 0 1 3370
box -9 -3 26 105
use FILL  FILL_2997
timestamp 1680363874
transform 1 0 3888 0 1 3370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1680363874
transform 1 0 3896 0 1 3370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1680363874
transform 1 0 3904 0 1 3370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1680363874
transform 1 0 3912 0 1 3370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1680363874
transform 1 0 3920 0 1 3370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1680363874
transform 1 0 3928 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_122
timestamp 1680363874
transform -1 0 3976 0 1 3370
box -8 -3 46 105
use FILL  FILL_3009
timestamp 1680363874
transform 1 0 3976 0 1 3370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1680363874
transform 1 0 3984 0 1 3370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1680363874
transform 1 0 3992 0 1 3370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1680363874
transform 1 0 4000 0 1 3370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1680363874
transform 1 0 4008 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_221
timestamp 1680363874
transform 1 0 4016 0 1 3370
box -9 -3 26 105
use FILL  FILL_3014
timestamp 1680363874
transform 1 0 4032 0 1 3370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1680363874
transform 1 0 4040 0 1 3370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1680363874
transform 1 0 4048 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_222
timestamp 1680363874
transform 1 0 4056 0 1 3370
box -9 -3 26 105
use FILL  FILL_3022
timestamp 1680363874
transform 1 0 4072 0 1 3370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1680363874
transform 1 0 4080 0 1 3370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1680363874
transform 1 0 4088 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2661
timestamp 1680363874
transform 1 0 4108 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_213
timestamp 1680363874
transform 1 0 4096 0 1 3370
box -8 -3 104 105
use FILL  FILL_3025
timestamp 1680363874
transform 1 0 4192 0 1 3370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1680363874
transform 1 0 4200 0 1 3370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1680363874
transform 1 0 4208 0 1 3370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1680363874
transform 1 0 4216 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_184
timestamp 1680363874
transform 1 0 4224 0 1 3370
box -8 -3 46 105
use FILL  FILL_3029
timestamp 1680363874
transform 1 0 4264 0 1 3370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1680363874
transform 1 0 4272 0 1 3370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1680363874
transform 1 0 4280 0 1 3370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1680363874
transform 1 0 4288 0 1 3370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1680363874
transform 1 0 4296 0 1 3370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1680363874
transform 1 0 4304 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_185
timestamp 1680363874
transform 1 0 4312 0 1 3370
box -8 -3 46 105
use FILL  FILL_3044
timestamp 1680363874
transform 1 0 4352 0 1 3370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1680363874
transform 1 0 4360 0 1 3370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1680363874
transform 1 0 4368 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_224
timestamp 1680363874
transform 1 0 4376 0 1 3370
box -9 -3 26 105
use FILL  FILL_3053
timestamp 1680363874
transform 1 0 4392 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2662
timestamp 1680363874
transform 1 0 4492 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_215
timestamp 1680363874
transform -1 0 4496 0 1 3370
box -8 -3 104 105
use FILL  FILL_3054
timestamp 1680363874
transform 1 0 4496 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2663
timestamp 1680363874
transform 1 0 4516 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_186
timestamp 1680363874
transform 1 0 4504 0 1 3370
box -8 -3 46 105
use FILL  FILL_3055
timestamp 1680363874
transform 1 0 4544 0 1 3370
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1680363874
transform 1 0 4552 0 1 3370
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1680363874
transform 1 0 4560 0 1 3370
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1680363874
transform 1 0 4568 0 1 3370
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1680363874
transform 1 0 4576 0 1 3370
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1680363874
transform 1 0 4584 0 1 3370
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1680363874
transform 1 0 4592 0 1 3370
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1680363874
transform 1 0 4600 0 1 3370
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1680363874
transform 1 0 4608 0 1 3370
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1680363874
transform 1 0 4616 0 1 3370
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1680363874
transform 1 0 4624 0 1 3370
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1680363874
transform 1 0 4632 0 1 3370
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1680363874
transform 1 0 4640 0 1 3370
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1680363874
transform 1 0 4648 0 1 3370
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1680363874
transform 1 0 4656 0 1 3370
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1680363874
transform 1 0 4664 0 1 3370
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1680363874
transform 1 0 4672 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1680363874
transform 1 0 4680 0 1 3370
box -9 -3 26 105
use FILL  FILL_3084
timestamp 1680363874
transform 1 0 4696 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_217
timestamp 1680363874
transform -1 0 4800 0 1 3370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_27
timestamp 1680363874
transform 1 0 4827 0 1 3370
box -10 -3 10 3
use M3_M2  M3_M2_2704
timestamp 1680363874
transform 1 0 140 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2977
timestamp 1680363874
transform 1 0 92 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1680363874
transform 1 0 180 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1680363874
transform 1 0 196 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1680363874
transform 1 0 140 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1680363874
transform 1 0 172 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1680363874
transform 1 0 188 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2830
timestamp 1680363874
transform 1 0 148 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1680363874
transform 1 0 196 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3083
timestamp 1680363874
transform 1 0 212 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2831
timestamp 1680363874
transform 1 0 204 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3189
timestamp 1680363874
transform 1 0 220 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2705
timestamp 1680363874
transform 1 0 260 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2980
timestamp 1680363874
transform 1 0 244 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1680363874
transform 1 0 260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1680363874
transform 1 0 276 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1680363874
transform 1 0 252 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1680363874
transform 1 0 268 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2782
timestamp 1680363874
transform 1 0 252 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1680363874
transform 1 0 268 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1680363874
transform 1 0 308 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2983
timestamp 1680363874
transform 1 0 316 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2677
timestamp 1680363874
transform 1 0 364 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1680363874
transform 1 0 356 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3086
timestamp 1680363874
transform 1 0 356 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1680363874
transform 1 0 412 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2678
timestamp 1680363874
transform 1 0 452 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2985
timestamp 1680363874
transform 1 0 436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1680363874
transform 1 0 452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1680363874
transform 1 0 428 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2816
timestamp 1680363874
transform 1 0 428 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2987
timestamp 1680363874
transform 1 0 532 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1680363874
transform 1 0 564 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2743
timestamp 1680363874
transform 1 0 572 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1680363874
transform 1 0 588 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2989
timestamp 1680363874
transform 1 0 580 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1680363874
transform 1 0 588 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1680363874
transform 1 0 548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1680363874
transform 1 0 556 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2762
timestamp 1680363874
transform 1 0 564 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3090
timestamp 1680363874
transform 1 0 572 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2783
timestamp 1680363874
transform 1 0 580 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1680363874
transform 1 0 580 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1680363874
transform 1 0 596 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1680363874
transform 1 0 652 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1680363874
transform 1 0 636 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2991
timestamp 1680363874
transform 1 0 636 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2744
timestamp 1680363874
transform 1 0 644 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1680363874
transform 1 0 660 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2992
timestamp 1680363874
transform 1 0 652 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1680363874
transform 1 0 660 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1680363874
transform 1 0 620 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1680363874
transform 1 0 644 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2784
timestamp 1680363874
transform 1 0 644 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3093
timestamp 1680363874
transform 1 0 660 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1680363874
transform 1 0 676 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2832
timestamp 1680363874
transform 1 0 676 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1680363874
transform 1 0 692 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1680363874
transform 1 0 732 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1680363874
transform 1 0 716 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1680363874
transform 1 0 740 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2994
timestamp 1680363874
transform 1 0 716 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1680363874
transform 1 0 732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1680363874
transform 1 0 740 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1680363874
transform 1 0 724 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2786
timestamp 1680363874
transform 1 0 716 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1680363874
transform 1 0 788 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3096
timestamp 1680363874
transform 1 0 788 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1680363874
transform 1 0 804 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1680363874
transform 1 0 812 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2818
timestamp 1680363874
transform 1 0 812 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1680363874
transform 1 0 844 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1680363874
transform 1 0 860 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3098
timestamp 1680363874
transform 1 0 868 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1680363874
transform 1 0 860 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2826
timestamp 1680363874
transform 1 0 868 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3192
timestamp 1680363874
transform 1 0 908 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1680363874
transform 1 0 940 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2680
timestamp 1680363874
transform 1 0 996 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2997
timestamp 1680363874
transform 1 0 996 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2763
timestamp 1680363874
transform 1 0 996 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1680363874
transform 1 0 988 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1680363874
transform 1 0 1036 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1680363874
transform 1 0 1060 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2998
timestamp 1680363874
transform 1 0 1044 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2746
timestamp 1680363874
transform 1 0 1052 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2999
timestamp 1680363874
transform 1 0 1060 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1680363874
transform 1 0 1036 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2788
timestamp 1680363874
transform 1 0 1028 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1680363874
transform 1 0 1044 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3100
timestamp 1680363874
transform 1 0 1052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1680363874
transform 1 0 1068 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2789
timestamp 1680363874
transform 1 0 1052 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1680363874
transform 1 0 1084 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3102
timestamp 1680363874
transform 1 0 1084 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2683
timestamp 1680363874
transform 1 0 1116 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1680363874
transform 1 0 1156 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1680363874
transform 1 0 1140 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3000
timestamp 1680363874
transform 1 0 1116 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1680363874
transform 1 0 1124 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1680363874
transform 1 0 1140 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1680363874
transform 1 0 1156 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1680363874
transform 1 0 1164 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1680363874
transform 1 0 1116 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2765
timestamp 1680363874
transform 1 0 1124 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3104
timestamp 1680363874
transform 1 0 1148 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2833
timestamp 1680363874
transform 1 0 1132 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1680363874
transform 1 0 1180 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1680363874
transform 1 0 1212 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1680363874
transform 1 0 1228 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3005
timestamp 1680363874
transform 1 0 1220 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1680363874
transform 1 0 1228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1680363874
transform 1 0 1212 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2766
timestamp 1680363874
transform 1 0 1220 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3106
timestamp 1680363874
transform 1 0 1228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1680363874
transform 1 0 1244 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2666
timestamp 1680363874
transform 1 0 1276 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1680363874
transform 1 0 1268 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3107
timestamp 1680363874
transform 1 0 1268 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2717
timestamp 1680363874
transform 1 0 1292 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3008
timestamp 1680363874
transform 1 0 1292 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1680363874
transform 1 0 1300 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2686
timestamp 1680363874
transform 1 0 1324 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3009
timestamp 1680363874
transform 1 0 1332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1680363874
transform 1 0 1340 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1680363874
transform 1 0 1380 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1680363874
transform 1 0 1404 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3010
timestamp 1680363874
transform 1 0 1428 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1680363874
transform 1 0 1380 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1680363874
transform 1 0 1428 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1680363874
transform 1 0 1516 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1680363874
transform 1 0 1476 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1680363874
transform 1 0 1492 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3011
timestamp 1680363874
transform 1 0 1540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1680363874
transform 1 0 1460 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1680363874
transform 1 0 1516 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2790
timestamp 1680363874
transform 1 0 1460 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3012
timestamp 1680363874
transform 1 0 1556 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2791
timestamp 1680363874
transform 1 0 1556 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1680363874
transform 1 0 1604 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_3113
timestamp 1680363874
transform 1 0 1596 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1680363874
transform 1 0 1604 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2720
timestamp 1680363874
transform 1 0 1628 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1680363874
transform 1 0 1644 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3014
timestamp 1680363874
transform 1 0 1628 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1680363874
transform 1 0 1644 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1680363874
transform 1 0 1612 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1680363874
transform 1 0 1620 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1680363874
transform 1 0 1636 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2792
timestamp 1680363874
transform 1 0 1612 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1680363874
transform 1 0 1636 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1680363874
transform 1 0 1620 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_3117
timestamp 1680363874
transform 1 0 1652 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2820
timestamp 1680363874
transform 1 0 1652 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1680363874
transform 1 0 1652 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1680363874
transform 1 0 1708 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1680363874
transform 1 0 1676 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1680363874
transform 1 0 1692 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1680363874
transform 1 0 1708 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1680363874
transform 1 0 1684 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1680363874
transform 1 0 1700 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2835
timestamp 1680363874
transform 1 0 1676 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3120
timestamp 1680363874
transform 1 0 1716 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2821
timestamp 1680363874
transform 1 0 1708 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_3019
timestamp 1680363874
transform 1 0 1748 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1680363874
transform 1 0 1756 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1680363874
transform 1 0 1788 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1680363874
transform 1 0 1828 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1680363874
transform 1 0 1844 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1680363874
transform 1 0 1852 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1680363874
transform 1 0 1876 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1680363874
transform 1 0 1884 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1680363874
transform 1 0 1948 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1680363874
transform 1 0 1964 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1680363874
transform 1 0 1980 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1680363874
transform 1 0 1988 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2794
timestamp 1680363874
transform 1 0 1988 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3025
timestamp 1680363874
transform 1 0 2004 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1680363874
transform 1 0 2004 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2795
timestamp 1680363874
transform 1 0 2004 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3026
timestamp 1680363874
transform 1 0 2044 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1680363874
transform 1 0 2052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1680363874
transform 1 0 2060 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1680363874
transform 1 0 2148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1680363874
transform 1 0 2100 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2768
timestamp 1680363874
transform 1 0 2148 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1680363874
transform 1 0 2076 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3130
timestamp 1680363874
transform 1 0 2164 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2797
timestamp 1680363874
transform 1 0 2164 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1680363874
transform 1 0 2204 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3028
timestamp 1680363874
transform 1 0 2204 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1680363874
transform 1 0 2220 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2769
timestamp 1680363874
transform 1 0 2212 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3131
timestamp 1680363874
transform 1 0 2228 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2687
timestamp 1680363874
transform 1 0 2244 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3132
timestamp 1680363874
transform 1 0 2244 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1680363874
transform 1 0 2252 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2751
timestamp 1680363874
transform 1 0 2276 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3031
timestamp 1680363874
transform 1 0 2292 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1680363874
transform 1 0 2284 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2688
timestamp 1680363874
transform 1 0 2300 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1680363874
transform 1 0 2316 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_3134
timestamp 1680363874
transform 1 0 2308 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2798
timestamp 1680363874
transform 1 0 2308 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3135
timestamp 1680363874
transform 1 0 2332 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2836
timestamp 1680363874
transform 1 0 2332 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1680363874
transform 1 0 2356 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3032
timestamp 1680363874
transform 1 0 2356 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2770
timestamp 1680363874
transform 1 0 2356 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1680363874
transform 1 0 2388 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3033
timestamp 1680363874
transform 1 0 2380 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1680363874
transform 1 0 2396 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1680363874
transform 1 0 2388 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2724
timestamp 1680363874
transform 1 0 2484 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1680363874
transform 1 0 2500 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3035
timestamp 1680363874
transform 1 0 2452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1680363874
transform 1 0 2540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1680363874
transform 1 0 2500 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1680363874
transform 1 0 2532 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2799
timestamp 1680363874
transform 1 0 2484 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1680363874
transform 1 0 2516 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1680363874
transform 1 0 2564 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1680363874
transform 1 0 2580 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1680363874
transform 1 0 2588 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3037
timestamp 1680363874
transform 1 0 2588 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1680363874
transform 1 0 2580 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1680363874
transform 1 0 2596 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2692
timestamp 1680363874
transform 1 0 2620 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1680363874
transform 1 0 2628 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3038
timestamp 1680363874
transform 1 0 2644 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2771
timestamp 1680363874
transform 1 0 2660 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1680363874
transform 1 0 2732 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3039
timestamp 1680363874
transform 1 0 2684 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1680363874
transform 1 0 2732 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2838
timestamp 1680363874
transform 1 0 2740 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3040
timestamp 1680363874
transform 1 0 2772 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2693
timestamp 1680363874
transform 1 0 2788 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3142
timestamp 1680363874
transform 1 0 2780 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2800
timestamp 1680363874
transform 1 0 2772 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1680363874
transform 1 0 2796 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1680363874
transform 1 0 2820 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1680363874
transform 1 0 2812 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3041
timestamp 1680363874
transform 1 0 2820 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1680363874
transform 1 0 2836 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1680363874
transform 1 0 2812 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2773
timestamp 1680363874
transform 1 0 2820 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3144
timestamp 1680363874
transform 1 0 2828 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2801
timestamp 1680363874
transform 1 0 2812 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3145
timestamp 1680363874
transform 1 0 2844 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1680363874
transform 1 0 2852 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2802
timestamp 1680363874
transform 1 0 2844 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1680363874
transform 1 0 2884 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1680363874
transform 1 0 2892 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1680363874
transform 1 0 2892 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3044
timestamp 1680363874
transform 1 0 2892 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1680363874
transform 1 0 2908 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1680363874
transform 1 0 2900 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1680363874
transform 1 0 2964 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2695
timestamp 1680363874
transform 1 0 3052 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1680363874
transform 1 0 3012 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3046
timestamp 1680363874
transform 1 0 3052 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1680363874
transform 1 0 3012 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2774
timestamp 1680363874
transform 1 0 3052 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3047
timestamp 1680363874
transform 1 0 3068 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2839
timestamp 1680363874
transform 1 0 3068 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3149
timestamp 1680363874
transform 1 0 3092 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1680363874
transform 1 0 3100 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2775
timestamp 1680363874
transform 1 0 3116 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3195
timestamp 1680363874
transform 1 0 3156 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1680363874
transform 1 0 3212 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2827
timestamp 1680363874
transform 1 0 3220 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3151
timestamp 1680363874
transform 1 0 3252 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2696
timestamp 1680363874
transform 1 0 3260 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1680363874
transform 1 0 3260 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3049
timestamp 1680363874
transform 1 0 3260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1680363874
transform 1 0 3268 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2803
timestamp 1680363874
transform 1 0 3268 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1680363874
transform 1 0 3292 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1680363874
transform 1 0 3284 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3051
timestamp 1680363874
transform 1 0 3284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1680363874
transform 1 0 3332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1680363874
transform 1 0 3300 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1680363874
transform 1 0 3308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1680363874
transform 1 0 3324 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2822
timestamp 1680363874
transform 1 0 3300 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1680363874
transform 1 0 3324 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1680363874
transform 1 0 3452 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1680363874
transform 1 0 3396 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1680363874
transform 1 0 3388 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3155
timestamp 1680363874
transform 1 0 3380 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1680363874
transform 1 0 3388 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2828
timestamp 1680363874
transform 1 0 3372 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3053
timestamp 1680363874
transform 1 0 3476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1680363874
transform 1 0 3428 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2823
timestamp 1680363874
transform 1 0 3428 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1680363874
transform 1 0 3428 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3054
timestamp 1680363874
transform 1 0 3508 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1680363874
transform 1 0 3556 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1680363874
transform 1 0 3604 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2805
timestamp 1680363874
transform 1 0 3604 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3160
timestamp 1680363874
transform 1 0 3620 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2734
timestamp 1680363874
transform 1 0 3636 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3055
timestamp 1680363874
transform 1 0 3636 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2755
timestamp 1680363874
transform 1 0 3644 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3056
timestamp 1680363874
transform 1 0 3652 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1680363874
transform 1 0 3644 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2776
timestamp 1680363874
transform 1 0 3652 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1680363874
transform 1 0 3676 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1680363874
transform 1 0 3668 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3162
timestamp 1680363874
transform 1 0 3660 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2840
timestamp 1680363874
transform 1 0 3644 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1680363874
transform 1 0 3660 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3163
timestamp 1680363874
transform 1 0 3676 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1680363874
transform 1 0 3692 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1680363874
transform 1 0 3748 0 1 3345
box -2 -2 2 2
use M3_M2  M3_M2_2671
timestamp 1680363874
transform 1 0 3812 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1680363874
transform 1 0 3812 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1680363874
transform 1 0 3788 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3058
timestamp 1680363874
transform 1 0 3788 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1680363874
transform 1 0 3796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1680363874
transform 1 0 3812 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1680363874
transform 1 0 3804 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1680363874
transform 1 0 3820 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2806
timestamp 1680363874
transform 1 0 3812 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1680363874
transform 1 0 3892 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1680363874
transform 1 0 3884 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1680363874
transform 1 0 4012 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1680363874
transform 1 0 3964 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1680363874
transform 1 0 3964 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3061
timestamp 1680363874
transform 1 0 4012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1680363874
transform 1 0 3932 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1680363874
transform 1 0 3988 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2842
timestamp 1680363874
transform 1 0 4004 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1680363874
transform 1 0 4028 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3168
timestamp 1680363874
transform 1 0 4044 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2738
timestamp 1680363874
transform 1 0 4084 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3062
timestamp 1680363874
transform 1 0 4084 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1680363874
transform 1 0 4100 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1680363874
transform 1 0 4108 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1680363874
transform 1 0 4092 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2739
timestamp 1680363874
transform 1 0 4132 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3170
timestamp 1680363874
transform 1 0 4132 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2807
timestamp 1680363874
transform 1 0 4132 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3171
timestamp 1680363874
transform 1 0 4148 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2673
timestamp 1680363874
transform 1 0 4220 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1680363874
transform 1 0 4220 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3065
timestamp 1680363874
transform 1 0 4172 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2758
timestamp 1680363874
transform 1 0 4212 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3172
timestamp 1680363874
transform 1 0 4212 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2674
timestamp 1680363874
transform 1 0 4316 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1680363874
transform 1 0 4316 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3066
timestamp 1680363874
transform 1 0 4300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1680363874
transform 1 0 4316 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1680363874
transform 1 0 4324 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1680363874
transform 1 0 4292 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1680363874
transform 1 0 4308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1680363874
transform 1 0 4324 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2808
timestamp 1680363874
transform 1 0 4292 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1680363874
transform 1 0 4348 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1680363874
transform 1 0 4364 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3069
timestamp 1680363874
transform 1 0 4372 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2809
timestamp 1680363874
transform 1 0 4372 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1680363874
transform 1 0 4404 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1680363874
transform 1 0 4396 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_3070
timestamp 1680363874
transform 1 0 4404 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1680363874
transform 1 0 4396 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2676
timestamp 1680363874
transform 1 0 4436 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_3071
timestamp 1680363874
transform 1 0 4420 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1680363874
transform 1 0 4436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1680363874
transform 1 0 4412 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2777
timestamp 1680363874
transform 1 0 4420 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3178
timestamp 1680363874
transform 1 0 4428 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1680363874
transform 1 0 4444 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2810
timestamp 1680363874
transform 1 0 4428 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1680363874
transform 1 0 4444 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_3073
timestamp 1680363874
transform 1 0 4484 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2703
timestamp 1680363874
transform 1 0 4524 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3074
timestamp 1680363874
transform 1 0 4516 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1680363874
transform 1 0 4524 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1680363874
transform 1 0 4508 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2778
timestamp 1680363874
transform 1 0 4516 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3076
timestamp 1680363874
transform 1 0 4572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1680363874
transform 1 0 4548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1680363874
transform 1 0 4556 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1680363874
transform 1 0 4596 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1680363874
transform 1 0 4652 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2811
timestamp 1680363874
transform 1 0 4548 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1680363874
transform 1 0 4596 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1680363874
transform 1 0 4660 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3077
timestamp 1680363874
transform 1 0 4684 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1680363874
transform 1 0 4700 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1680363874
transform 1 0 4708 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1680363874
transform 1 0 4676 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2780
timestamp 1680363874
transform 1 0 4684 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3186
timestamp 1680363874
transform 1 0 4692 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2781
timestamp 1680363874
transform 1 0 4708 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3187
timestamp 1680363874
transform 1 0 4716 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2813
timestamp 1680363874
transform 1 0 4676 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1680363874
transform 1 0 4724 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3188
timestamp 1680363874
transform 1 0 4756 0 1 3325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_28
timestamp 1680363874
transform 1 0 24 0 1 3270
box -10 -3 10 3
use FILL  FILL_2553
timestamp 1680363874
transform 1 0 72 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1680363874
transform 1 0 80 0 -1 3370
box -8 -3 104 105
use NAND2X1  NAND2X1_14
timestamp 1680363874
transform 1 0 176 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2563
timestamp 1680363874
transform 1 0 200 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1680363874
transform 1 0 208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1680363874
transform 1 0 216 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1680363874
transform 1 0 224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1680363874
transform 1 0 232 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_159
timestamp 1680363874
transform 1 0 240 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2570
timestamp 1680363874
transform 1 0 280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1680363874
transform 1 0 288 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1680363874
transform 1 0 296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1680363874
transform 1 0 304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1680363874
transform 1 0 312 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_197
timestamp 1680363874
transform 1 0 320 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2576
timestamp 1680363874
transform 1 0 336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1680363874
transform 1 0 344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1680363874
transform 1 0 352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1680363874
transform 1 0 360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1680363874
transform 1 0 368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1680363874
transform 1 0 376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1680363874
transform 1 0 384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1680363874
transform 1 0 392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1680363874
transform 1 0 400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1680363874
transform 1 0 408 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_161
timestamp 1680363874
transform -1 0 456 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2592
timestamp 1680363874
transform 1 0 456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1680363874
transform 1 0 464 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1680363874
transform 1 0 472 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_199
timestamp 1680363874
transform -1 0 496 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2595
timestamp 1680363874
transform 1 0 496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1680363874
transform 1 0 504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1680363874
transform 1 0 512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1680363874
transform 1 0 520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1680363874
transform 1 0 528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1680363874
transform 1 0 536 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_162
timestamp 1680363874
transform 1 0 544 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2607
timestamp 1680363874
transform 1 0 584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1680363874
transform 1 0 592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1680363874
transform 1 0 600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1680363874
transform 1 0 608 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_164
timestamp 1680363874
transform 1 0 616 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2615
timestamp 1680363874
transform 1 0 656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1680363874
transform 1 0 664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1680363874
transform 1 0 672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1680363874
transform 1 0 680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1680363874
transform 1 0 688 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_165
timestamp 1680363874
transform 1 0 696 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2627
timestamp 1680363874
transform 1 0 736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1680363874
transform 1 0 744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1680363874
transform 1 0 752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1680363874
transform 1 0 760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1680363874
transform 1 0 768 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_78
timestamp 1680363874
transform 1 0 776 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2638
timestamp 1680363874
transform 1 0 808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1680363874
transform 1 0 816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1680363874
transform 1 0 824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1680363874
transform 1 0 832 0 -1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_18
timestamp 1680363874
transform 1 0 840 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2646
timestamp 1680363874
transform 1 0 864 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1680363874
transform 1 0 872 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1680363874
transform 1 0 880 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1680363874
transform 1 0 888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1680363874
transform 1 0 896 0 -1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_19
timestamp 1680363874
transform -1 0 928 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2656
timestamp 1680363874
transform 1 0 928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1680363874
transform 1 0 936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1680363874
transform 1 0 944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1680363874
transform 1 0 952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1680363874
transform 1 0 960 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_80
timestamp 1680363874
transform -1 0 1000 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2669
timestamp 1680363874
transform 1 0 1000 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1680363874
transform 1 0 1008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1680363874
transform 1 0 1016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1680363874
transform 1 0 1024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1680363874
transform 1 0 1032 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_166
timestamp 1680363874
transform 1 0 1040 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2684
timestamp 1680363874
transform 1 0 1080 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1680363874
transform 1 0 1088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1680363874
transform 1 0 1096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1680363874
transform 1 0 1104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1680363874
transform 1 0 1112 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_167
timestamp 1680363874
transform 1 0 1120 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2697
timestamp 1680363874
transform 1 0 1160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1680363874
transform 1 0 1168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1680363874
transform 1 0 1176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1680363874
transform 1 0 1184 0 -1 3370
box -8 -3 16 105
use BUFX2  BUFX2_4
timestamp 1680363874
transform -1 0 1216 0 -1 3370
box -5 -3 28 105
use FILL  FILL_2726
timestamp 1680363874
transform 1 0 1216 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_203
timestamp 1680363874
transform 1 0 1224 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2727
timestamp 1680363874
transform 1 0 1240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1680363874
transform 1 0 1248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1680363874
transform 1 0 1256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1680363874
transform 1 0 1264 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_170
timestamp 1680363874
transform 1 0 1272 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2731
timestamp 1680363874
transform 1 0 1312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1680363874
transform 1 0 1320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1680363874
transform 1 0 1328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1680363874
transform 1 0 1336 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_198
timestamp 1680363874
transform -1 0 1440 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2735
timestamp 1680363874
transform 1 0 1440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1680363874
transform 1 0 1448 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_199
timestamp 1680363874
transform -1 0 1552 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2737
timestamp 1680363874
transform 1 0 1552 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1680363874
transform 1 0 1560 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1680363874
transform 1 0 1568 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_204
timestamp 1680363874
transform 1 0 1576 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2740
timestamp 1680363874
transform 1 0 1592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1680363874
transform 1 0 1600 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_171
timestamp 1680363874
transform 1 0 1608 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2742
timestamp 1680363874
transform 1 0 1648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1680363874
transform 1 0 1656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1680363874
transform 1 0 1664 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_172
timestamp 1680363874
transform 1 0 1672 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2745
timestamp 1680363874
transform 1 0 1712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1680363874
transform 1 0 1720 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_205
timestamp 1680363874
transform -1 0 1744 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2748
timestamp 1680363874
transform 1 0 1744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1680363874
transform 1 0 1752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1680363874
transform 1 0 1760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1680363874
transform 1 0 1768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1680363874
transform 1 0 1776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1680363874
transform 1 0 1784 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_82
timestamp 1680363874
transform -1 0 1824 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2760
timestamp 1680363874
transform 1 0 1824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1680363874
transform 1 0 1832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1680363874
transform 1 0 1840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1680363874
transform 1 0 1848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1680363874
transform 1 0 1856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1680363874
transform 1 0 1864 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_207
timestamp 1680363874
transform 1 0 1872 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2775
timestamp 1680363874
transform 1 0 1888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1680363874
transform 1 0 1896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1680363874
transform 1 0 1904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1680363874
transform 1 0 1912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1680363874
transform 1 0 1920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1680363874
transform 1 0 1928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1680363874
transform 1 0 1936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1680363874
transform 1 0 1944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1680363874
transform 1 0 1952 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_174
timestamp 1680363874
transform 1 0 1960 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2784
timestamp 1680363874
transform 1 0 2000 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1680363874
transform 1 0 2008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1680363874
transform 1 0 2016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1680363874
transform 1 0 2024 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_208
timestamp 1680363874
transform -1 0 2048 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2788
timestamp 1680363874
transform 1 0 2048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1680363874
transform 1 0 2056 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1680363874
transform -1 0 2160 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2800
timestamp 1680363874
transform 1 0 2160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1680363874
transform 1 0 2168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1680363874
transform 1 0 2176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1680363874
transform 1 0 2184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1680363874
transform 1 0 2192 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_175
timestamp 1680363874
transform 1 0 2200 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2805
timestamp 1680363874
transform 1 0 2240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1680363874
transform 1 0 2248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1680363874
transform 1 0 2256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1680363874
transform 1 0 2264 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_211
timestamp 1680363874
transform -1 0 2288 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2813
timestamp 1680363874
transform 1 0 2288 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1680363874
transform 1 0 2296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1680363874
transform 1 0 2304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1680363874
transform 1 0 2312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1680363874
transform 1 0 2320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1680363874
transform 1 0 2328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1680363874
transform 1 0 2336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1680363874
transform 1 0 2344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1680363874
transform 1 0 2352 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_177
timestamp 1680363874
transform 1 0 2360 0 -1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2844
timestamp 1680363874
transform 1 0 2412 0 1 3275
box -3 -3 3 3
use FILL  FILL_2834
timestamp 1680363874
transform 1 0 2400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1680363874
transform 1 0 2408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1680363874
transform 1 0 2416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1680363874
transform 1 0 2424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1680363874
transform 1 0 2432 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_204
timestamp 1680363874
transform 1 0 2440 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2839
timestamp 1680363874
transform 1 0 2536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1680363874
transform 1 0 2544 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1680363874
transform 1 0 2552 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1680363874
transform 1 0 2560 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_179
timestamp 1680363874
transform 1 0 2568 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2850
timestamp 1680363874
transform 1 0 2608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1680363874
transform 1 0 2616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1680363874
transform 1 0 2624 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1680363874
transform 1 0 2632 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1680363874
transform 1 0 2640 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1680363874
transform 1 0 2648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1680363874
transform 1 0 2656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1680363874
transform 1 0 2664 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1680363874
transform 1 0 2672 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2868
timestamp 1680363874
transform 1 0 2768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1680363874
transform 1 0 2776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1680363874
transform 1 0 2784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1680363874
transform 1 0 2792 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_182
timestamp 1680363874
transform 1 0 2800 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2877
timestamp 1680363874
transform 1 0 2840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1680363874
transform 1 0 2848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1680363874
transform 1 0 2856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1680363874
transform 1 0 2864 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_183
timestamp 1680363874
transform 1 0 2872 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2886
timestamp 1680363874
transform 1 0 2912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1680363874
transform 1 0 2920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1680363874
transform 1 0 2928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1680363874
transform 1 0 2936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1680363874
transform 1 0 2944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1680363874
transform 1 0 2952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1680363874
transform 1 0 2960 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1680363874
transform -1 0 3064 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2905
timestamp 1680363874
transform 1 0 3064 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1680363874
transform 1 0 3072 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1680363874
transform 1 0 3080 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1680363874
transform 1 0 3088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1680363874
transform 1 0 3096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1680363874
transform 1 0 3104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1680363874
transform 1 0 3112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1680363874
transform 1 0 3120 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_85
timestamp 1680363874
transform 1 0 3128 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2922
timestamp 1680363874
transform 1 0 3160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1680363874
transform 1 0 3168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1680363874
transform 1 0 3176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1680363874
transform 1 0 3184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1680363874
transform 1 0 3192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1680363874
transform 1 0 3200 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1680363874
transform -1 0 3240 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2928
timestamp 1680363874
transform 1 0 3240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1680363874
transform 1 0 3248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1680363874
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_218
timestamp 1680363874
transform 1 0 3264 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2931
timestamp 1680363874
transform 1 0 3280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1680363874
transform 1 0 3288 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1680363874
transform 1 0 3296 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_119
timestamp 1680363874
transform -1 0 3344 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2937
timestamp 1680363874
transform 1 0 3344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1680363874
transform 1 0 3352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1680363874
transform 1 0 3360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1680363874
transform 1 0 3368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1680363874
transform 1 0 3376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1680363874
transform 1 0 3384 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1680363874
transform -1 0 3488 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2955
timestamp 1680363874
transform 1 0 3488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1680363874
transform 1 0 3496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1680363874
transform 1 0 3504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1680363874
transform 1 0 3512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1680363874
transform 1 0 3520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1680363874
transform 1 0 3528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1680363874
transform 1 0 3536 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2845
timestamp 1680363874
transform 1 0 3564 0 1 3275
box -3 -3 3 3
use AND2X2  AND2X2_4
timestamp 1680363874
transform 1 0 3544 0 -1 3370
box -8 -3 40 105
use FILL  FILL_2962
timestamp 1680363874
transform 1 0 3576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1680363874
transform 1 0 3584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1680363874
transform 1 0 3592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1680363874
transform 1 0 3600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1680363874
transform 1 0 3608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1680363874
transform 1 0 3616 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_120
timestamp 1680363874
transform -1 0 3664 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2974
timestamp 1680363874
transform 1 0 3664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1680363874
transform 1 0 3672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1680363874
transform 1 0 3680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1680363874
transform 1 0 3688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1680363874
transform 1 0 3696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1680363874
transform 1 0 3704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1680363874
transform 1 0 3712 0 -1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_27
timestamp 1680363874
transform -1 0 3744 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2981
timestamp 1680363874
transform 1 0 3744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1680363874
transform 1 0 3752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1680363874
transform 1 0 3760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1680363874
transform 1 0 3768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1680363874
transform 1 0 3776 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_121
timestamp 1680363874
transform -1 0 3824 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2986
timestamp 1680363874
transform 1 0 3824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1680363874
transform 1 0 3832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1680363874
transform 1 0 3840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1680363874
transform 1 0 3848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1680363874
transform 1 0 3856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1680363874
transform 1 0 3864 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1680363874
transform 1 0 3872 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1680363874
transform 1 0 3880 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1680363874
transform 1 0 3888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1680363874
transform 1 0 3896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1680363874
transform 1 0 3904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1680363874
transform 1 0 3912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1680363874
transform 1 0 3920 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1680363874
transform -1 0 4024 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3016
timestamp 1680363874
transform 1 0 4024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1680363874
transform 1 0 4032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1680363874
transform 1 0 4040 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1680363874
transform 1 0 4048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1680363874
transform 1 0 4056 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1680363874
transform 1 0 4064 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_123
timestamp 1680363874
transform 1 0 4072 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3032
timestamp 1680363874
transform 1 0 4112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1680363874
transform 1 0 4120 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_223
timestamp 1680363874
transform 1 0 4128 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3034
timestamp 1680363874
transform 1 0 4144 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1680363874
transform 1 0 4152 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1680363874
transform 1 0 4160 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3036
timestamp 1680363874
transform 1 0 4256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1680363874
transform 1 0 4264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1680363874
transform 1 0 4272 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1680363874
transform 1 0 4280 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_124
timestamp 1680363874
transform -1 0 4328 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3046
timestamp 1680363874
transform 1 0 4328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1680363874
transform 1 0 4336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1680363874
transform 1 0 4344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1680363874
transform 1 0 4352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1680363874
transform 1 0 4360 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_225
timestamp 1680363874
transform 1 0 4368 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3070
timestamp 1680363874
transform 1 0 4384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1680363874
transform 1 0 4392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1680363874
transform 1 0 4400 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_125
timestamp 1680363874
transform 1 0 4408 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3073
timestamp 1680363874
transform 1 0 4448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1680363874
transform 1 0 4456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1680363874
transform 1 0 4464 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1680363874
transform 1 0 4472 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1680363874
transform 1 0 4480 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_126
timestamp 1680363874
transform -1 0 4528 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3078
timestamp 1680363874
transform 1 0 4528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1680363874
transform 1 0 4536 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_226
timestamp 1680363874
transform 1 0 4544 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1680363874
transform 1 0 4560 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3080
timestamp 1680363874
transform 1 0 4656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1680363874
transform 1 0 4664 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_127
timestamp 1680363874
transform 1 0 4672 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3085
timestamp 1680363874
transform 1 0 4712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1680363874
transform 1 0 4720 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1680363874
transform 1 0 4728 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_228
timestamp 1680363874
transform 1 0 4736 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3088
timestamp 1680363874
transform 1 0 4752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1680363874
transform 1 0 4760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1680363874
transform 1 0 4768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1680363874
transform 1 0 4776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1680363874
transform 1 0 4784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1680363874
transform 1 0 4792 0 -1 3370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_29
timestamp 1680363874
transform 1 0 4851 0 1 3270
box -10 -3 10 3
use M3_M2  M3_M2_2846
timestamp 1680363874
transform 1 0 92 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1680363874
transform 1 0 156 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1680363874
transform 1 0 180 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3219
timestamp 1680363874
transform 1 0 116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1680363874
transform 1 0 172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1680363874
transform 1 0 180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1680363874
transform 1 0 84 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1680363874
transform 1 0 172 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2945
timestamp 1680363874
transform 1 0 180 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3311
timestamp 1680363874
transform 1 0 188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1680363874
transform 1 0 220 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2946
timestamp 1680363874
transform 1 0 212 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3222
timestamp 1680363874
transform 1 0 268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1680363874
transform 1 0 284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1680363874
transform 1 0 276 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2961
timestamp 1680363874
transform 1 0 276 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3313
timestamp 1680363874
transform 1 0 292 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2962
timestamp 1680363874
transform 1 0 292 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3199
timestamp 1680363874
transform 1 0 316 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2928
timestamp 1680363874
transform 1 0 316 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3200
timestamp 1680363874
transform 1 0 332 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2963
timestamp 1680363874
transform 1 0 324 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1680363874
transform 1 0 340 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3314
timestamp 1680363874
transform 1 0 340 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1680363874
transform 1 0 356 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2947
timestamp 1680363874
transform 1 0 364 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1680363874
transform 1 0 388 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3316
timestamp 1680363874
transform 1 0 380 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1680363874
transform 1 0 388 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2847
timestamp 1680363874
transform 1 0 436 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1680363874
transform 1 0 428 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3224
timestamp 1680363874
transform 1 0 404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1680363874
transform 1 0 420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1680363874
transform 1 0 396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1680363874
transform 1 0 428 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1680363874
transform 1 0 444 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1680363874
transform 1 0 452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1680363874
transform 1 0 476 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2930
timestamp 1680363874
transform 1 0 476 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1680363874
transform 1 0 492 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3320
timestamp 1680363874
transform 1 0 484 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2964
timestamp 1680363874
transform 1 0 476 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1680363874
transform 1 0 524 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3204
timestamp 1680363874
transform 1 0 572 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1680363874
transform 1 0 564 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2848
timestamp 1680363874
transform 1 0 620 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1680363874
transform 1 0 612 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1680363874
transform 1 0 636 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3226
timestamp 1680363874
transform 1 0 604 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2893
timestamp 1680363874
transform 1 0 620 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3227
timestamp 1680363874
transform 1 0 620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1680363874
transform 1 0 636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1680363874
transform 1 0 652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1680363874
transform 1 0 628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1680363874
transform 1 0 644 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2966
timestamp 1680363874
transform 1 0 628 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1680363874
transform 1 0 660 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3230
timestamp 1680363874
transform 1 0 708 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2948
timestamp 1680363874
transform 1 0 708 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1680363874
transform 1 0 724 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1680363874
transform 1 0 724 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3324
timestamp 1680363874
transform 1 0 740 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1680363874
transform 1 0 748 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2996
timestamp 1680363874
transform 1 0 740 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3205
timestamp 1680363874
transform 1 0 764 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1680363874
transform 1 0 764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1680363874
transform 1 0 804 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1680363874
transform 1 0 828 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2967
timestamp 1680363874
transform 1 0 828 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1680363874
transform 1 0 868 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1680363874
transform 1 0 860 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1680363874
transform 1 0 852 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3231
timestamp 1680363874
transform 1 0 844 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2949
timestamp 1680363874
transform 1 0 844 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3232
timestamp 1680363874
transform 1 0 868 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2897
timestamp 1680363874
transform 1 0 884 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3207
timestamp 1680363874
transform 1 0 892 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1680363874
transform 1 0 892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1680363874
transform 1 0 908 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2968
timestamp 1680363874
transform 1 0 908 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3208
timestamp 1680363874
transform 1 0 940 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1680363874
transform 1 0 956 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2932
timestamp 1680363874
transform 1 0 948 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1680363874
transform 1 0 948 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3329
timestamp 1680363874
transform 1 0 996 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2997
timestamp 1680363874
transform 1 0 980 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1680363874
transform 1 0 1012 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1680363874
transform 1 0 1068 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3234
timestamp 1680363874
transform 1 0 1044 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1680363874
transform 1 0 1052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1680363874
transform 1 0 1068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1680363874
transform 1 0 1044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1680363874
transform 1 0 1060 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2950
timestamp 1680363874
transform 1 0 1068 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1680363874
transform 1 0 1044 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3237
timestamp 1680363874
transform 1 0 1084 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1680363874
transform 1 0 1092 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2971
timestamp 1680363874
transform 1 0 1084 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1680363874
transform 1 0 1092 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1680363874
transform 1 0 1156 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1680363874
transform 1 0 1132 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1680363874
transform 1 0 1148 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3333
timestamp 1680363874
transform 1 0 1124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1680363874
transform 1 0 1156 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1680363874
transform 1 0 1148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1680363874
transform 1 0 1172 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2972
timestamp 1680363874
transform 1 0 1172 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3335
timestamp 1680363874
transform 1 0 1196 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2973
timestamp 1680363874
transform 1 0 1196 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1680363874
transform 1 0 1220 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3240
timestamp 1680363874
transform 1 0 1220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1680363874
transform 1 0 1220 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2878
timestamp 1680363874
transform 1 0 1260 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3241
timestamp 1680363874
transform 1 0 1260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1680363874
transform 1 0 1236 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1680363874
transform 1 0 1252 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1680363874
transform 1 0 1268 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2974
timestamp 1680363874
transform 1 0 1228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1680363874
transform 1 0 1268 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1680363874
transform 1 0 1284 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3242
timestamp 1680363874
transform 1 0 1284 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2879
timestamp 1680363874
transform 1 0 1300 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3340
timestamp 1680363874
transform 1 0 1332 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1680363874
transform 1 0 1340 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2855
timestamp 1680363874
transform 1 0 1372 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1680363874
transform 1 0 1388 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3243
timestamp 1680363874
transform 1 0 1372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1680363874
transform 1 0 1388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1680363874
transform 1 0 1380 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1680363874
transform 1 0 1396 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2976
timestamp 1680363874
transform 1 0 1380 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1680363874
transform 1 0 1388 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3245
timestamp 1680363874
transform 1 0 1468 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1680363874
transform 1 0 1444 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2977
timestamp 1680363874
transform 1 0 1468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1680363874
transform 1 0 1540 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3246
timestamp 1680363874
transform 1 0 1532 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1680363874
transform 1 0 1540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1680363874
transform 1 0 1548 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3000
timestamp 1680363874
transform 1 0 1548 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3346
timestamp 1680363874
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2905
timestamp 1680363874
transform 1 0 1612 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1680363874
transform 1 0 1636 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3248
timestamp 1680363874
transform 1 0 1612 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1680363874
transform 1 0 1620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1680363874
transform 1 0 1636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1680363874
transform 1 0 1612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1680363874
transform 1 0 1628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1680363874
transform 1 0 1644 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2978
timestamp 1680363874
transform 1 0 1612 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1680363874
transform 1 0 1660 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1680363874
transform 1 0 1692 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3251
timestamp 1680363874
transform 1 0 1692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1680363874
transform 1 0 1708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1680363874
transform 1 0 1684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1680363874
transform 1 0 1700 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2951
timestamp 1680363874
transform 1 0 1708 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1680363874
transform 1 0 1724 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3352
timestamp 1680363874
transform 1 0 1716 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2980
timestamp 1680363874
transform 1 0 1684 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1680363874
transform 1 0 1780 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3253
timestamp 1680363874
transform 1 0 1748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1680363874
transform 1 0 1780 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2934
timestamp 1680363874
transform 1 0 1788 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1680363874
transform 1 0 1828 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1680363874
transform 1 0 1756 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3353
timestamp 1680363874
transform 1 0 1828 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2981
timestamp 1680363874
transform 1 0 1828 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1680363874
transform 1 0 1796 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3255
timestamp 1680363874
transform 1 0 1852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1680363874
transform 1 0 1900 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1680363874
transform 1 0 1932 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2982
timestamp 1680363874
transform 1 0 1932 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1680363874
transform 1 0 1948 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1680363874
transform 1 0 2020 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1680363874
transform 1 0 1964 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3257
timestamp 1680363874
transform 1 0 1988 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2936
timestamp 1680363874
transform 1 0 2028 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1680363874
transform 1 0 2060 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1680363874
transform 1 0 2052 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3258
timestamp 1680363874
transform 1 0 2044 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1680363874
transform 1 0 2052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1680363874
transform 1 0 1964 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2983
timestamp 1680363874
transform 1 0 1964 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1680363874
transform 1 0 2084 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3260
timestamp 1680363874
transform 1 0 2076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1680363874
transform 1 0 2108 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2937
timestamp 1680363874
transform 1 0 2116 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3356
timestamp 1680363874
transform 1 0 2084 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1680363874
transform 1 0 2100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1680363874
transform 1 0 2116 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1680363874
transform 1 0 2148 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1680363874
transform 1 0 2172 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2984
timestamp 1680363874
transform 1 0 2172 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1680363874
transform 1 0 2196 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1680363874
transform 1 0 2268 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1680363874
transform 1 0 2284 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3263
timestamp 1680363874
transform 1 0 2236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1680363874
transform 1 0 2292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1680363874
transform 1 0 2212 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2986
timestamp 1680363874
transform 1 0 2228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1680363874
transform 1 0 2204 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1680363874
transform 1 0 2260 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1680363874
transform 1 0 2292 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3361
timestamp 1680363874
transform 1 0 2308 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2859
timestamp 1680363874
transform 1 0 2340 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3210
timestamp 1680363874
transform 1 0 2356 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1680363874
transform 1 0 2340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1680363874
transform 1 0 2356 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2851
timestamp 1680363874
transform 1 0 2380 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3211
timestamp 1680363874
transform 1 0 2388 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2911
timestamp 1680363874
transform 1 0 2396 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1680363874
transform 1 0 2388 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3362
timestamp 1680363874
transform 1 0 2388 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2912
timestamp 1680363874
transform 1 0 2412 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3267
timestamp 1680363874
transform 1 0 2404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1680363874
transform 1 0 2412 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2882
timestamp 1680363874
transform 1 0 2428 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1680363874
transform 1 0 2428 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1680363874
transform 1 0 2420 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1680363874
transform 1 0 2452 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3212
timestamp 1680363874
transform 1 0 2460 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1680363874
transform 1 0 2452 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2987
timestamp 1680363874
transform 1 0 2460 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1680363874
transform 1 0 2460 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1680363874
transform 1 0 2484 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3399
timestamp 1680363874
transform 1 0 2476 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1680363874
transform 1 0 2500 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2939
timestamp 1680363874
transform 1 0 2500 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1680363874
transform 1 0 2500 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1680363874
transform 1 0 2540 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3365
timestamp 1680363874
transform 1 0 2556 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2915
timestamp 1680363874
transform 1 0 2572 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1680363874
transform 1 0 2588 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3268
timestamp 1680363874
transform 1 0 2588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1680363874
transform 1 0 2596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1680363874
transform 1 0 2612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1680363874
transform 1 0 2628 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2916
timestamp 1680363874
transform 1 0 2644 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1680363874
transform 1 0 2684 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3271
timestamp 1680363874
transform 1 0 2692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1680363874
transform 1 0 2740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1680363874
transform 1 0 2644 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2955
timestamp 1680363874
transform 1 0 2692 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1680363874
transform 1 0 2724 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1680363874
transform 1 0 2756 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1680363874
transform 1 0 2852 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3273
timestamp 1680363874
transform 1 0 2820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1680363874
transform 1 0 2788 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2988
timestamp 1680363874
transform 1 0 2860 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1680363874
transform 1 0 2876 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3274
timestamp 1680363874
transform 1 0 2916 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2989
timestamp 1680363874
transform 1 0 2932 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1680363874
transform 1 0 2972 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3214
timestamp 1680363874
transform 1 0 2972 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1680363874
transform 1 0 2956 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2990
timestamp 1680363874
transform 1 0 2956 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1680363874
transform 1 0 2988 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1680363874
transform 1 0 3028 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1680363874
transform 1 0 3012 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3276
timestamp 1680363874
transform 1 0 3028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1680363874
transform 1 0 3012 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2940
timestamp 1680363874
transform 1 0 3036 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3370
timestamp 1680363874
transform 1 0 3052 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1680363874
transform 1 0 3060 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1680363874
transform 1 0 3044 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2884
timestamp 1680363874
transform 1 0 3076 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1680363874
transform 1 0 3076 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3277
timestamp 1680363874
transform 1 0 3076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1680363874
transform 1 0 3076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1680363874
transform 1 0 3092 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2873
timestamp 1680363874
transform 1 0 3116 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1680363874
transform 1 0 3132 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1680363874
transform 1 0 3132 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3215
timestamp 1680363874
transform 1 0 3132 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1680363874
transform 1 0 3140 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2863
timestamp 1680363874
transform 1 0 3164 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1680363874
transform 1 0 3156 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1680363874
transform 1 0 3188 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1680363874
transform 1 0 3180 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3279
timestamp 1680363874
transform 1 0 3180 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2957
timestamp 1680363874
transform 1 0 3180 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3373
timestamp 1680363874
transform 1 0 3188 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2887
timestamp 1680363874
transform 1 0 3212 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1680363874
transform 1 0 3212 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3280
timestamp 1680363874
transform 1 0 3212 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2992
timestamp 1680363874
transform 1 0 3204 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3281
timestamp 1680363874
transform 1 0 3244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1680363874
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1680363874
transform 1 0 3268 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3008
timestamp 1680363874
transform 1 0 3268 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1680363874
transform 1 0 3284 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1680363874
transform 1 0 3324 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3282
timestamp 1680363874
transform 1 0 3284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1680363874
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1680363874
transform 1 0 3324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1680363874
transform 1 0 3372 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3009
timestamp 1680363874
transform 1 0 3284 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1680363874
transform 1 0 3380 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1680363874
transform 1 0 3420 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3285
timestamp 1680363874
transform 1 0 3428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1680363874
transform 1 0 3420 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1680363874
transform 1 0 3452 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1680363874
transform 1 0 3460 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_3011
timestamp 1680363874
transform 1 0 3460 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3288
timestamp 1680363874
transform 1 0 3492 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1680363874
transform 1 0 3484 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3012
timestamp 1680363874
transform 1 0 3492 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1680363874
transform 1 0 3508 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1680363874
transform 1 0 3548 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3289
timestamp 1680363874
transform 1 0 3548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1680363874
transform 1 0 3540 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2876
timestamp 1680363874
transform 1 0 3588 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3217
timestamp 1680363874
transform 1 0 3588 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1680363874
transform 1 0 3588 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1680363874
transform 1 0 3580 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1680363874
transform 1 0 3620 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1680363874
transform 1 0 3652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1680363874
transform 1 0 3668 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1680363874
transform 1 0 3684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1680363874
transform 1 0 3716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1680363874
transform 1 0 3708 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2864
timestamp 1680363874
transform 1 0 3748 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3292
timestamp 1680363874
transform 1 0 3748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1680363874
transform 1 0 3740 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3013
timestamp 1680363874
transform 1 0 3740 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3293
timestamp 1680363874
transform 1 0 3796 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1680363874
transform 1 0 3836 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1680363874
transform 1 0 3876 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3014
timestamp 1680363874
transform 1 0 3844 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3387
timestamp 1680363874
transform 1 0 3932 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1680363874
transform 1 0 3948 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1680363874
transform 1 0 3964 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1680363874
transform 1 0 3956 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1680363874
transform 1 0 3980 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2958
timestamp 1680363874
transform 1 0 3980 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1680363874
transform 1 0 4028 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3389
timestamp 1680363874
transform 1 0 4028 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1680363874
transform 1 0 4036 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2925
timestamp 1680363874
transform 1 0 4052 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3298
timestamp 1680363874
transform 1 0 4052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1680363874
transform 1 0 4060 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1680363874
transform 1 0 4092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1680363874
transform 1 0 4148 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1680363874
transform 1 0 4172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1680363874
transform 1 0 4188 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2993
timestamp 1680363874
transform 1 0 4188 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3392
timestamp 1680363874
transform 1 0 4228 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1680363874
transform 1 0 4244 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1680363874
transform 1 0 4436 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1680363874
transform 1 0 4452 0 1 3235
box -2 -2 2 2
use M3_M2  M3_M2_2943
timestamp 1680363874
transform 1 0 4468 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1680363874
transform 1 0 4508 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1680363874
transform 1 0 4484 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3302
timestamp 1680363874
transform 1 0 4492 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2944
timestamp 1680363874
transform 1 0 4500 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3303
timestamp 1680363874
transform 1 0 4508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1680363874
transform 1 0 4484 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1680363874
transform 1 0 4500 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3015
timestamp 1680363874
transform 1 0 4492 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1680363874
transform 1 0 4532 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1680363874
transform 1 0 4532 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1680363874
transform 1 0 4556 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1680363874
transform 1 0 4588 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3395
timestamp 1680363874
transform 1 0 4548 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2994
timestamp 1680363874
transform 1 0 4548 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1680363874
transform 1 0 4644 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3304
timestamp 1680363874
transform 1 0 4588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1680363874
transform 1 0 4644 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1680363874
transform 1 0 4660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1680363874
transform 1 0 4564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1680363874
transform 1 0 4652 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1680363874
transform 1 0 4676 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1680363874
transform 1 0 4676 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3218
timestamp 1680363874
transform 1 0 4700 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1680363874
transform 1 0 4756 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2960
timestamp 1680363874
transform 1 0 4748 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3398
timestamp 1680363874
transform 1 0 4788 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_3016
timestamp 1680363874
transform 1 0 4804 0 1 3185
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_30
timestamp 1680363874
transform 1 0 48 0 1 3170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_218
timestamp 1680363874
transform 1 0 72 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_229
timestamp 1680363874
transform 1 0 168 0 1 3170
box -9 -3 26 105
use NAND2X1  NAND2X1_20
timestamp 1680363874
transform 1 0 184 0 1 3170
box -8 -3 32 105
use FILL  FILL_3094
timestamp 1680363874
transform 1 0 208 0 1 3170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1680363874
transform 1 0 216 0 1 3170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1680363874
transform 1 0 224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1680363874
transform 1 0 232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1680363874
transform 1 0 240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1680363874
transform 1 0 248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1680363874
transform 1 0 256 0 1 3170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1680363874
transform 1 0 264 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_22
timestamp 1680363874
transform 1 0 272 0 1 3170
box -8 -3 32 105
use FILL  FILL_3105
timestamp 1680363874
transform 1 0 296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1680363874
transform 1 0 304 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_23
timestamp 1680363874
transform 1 0 312 0 1 3170
box -8 -3 32 105
use FILL  FILL_3107
timestamp 1680363874
transform 1 0 336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1680363874
transform 1 0 344 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3017
timestamp 1680363874
transform 1 0 372 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1680363874
transform 1 0 388 0 1 3175
box -3 -3 3 3
use OAI21X1  OAI21X1_89
timestamp 1680363874
transform 1 0 352 0 1 3170
box -8 -3 34 105
use FILL  FILL_3114
timestamp 1680363874
transform 1 0 384 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3019
timestamp 1680363874
transform 1 0 428 0 1 3175
box -3 -3 3 3
use OAI21X1  OAI21X1_91
timestamp 1680363874
transform 1 0 392 0 1 3170
box -8 -3 34 105
use FILL  FILL_3115
timestamp 1680363874
transform 1 0 424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1680363874
transform 1 0 432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1680363874
transform 1 0 440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1680363874
transform 1 0 448 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_26
timestamp 1680363874
transform 1 0 456 0 1 3170
box -8 -3 32 105
use FILL  FILL_3119
timestamp 1680363874
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1680363874
transform 1 0 488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1680363874
transform 1 0 496 0 1 3170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1680363874
transform 1 0 504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1680363874
transform 1 0 512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1680363874
transform 1 0 520 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_92
timestamp 1680363874
transform 1 0 528 0 1 3170
box -8 -3 34 105
use M3_M2  M3_M2_3020
timestamp 1680363874
transform 1 0 572 0 1 3175
box -3 -3 3 3
use FILL  FILL_3134
timestamp 1680363874
transform 1 0 560 0 1 3170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1680363874
transform 1 0 568 0 1 3170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1680363874
transform 1 0 576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1680363874
transform 1 0 584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1680363874
transform 1 0 592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1680363874
transform 1 0 600 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3021
timestamp 1680363874
transform 1 0 636 0 1 3175
box -3 -3 3 3
use OAI22X1  OAI22X1_187
timestamp 1680363874
transform 1 0 608 0 1 3170
box -8 -3 46 105
use FILL  FILL_3146
timestamp 1680363874
transform 1 0 648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1680363874
transform 1 0 656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1680363874
transform 1 0 664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1680363874
transform 1 0 672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1680363874
transform 1 0 680 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_234
timestamp 1680363874
transform -1 0 704 0 1 3170
box -9 -3 26 105
use FILL  FILL_3157
timestamp 1680363874
transform 1 0 704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1680363874
transform 1 0 712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1680363874
transform 1 0 720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1680363874
transform 1 0 728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1680363874
transform 1 0 736 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3022
timestamp 1680363874
transform 1 0 764 0 1 3175
box -3 -3 3 3
use NAND2X1  NAND2X1_28
timestamp 1680363874
transform 1 0 744 0 1 3170
box -8 -3 32 105
use FILL  FILL_3165
timestamp 1680363874
transform 1 0 768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1680363874
transform 1 0 776 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3023
timestamp 1680363874
transform 1 0 796 0 1 3175
box -3 -3 3 3
use FILL  FILL_3167
timestamp 1680363874
transform 1 0 784 0 1 3170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1680363874
transform 1 0 792 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_95
timestamp 1680363874
transform -1 0 832 0 1 3170
box -8 -3 34 105
use FILL  FILL_3169
timestamp 1680363874
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1680363874
transform 1 0 840 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_235
timestamp 1680363874
transform -1 0 864 0 1 3170
box -9 -3 26 105
use FILL  FILL_3171
timestamp 1680363874
transform 1 0 864 0 1 3170
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1680363874
transform 1 0 872 0 1 3170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1680363874
transform 1 0 880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1680363874
transform 1 0 888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1680363874
transform 1 0 896 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_29
timestamp 1680363874
transform -1 0 928 0 1 3170
box -8 -3 32 105
use FILL  FILL_3180
timestamp 1680363874
transform 1 0 928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1680363874
transform 1 0 936 0 1 3170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1680363874
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1680363874
transform 1 0 952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1680363874
transform 1 0 960 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_96
timestamp 1680363874
transform -1 0 1000 0 1 3170
box -8 -3 34 105
use FILL  FILL_3185
timestamp 1680363874
transform 1 0 1000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1680363874
transform 1 0 1008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1680363874
transform 1 0 1016 0 1 3170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1680363874
transform 1 0 1024 0 1 3170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1680363874
transform 1 0 1032 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_188
timestamp 1680363874
transform 1 0 1040 0 1 3170
box -8 -3 46 105
use FILL  FILL_3198
timestamp 1680363874
transform 1 0 1080 0 1 3170
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1680363874
transform 1 0 1088 0 1 3170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1680363874
transform 1 0 1096 0 1 3170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1680363874
transform 1 0 1104 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3024
timestamp 1680363874
transform 1 0 1124 0 1 3175
box -3 -3 3 3
use FILL  FILL_3206
timestamp 1680363874
transform 1 0 1112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1680363874
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_190
timestamp 1680363874
transform 1 0 1128 0 1 3170
box -8 -3 46 105
use FILL  FILL_3210
timestamp 1680363874
transform 1 0 1168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1680363874
transform 1 0 1176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1680363874
transform 1 0 1184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1680363874
transform 1 0 1192 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_239
timestamp 1680363874
transform -1 0 1216 0 1 3170
box -9 -3 26 105
use FILL  FILL_3214
timestamp 1680363874
transform 1 0 1216 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3025
timestamp 1680363874
transform 1 0 1236 0 1 3175
box -3 -3 3 3
use FILL  FILL_3215
timestamp 1680363874
transform 1 0 1224 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_191
timestamp 1680363874
transform 1 0 1232 0 1 3170
box -8 -3 46 105
use FILL  FILL_3216
timestamp 1680363874
transform 1 0 1272 0 1 3170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1680363874
transform 1 0 1280 0 1 3170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1680363874
transform 1 0 1288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1680363874
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1680363874
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1680363874
transform 1 0 1312 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_240
timestamp 1680363874
transform -1 0 1336 0 1 3170
box -9 -3 26 105
use FILL  FILL_3222
timestamp 1680363874
transform 1 0 1336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1680363874
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1680363874
transform 1 0 1352 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_192
timestamp 1680363874
transform -1 0 1400 0 1 3170
box -8 -3 46 105
use FILL  FILL_3225
timestamp 1680363874
transform 1 0 1400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1680363874
transform 1 0 1408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1680363874
transform 1 0 1416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1680363874
transform 1 0 1424 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3026
timestamp 1680363874
transform 1 0 1508 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_223
timestamp 1680363874
transform 1 0 1432 0 1 3170
box -8 -3 104 105
use FILL  FILL_3233
timestamp 1680363874
transform 1 0 1528 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_242
timestamp 1680363874
transform -1 0 1552 0 1 3170
box -9 -3 26 105
use FILL  FILL_3234
timestamp 1680363874
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1680363874
transform 1 0 1560 0 1 3170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1680363874
transform 1 0 1568 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_243
timestamp 1680363874
transform 1 0 1576 0 1 3170
box -9 -3 26 105
use FILL  FILL_3237
timestamp 1680363874
transform 1 0 1592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1680363874
transform 1 0 1600 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_193
timestamp 1680363874
transform 1 0 1608 0 1 3170
box -8 -3 46 105
use FILL  FILL_3239
timestamp 1680363874
transform 1 0 1648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1680363874
transform 1 0 1656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1680363874
transform 1 0 1664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1680363874
transform 1 0 1672 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_194
timestamp 1680363874
transform -1 0 1720 0 1 3170
box -8 -3 46 105
use FILL  FILL_3243
timestamp 1680363874
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1680363874
transform 1 0 1728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1680363874
transform 1 0 1736 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1680363874
transform -1 0 1840 0 1 3170
box -8 -3 104 105
use FILL  FILL_3254
timestamp 1680363874
transform 1 0 1840 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1680363874
transform -1 0 1944 0 1 3170
box -8 -3 104 105
use FILL  FILL_3255
timestamp 1680363874
transform 1 0 1944 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1680363874
transform 1 0 1952 0 1 3170
box -8 -3 104 105
use FILL  FILL_3256
timestamp 1680363874
transform 1 0 2048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1680363874
transform 1 0 2056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1680363874
transform 1 0 2064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1680363874
transform 1 0 2072 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_198
timestamp 1680363874
transform 1 0 2080 0 1 3170
box -8 -3 46 105
use FILL  FILL_3284
timestamp 1680363874
transform 1 0 2120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1680363874
transform 1 0 2128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1680363874
transform 1 0 2136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1680363874
transform 1 0 2144 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_8
timestamp 1680363874
transform 1 0 2152 0 1 3170
box -5 -3 28 105
use FILL  FILL_3292
timestamp 1680363874
transform 1 0 2176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1680363874
transform 1 0 2184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1680363874
transform 1 0 2192 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1680363874
transform 1 0 2200 0 1 3170
box -8 -3 104 105
use FILL  FILL_3299
timestamp 1680363874
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1680363874
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1680363874
transform 1 0 2312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1680363874
transform 1 0 2320 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_97
timestamp 1680363874
transform 1 0 2328 0 1 3170
box -8 -3 34 105
use FILL  FILL_3312
timestamp 1680363874
transform 1 0 2360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1680363874
transform 1 0 2368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1680363874
transform 1 0 2376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1680363874
transform 1 0 2384 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_247
timestamp 1680363874
transform -1 0 2408 0 1 3170
box -9 -3 26 105
use FILL  FILL_3322
timestamp 1680363874
transform 1 0 2408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1680363874
transform 1 0 2416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1680363874
transform 1 0 2424 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3027
timestamp 1680363874
transform 1 0 2452 0 1 3175
box -3 -3 3 3
use NAND2X1  NAND2X1_30
timestamp 1680363874
transform 1 0 2432 0 1 3170
box -8 -3 32 105
use FILL  FILL_3329
timestamp 1680363874
transform 1 0 2456 0 1 3170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1680363874
transform 1 0 2464 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3028
timestamp 1680363874
transform 1 0 2492 0 1 3175
box -3 -3 3 3
use NOR2X1  NOR2X1_28
timestamp 1680363874
transform 1 0 2472 0 1 3170
box -8 -3 32 105
use FILL  FILL_3331
timestamp 1680363874
transform 1 0 2496 0 1 3170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1680363874
transform 1 0 2504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1680363874
transform 1 0 2512 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3029
timestamp 1680363874
transform 1 0 2548 0 1 3175
box -3 -3 3 3
use OAI21X1  OAI21X1_98
timestamp 1680363874
transform -1 0 2552 0 1 3170
box -8 -3 34 105
use FILL  FILL_3334
timestamp 1680363874
transform 1 0 2552 0 1 3170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1680363874
transform 1 0 2560 0 1 3170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1680363874
transform 1 0 2568 0 1 3170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1680363874
transform 1 0 2576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1680363874
transform 1 0 2584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1680363874
transform 1 0 2592 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3030
timestamp 1680363874
transform 1 0 2612 0 1 3175
box -3 -3 3 3
use INVX2  INVX2_249
timestamp 1680363874
transform -1 0 2616 0 1 3170
box -9 -3 26 105
use FILL  FILL_3348
timestamp 1680363874
transform 1 0 2616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1680363874
transform 1 0 2624 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1680363874
transform 1 0 2632 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_250
timestamp 1680363874
transform 1 0 2728 0 1 3170
box -9 -3 26 105
use FILL  FILL_3350
timestamp 1680363874
transform 1 0 2744 0 1 3170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1680363874
transform 1 0 2752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1680363874
transform 1 0 2760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1680363874
transform 1 0 2768 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1680363874
transform 1 0 2776 0 1 3170
box -8 -3 104 105
use FILL  FILL_3367
timestamp 1680363874
transform 1 0 2872 0 1 3170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1680363874
transform 1 0 2880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1680363874
transform 1 0 2888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1680363874
transform 1 0 2896 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_251
timestamp 1680363874
transform 1 0 2904 0 1 3170
box -9 -3 26 105
use FILL  FILL_3379
timestamp 1680363874
transform 1 0 2920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1680363874
transform 1 0 2928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1680363874
transform 1 0 2936 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_99
timestamp 1680363874
transform 1 0 2944 0 1 3170
box -8 -3 34 105
use FILL  FILL_3385
timestamp 1680363874
transform 1 0 2976 0 1 3170
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1680363874
transform 1 0 2984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1680363874
transform 1 0 2992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1680363874
transform 1 0 3000 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_100
timestamp 1680363874
transform -1 0 3040 0 1 3170
box -8 -3 34 105
use FILL  FILL_3392
timestamp 1680363874
transform 1 0 3040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1680363874
transform 1 0 3048 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_29
timestamp 1680363874
transform 1 0 3056 0 1 3170
box -8 -3 32 105
use FILL  FILL_3399
timestamp 1680363874
transform 1 0 3080 0 1 3170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1680363874
transform 1 0 3088 0 1 3170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1680363874
transform 1 0 3096 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_101
timestamp 1680363874
transform 1 0 3104 0 1 3170
box -8 -3 34 105
use FILL  FILL_3408
timestamp 1680363874
transform 1 0 3136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1680363874
transform 1 0 3144 0 1 3170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1680363874
transform 1 0 3152 0 1 3170
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1680363874
transform 1 0 3160 0 1 3170
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1680363874
transform 1 0 3168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1680363874
transform 1 0 3176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1680363874
transform 1 0 3184 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_102
timestamp 1680363874
transform -1 0 3224 0 1 3170
box -8 -3 34 105
use FILL  FILL_3420
timestamp 1680363874
transform 1 0 3224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1680363874
transform 1 0 3232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1680363874
transform 1 0 3240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1680363874
transform 1 0 3248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1680363874
transform 1 0 3256 0 1 3170
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1680363874
transform 1 0 3264 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_254
timestamp 1680363874
transform 1 0 3272 0 1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1680363874
transform -1 0 3384 0 1 3170
box -8 -3 104 105
use FILL  FILL_3436
timestamp 1680363874
transform 1 0 3384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1680363874
transform 1 0 3392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1680363874
transform 1 0 3400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1680363874
transform 1 0 3408 0 1 3170
box -8 -3 16 105
use AND2X2  AND2X2_8
timestamp 1680363874
transform 1 0 3416 0 1 3170
box -8 -3 40 105
use FILL  FILL_3451
timestamp 1680363874
transform 1 0 3448 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3031
timestamp 1680363874
transform 1 0 3468 0 1 3175
box -3 -3 3 3
use FILL  FILL_3455
timestamp 1680363874
transform 1 0 3456 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_11
timestamp 1680363874
transform 1 0 3464 0 1 3170
box -5 -3 28 105
use FILL  FILL_3457
timestamp 1680363874
transform 1 0 3488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1680363874
transform 1 0 3496 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3032
timestamp 1680363874
transform 1 0 3516 0 1 3175
box -3 -3 3 3
use FILL  FILL_3459
timestamp 1680363874
transform 1 0 3504 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_12
timestamp 1680363874
transform 1 0 3512 0 1 3170
box -5 -3 28 105
use FILL  FILL_3460
timestamp 1680363874
transform 1 0 3536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1680363874
transform 1 0 3544 0 1 3170
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1680363874
transform 1 0 3552 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_30
timestamp 1680363874
transform -1 0 3584 0 1 3170
box -8 -3 32 105
use FILL  FILL_3469
timestamp 1680363874
transform 1 0 3584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1680363874
transform 1 0 3592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1680363874
transform 1 0 3600 0 1 3170
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1680363874
transform 1 0 3608 0 1 3170
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1680363874
transform 1 0 3616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1680363874
transform 1 0 3624 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3033
timestamp 1680363874
transform 1 0 3660 0 1 3175
box -3 -3 3 3
use OAI21X1  OAI21X1_103
timestamp 1680363874
transform -1 0 3664 0 1 3170
box -8 -3 34 105
use FILL  FILL_3480
timestamp 1680363874
transform 1 0 3664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1680363874
transform 1 0 3672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1680363874
transform 1 0 3680 0 1 3170
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1680363874
transform 1 0 3688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1680363874
transform 1 0 3696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1680363874
transform 1 0 3704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1680363874
transform 1 0 3712 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_204
timestamp 1680363874
transform 1 0 3720 0 1 3170
box -8 -3 46 105
use FILL  FILL_3487
timestamp 1680363874
transform 1 0 3760 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3034
timestamp 1680363874
transform 1 0 3780 0 1 3175
box -3 -3 3 3
use FILL  FILL_3488
timestamp 1680363874
transform 1 0 3768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1680363874
transform 1 0 3776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1680363874
transform 1 0 3784 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_235
timestamp 1680363874
transform -1 0 3888 0 1 3170
box -8 -3 104 105
use FILL  FILL_3497
timestamp 1680363874
transform 1 0 3888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1680363874
transform 1 0 3896 0 1 3170
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1680363874
transform 1 0 3904 0 1 3170
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1680363874
transform 1 0 3912 0 1 3170
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1680363874
transform 1 0 3920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1680363874
transform 1 0 3928 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_205
timestamp 1680363874
transform -1 0 3976 0 1 3170
box -8 -3 46 105
use FILL  FILL_3513
timestamp 1680363874
transform 1 0 3976 0 1 3170
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1680363874
transform 1 0 3984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1680363874
transform 1 0 3992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1680363874
transform 1 0 4000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1680363874
transform 1 0 4008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1680363874
transform 1 0 4016 0 1 3170
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1680363874
transform 1 0 4024 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_32
timestamp 1680363874
transform -1 0 4056 0 1 3170
box -8 -3 32 105
use FILL  FILL_3525
timestamp 1680363874
transform 1 0 4056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1680363874
transform 1 0 4064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1680363874
transform 1 0 4072 0 1 3170
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1680363874
transform 1 0 4080 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1680363874
transform -1 0 4184 0 1 3170
box -8 -3 104 105
use FILL  FILL_3535
timestamp 1680363874
transform 1 0 4184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1680363874
transform 1 0 4192 0 1 3170
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1680363874
transform 1 0 4200 0 1 3170
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1680363874
transform 1 0 4208 0 1 3170
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1680363874
transform 1 0 4216 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_33
timestamp 1680363874
transform -1 0 4248 0 1 3170
box -8 -3 32 105
use FILL  FILL_3540
timestamp 1680363874
transform 1 0 4248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1680363874
transform 1 0 4256 0 1 3170
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1680363874
transform 1 0 4264 0 1 3170
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1680363874
transform 1 0 4272 0 1 3170
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1680363874
transform 1 0 4280 0 1 3170
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1680363874
transform 1 0 4288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1680363874
transform 1 0 4296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1680363874
transform 1 0 4304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1680363874
transform 1 0 4312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1680363874
transform 1 0 4320 0 1 3170
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1680363874
transform 1 0 4328 0 1 3170
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1680363874
transform 1 0 4336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1680363874
transform 1 0 4344 0 1 3170
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1680363874
transform 1 0 4352 0 1 3170
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1680363874
transform 1 0 4360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1680363874
transform 1 0 4368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1680363874
transform 1 0 4376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1680363874
transform 1 0 4384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1680363874
transform 1 0 4392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1680363874
transform 1 0 4400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1680363874
transform 1 0 4408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1680363874
transform 1 0 4416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1680363874
transform 1 0 4424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1680363874
transform 1 0 4432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1680363874
transform 1 0 4440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1680363874
transform 1 0 4448 0 1 3170
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1680363874
transform 1 0 4456 0 1 3170
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1680363874
transform 1 0 4464 0 1 3170
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1680363874
transform 1 0 4472 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_207
timestamp 1680363874
transform 1 0 4480 0 1 3170
box -8 -3 46 105
use FILL  FILL_3590
timestamp 1680363874
transform 1 0 4520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1680363874
transform 1 0 4528 0 1 3170
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1680363874
transform 1 0 4536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1680363874
transform 1 0 4544 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_237
timestamp 1680363874
transform 1 0 4552 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_258
timestamp 1680363874
transform 1 0 4648 0 1 3170
box -9 -3 26 105
use FILL  FILL_3594
timestamp 1680363874
transform 1 0 4664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1680363874
transform 1 0 4672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1680363874
transform 1 0 4680 0 1 3170
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1680363874
transform 1 0 4688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1680363874
transform 1 0 4696 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1680363874
transform -1 0 4800 0 1 3170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_31
timestamp 1680363874
transform 1 0 4827 0 1 3170
box -10 -3 10 3
use M2_M1  M2_M1_3410
timestamp 1680363874
transform 1 0 84 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1680363874
transform 1 0 132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1680363874
transform 1 0 196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1680363874
transform 1 0 220 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3160
timestamp 1680363874
transform 1 0 220 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3411
timestamp 1680363874
transform 1 0 236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1680363874
transform 1 0 244 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3129
timestamp 1680363874
transform 1 0 244 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1680363874
transform 1 0 236 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3600
timestamp 1680363874
transform 1 0 244 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1680363874
transform 1 0 284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1680363874
transform 1 0 276 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3147
timestamp 1680363874
transform 1 0 284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1680363874
transform 1 0 276 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1680363874
transform 1 0 300 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1680363874
transform 1 0 332 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1680363874
transform 1 0 324 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3413
timestamp 1680363874
transform 1 0 300 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3107
timestamp 1680363874
transform 1 0 308 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3414
timestamp 1680363874
transform 1 0 316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1680363874
transform 1 0 308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1680363874
transform 1 0 324 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3148
timestamp 1680363874
transform 1 0 332 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1680363874
transform 1 0 348 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3415
timestamp 1680363874
transform 1 0 348 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1680363874
transform 1 0 356 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3071
timestamp 1680363874
transform 1 0 388 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3417
timestamp 1680363874
transform 1 0 380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1680363874
transform 1 0 388 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3130
timestamp 1680363874
transform 1 0 380 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3603
timestamp 1680363874
transform 1 0 380 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1680363874
transform 1 0 396 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1680363874
transform 1 0 436 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3058
timestamp 1680363874
transform 1 0 452 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1680363874
transform 1 0 444 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1680363874
transform 1 0 468 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3420
timestamp 1680363874
transform 1 0 468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1680363874
transform 1 0 452 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1680363874
transform 1 0 460 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3162
timestamp 1680363874
transform 1 0 460 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1680363874
transform 1 0 484 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3508
timestamp 1680363874
transform 1 0 492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1680363874
transform 1 0 516 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3163
timestamp 1680363874
transform 1 0 516 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1680363874
transform 1 0 524 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3421
timestamp 1680363874
transform 1 0 540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1680363874
transform 1 0 556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1680363874
transform 1 0 604 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3109
timestamp 1680363874
transform 1 0 612 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3605
timestamp 1680363874
transform 1 0 636 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3164
timestamp 1680363874
transform 1 0 636 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1680363874
transform 1 0 660 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3424
timestamp 1680363874
transform 1 0 660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1680363874
transform 1 0 652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1680363874
transform 1 0 676 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1680363874
transform 1 0 724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1680363874
transform 1 0 732 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3038
timestamp 1680363874
transform 1 0 740 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3425
timestamp 1680363874
transform 1 0 740 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3165
timestamp 1680363874
transform 1 0 732 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3426
timestamp 1680363874
transform 1 0 756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1680363874
transform 1 0 844 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1680363874
transform 1 0 868 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1680363874
transform 1 0 764 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1680363874
transform 1 0 812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1680363874
transform 1 0 860 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3149
timestamp 1680363874
transform 1 0 892 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3429
timestamp 1680363874
transform 1 0 924 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3110
timestamp 1680363874
transform 1 0 940 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3430
timestamp 1680363874
transform 1 0 972 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1680363874
transform 1 0 940 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1680363874
transform 1 0 948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1680363874
transform 1 0 964 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3150
timestamp 1680363874
transform 1 0 964 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3517
timestamp 1680363874
transform 1 0 980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1680363874
transform 1 0 1004 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3151
timestamp 1680363874
transform 1 0 1004 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1680363874
transform 1 0 1052 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3431
timestamp 1680363874
transform 1 0 1036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1680363874
transform 1 0 1044 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1680363874
transform 1 0 1028 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3152
timestamp 1680363874
transform 1 0 1036 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1680363874
transform 1 0 1084 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3433
timestamp 1680363874
transform 1 0 1068 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3111
timestamp 1680363874
transform 1 0 1076 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3520
timestamp 1680363874
transform 1 0 1060 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1680363874
transform 1 0 1076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1680363874
transform 1 0 1092 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3074
timestamp 1680363874
transform 1 0 1116 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1680363874
transform 1 0 1116 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1680363874
transform 1 0 1244 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1680363874
transform 1 0 1132 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1680363874
transform 1 0 1212 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1680363874
transform 1 0 1228 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3435
timestamp 1680363874
transform 1 0 1140 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3076
timestamp 1680363874
transform 1 0 1252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1680363874
transform 1 0 1284 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3436
timestamp 1680363874
transform 1 0 1236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1680363874
transform 1 0 1252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1680363874
transform 1 0 1164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1680363874
transform 1 0 1220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1680363874
transform 1 0 1228 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3154
timestamp 1680363874
transform 1 0 1140 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1680363874
transform 1 0 1212 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3525
timestamp 1680363874
transform 1 0 1284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1680363874
transform 1 0 1332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1680363874
transform 1 0 1348 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3156
timestamp 1680363874
transform 1 0 1252 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3607
timestamp 1680363874
transform 1 0 1340 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3195
timestamp 1680363874
transform 1 0 1268 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3613
timestamp 1680363874
transform 1 0 1356 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1680363874
transform 1 0 1372 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1680363874
transform 1 0 1380 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3040
timestamp 1680363874
transform 1 0 1396 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3438
timestamp 1680363874
transform 1 0 1420 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3132
timestamp 1680363874
transform 1 0 1420 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3610
timestamp 1680363874
transform 1 0 1412 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1680363874
transform 1 0 1396 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1680363874
transform 1 0 1436 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1680363874
transform 1 0 1476 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1680363874
transform 1 0 1468 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3166
timestamp 1680363874
transform 1 0 1468 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3529
timestamp 1680363874
transform 1 0 1500 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3167
timestamp 1680363874
transform 1 0 1500 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1680363874
transform 1 0 1580 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1680363874
transform 1 0 1604 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1680363874
transform 1 0 1572 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3440
timestamp 1680363874
transform 1 0 1524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1680363874
transform 1 0 1572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1680363874
transform 1 0 1604 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3168
timestamp 1680363874
transform 1 0 1524 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1680363874
transform 1 0 1628 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1680363874
transform 1 0 1692 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3441
timestamp 1680363874
transform 1 0 1628 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3112
timestamp 1680363874
transform 1 0 1676 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1680363874
transform 1 0 1700 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3532
timestamp 1680363874
transform 1 0 1676 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3169
timestamp 1680363874
transform 1 0 1628 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1680363874
transform 1 0 1676 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1680363874
transform 1 0 1660 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1680363874
transform 1 0 1724 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1680363874
transform 1 0 1716 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1680363874
transform 1 0 1748 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3533
timestamp 1680363874
transform 1 0 1748 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1680363874
transform 1 0 1756 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3043
timestamp 1680363874
transform 1 0 1796 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3442
timestamp 1680363874
transform 1 0 1796 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3115
timestamp 1680363874
transform 1 0 1804 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3443
timestamp 1680363874
transform 1 0 1812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1680363874
transform 1 0 1828 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1680363874
transform 1 0 1804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1680363874
transform 1 0 1820 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3170
timestamp 1680363874
transform 1 0 1796 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1680363874
transform 1 0 1820 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1680363874
transform 1 0 1804 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1680363874
transform 1 0 1844 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1680363874
transform 1 0 1868 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1680363874
transform 1 0 1876 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1680363874
transform 1 0 1916 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3445
timestamp 1680363874
transform 1 0 1876 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1680363874
transform 1 0 1892 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1680363874
transform 1 0 1908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1680363874
transform 1 0 1916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1680363874
transform 1 0 1884 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1680363874
transform 1 0 1908 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3173
timestamp 1680363874
transform 1 0 1900 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1680363874
transform 1 0 1908 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1680363874
transform 1 0 1924 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3539
timestamp 1680363874
transform 1 0 1948 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3116
timestamp 1680363874
transform 1 0 1972 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1680363874
transform 1 0 2020 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1680363874
transform 1 0 2012 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3449
timestamp 1680363874
transform 1 0 1980 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3117
timestamp 1680363874
transform 1 0 1988 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3450
timestamp 1680363874
transform 1 0 1996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1680363874
transform 1 0 2012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1680363874
transform 1 0 2004 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3174
timestamp 1680363874
transform 1 0 2004 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1680363874
transform 1 0 2036 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1680363874
transform 1 0 2076 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1680363874
transform 1 0 2092 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1680363874
transform 1 0 2116 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1680363874
transform 1 0 2116 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3452
timestamp 1680363874
transform 1 0 2084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1680363874
transform 1 0 2100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1680363874
transform 1 0 2116 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1680363874
transform 1 0 2076 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3133
timestamp 1680363874
transform 1 0 2084 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3542
timestamp 1680363874
transform 1 0 2108 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3134
timestamp 1680363874
transform 1 0 2116 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1680363874
transform 1 0 2108 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3543
timestamp 1680363874
transform 1 0 2132 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3177
timestamp 1680363874
transform 1 0 2132 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3455
timestamp 1680363874
transform 1 0 2172 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3119
timestamp 1680363874
transform 1 0 2196 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3544
timestamp 1680363874
transform 1 0 2188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1680363874
transform 1 0 2196 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3178
timestamp 1680363874
transform 1 0 2204 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1680363874
transform 1 0 2220 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1680363874
transform 1 0 2252 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3456
timestamp 1680363874
transform 1 0 2220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1680363874
transform 1 0 2236 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3120
timestamp 1680363874
transform 1 0 2244 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3458
timestamp 1680363874
transform 1 0 2252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1680363874
transform 1 0 2244 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1680363874
transform 1 0 2260 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3179
timestamp 1680363874
transform 1 0 2276 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1680363874
transform 1 0 2308 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3459
timestamp 1680363874
transform 1 0 2388 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3049
timestamp 1680363874
transform 1 0 2404 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1680363874
transform 1 0 2460 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1680363874
transform 1 0 2476 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3460
timestamp 1680363874
transform 1 0 2428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1680363874
transform 1 0 2476 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3180
timestamp 1680363874
transform 1 0 2428 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1680363874
transform 1 0 2468 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3461
timestamp 1680363874
transform 1 0 2556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1680363874
transform 1 0 2564 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3182
timestamp 1680363874
transform 1 0 2564 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1680363874
transform 1 0 2580 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3550
timestamp 1680363874
transform 1 0 2580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3210
timestamp 1680363874
transform 1 0 2596 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1680363874
transform 1 0 2628 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1680363874
transform 1 0 2620 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1680363874
transform 1 0 2636 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3462
timestamp 1680363874
transform 1 0 2620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1680363874
transform 1 0 2636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1680363874
transform 1 0 2644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1680363874
transform 1 0 2628 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3183
timestamp 1680363874
transform 1 0 2628 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1680363874
transform 1 0 2652 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1680363874
transform 1 0 2644 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3552
timestamp 1680363874
transform 1 0 2652 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3091
timestamp 1680363874
transform 1 0 2740 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3465
timestamp 1680363874
transform 1 0 2724 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1680363874
transform 1 0 2740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1680363874
transform 1 0 2732 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3124
timestamp 1680363874
transform 1 0 2748 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3467
timestamp 1680363874
transform 1 0 2756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1680363874
transform 1 0 2748 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3092
timestamp 1680363874
transform 1 0 2836 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3468
timestamp 1680363874
transform 1 0 2804 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1680363874
transform 1 0 2820 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1680363874
transform 1 0 2836 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1680363874
transform 1 0 2812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1680363874
transform 1 0 2828 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3136
timestamp 1680363874
transform 1 0 2836 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1680363874
transform 1 0 2812 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3471
timestamp 1680363874
transform 1 0 2884 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3093
timestamp 1680363874
transform 1 0 2908 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3557
timestamp 1680363874
transform 1 0 2892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1680363874
transform 1 0 2908 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3184
timestamp 1680363874
transform 1 0 2884 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1680363874
transform 1 0 2916 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1680363874
transform 1 0 2916 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3611
timestamp 1680363874
transform 1 0 2932 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1680363874
transform 1 0 2956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1680363874
transform 1 0 2988 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3051
timestamp 1680363874
transform 1 0 3076 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3560
timestamp 1680363874
transform 1 0 3092 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1680363874
transform 1 0 3100 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3212
timestamp 1680363874
transform 1 0 3100 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3562
timestamp 1680363874
transform 1 0 3116 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3185
timestamp 1680363874
transform 1 0 3124 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1680363874
transform 1 0 3132 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1680363874
transform 1 0 3132 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1680363874
transform 1 0 3148 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3473
timestamp 1680363874
transform 1 0 3148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1680363874
transform 1 0 3156 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1680363874
transform 1 0 3180 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3095
timestamp 1680363874
transform 1 0 3188 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3475
timestamp 1680363874
transform 1 0 3188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1680363874
transform 1 0 3188 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3186
timestamp 1680363874
transform 1 0 3188 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3565
timestamp 1680363874
transform 1 0 3212 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3052
timestamp 1680363874
transform 1 0 3260 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1680363874
transform 1 0 3252 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1680363874
transform 1 0 3292 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3476
timestamp 1680363874
transform 1 0 3276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1680363874
transform 1 0 3292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1680363874
transform 1 0 3268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1680363874
transform 1 0 3284 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3138
timestamp 1680363874
transform 1 0 3292 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3568
timestamp 1680363874
transform 1 0 3300 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3188
timestamp 1680363874
transform 1 0 3300 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3569
timestamp 1680363874
transform 1 0 3316 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3125
timestamp 1680363874
transform 1 0 3356 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1680363874
transform 1 0 3388 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3570
timestamp 1680363874
transform 1 0 3380 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3062
timestamp 1680363874
transform 1 0 3404 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3478
timestamp 1680363874
transform 1 0 3404 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3063
timestamp 1680363874
transform 1 0 3420 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1680363874
transform 1 0 3428 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3479
timestamp 1680363874
transform 1 0 3428 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3214
timestamp 1680363874
transform 1 0 3420 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1680363874
transform 1 0 3436 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3480
timestamp 1680363874
transform 1 0 3452 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3139
timestamp 1680363874
transform 1 0 3452 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3571
timestamp 1680363874
transform 1 0 3460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1680363874
transform 1 0 3468 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3097
timestamp 1680363874
transform 1 0 3508 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3481
timestamp 1680363874
transform 1 0 3492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1680363874
transform 1 0 3516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1680363874
transform 1 0 3508 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1680363874
transform 1 0 3524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1680363874
transform 1 0 3532 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3189
timestamp 1680363874
transform 1 0 3524 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1680363874
transform 1 0 3564 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1680363874
transform 1 0 3580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1680363874
transform 1 0 3620 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3483
timestamp 1680363874
transform 1 0 3604 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3140
timestamp 1680363874
transform 1 0 3604 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3484
timestamp 1680363874
transform 1 0 3628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1680363874
transform 1 0 3636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1680363874
transform 1 0 3620 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3216
timestamp 1680363874
transform 1 0 3636 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3576
timestamp 1680363874
transform 1 0 3652 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3203
timestamp 1680363874
transform 1 0 3652 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1680363874
transform 1 0 3732 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1680363874
transform 1 0 3716 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1680363874
transform 1 0 3732 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1680363874
transform 1 0 3700 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3486
timestamp 1680363874
transform 1 0 3764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1680363874
transform 1 0 3676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1680363874
transform 1 0 3684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1680363874
transform 1 0 3716 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3204
timestamp 1680363874
transform 1 0 3676 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1680363874
transform 1 0 3700 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1680363874
transform 1 0 3716 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1680363874
transform 1 0 3764 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1680363874
transform 1 0 3716 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3487
timestamp 1680363874
transform 1 0 3780 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3192
timestamp 1680363874
transform 1 0 3780 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1680363874
transform 1 0 3820 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3580
timestamp 1680363874
transform 1 0 3812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1680363874
transform 1 0 3820 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3218
timestamp 1680363874
transform 1 0 3828 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3405
timestamp 1680363874
transform 1 0 3860 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1680363874
transform 1 0 3860 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1680363874
transform 1 0 3868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1680363874
transform 1 0 3940 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3066
timestamp 1680363874
transform 1 0 3956 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1680363874
transform 1 0 3956 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3406
timestamp 1680363874
transform 1 0 3964 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1680363874
transform 1 0 3956 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1680363874
transform 1 0 3964 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1680363874
transform 1 0 3996 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_3101
timestamp 1680363874
transform 1 0 4012 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3584
timestamp 1680363874
transform 1 0 4004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1680363874
transform 1 0 4020 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1680363874
transform 1 0 4036 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3157
timestamp 1680363874
transform 1 0 4020 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1680363874
transform 1 0 4068 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3408
timestamp 1680363874
transform 1 0 4108 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1680363874
transform 1 0 4132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1680363874
transform 1 0 4140 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3103
timestamp 1680363874
transform 1 0 4172 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3491
timestamp 1680363874
transform 1 0 4172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1680363874
transform 1 0 4204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1680363874
transform 1 0 4236 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1680363874
transform 1 0 4236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1680363874
transform 1 0 4228 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3141
timestamp 1680363874
transform 1 0 4244 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1680363874
transform 1 0 4316 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3493
timestamp 1680363874
transform 1 0 4292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1680363874
transform 1 0 4308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1680363874
transform 1 0 4316 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3158
timestamp 1680363874
transform 1 0 4292 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1680363874
transform 1 0 4356 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3495
timestamp 1680363874
transform 1 0 4348 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3142
timestamp 1680363874
transform 1 0 4348 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1680363874
transform 1 0 4364 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3496
timestamp 1680363874
transform 1 0 4364 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3143
timestamp 1680363874
transform 1 0 4388 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3592
timestamp 1680363874
transform 1 0 4396 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1680363874
transform 1 0 4444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1680363874
transform 1 0 4452 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3159
timestamp 1680363874
transform 1 0 4444 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1680363874
transform 1 0 4356 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1680363874
transform 1 0 4412 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1680363874
transform 1 0 4492 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1680363874
transform 1 0 4540 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3497
timestamp 1680363874
transform 1 0 4540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1680363874
transform 1 0 4508 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3144
timestamp 1680363874
transform 1 0 4540 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1680363874
transform 1 0 4572 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3498
timestamp 1680363874
transform 1 0 4572 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3127
timestamp 1680363874
transform 1 0 4620 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1680363874
transform 1 0 4572 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1680363874
transform 1 0 4660 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3596
timestamp 1680363874
transform 1 0 4620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1680363874
transform 1 0 4652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1680363874
transform 1 0 4772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1680363874
transform 1 0 4692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1680363874
transform 1 0 4732 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3207
timestamp 1680363874
transform 1 0 4812 0 1 3095
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_32
timestamp 1680363874
transform 1 0 24 0 1 3070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_219
timestamp 1680363874
transform 1 0 72 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3095
timestamp 1680363874
transform 1 0 168 0 -1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_21
timestamp 1680363874
transform 1 0 176 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3096
timestamp 1680363874
transform 1 0 200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1680363874
transform 1 0 208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1680363874
transform 1 0 216 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_230
timestamp 1680363874
transform -1 0 240 0 -1 3170
box -9 -3 26 105
use OAI21X1  OAI21X1_88
timestamp 1680363874
transform -1 0 272 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3110
timestamp 1680363874
transform 1 0 272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1680363874
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1680363874
transform 1 0 288 0 -1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_24
timestamp 1680363874
transform -1 0 320 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1680363874
transform -1 0 344 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3113
timestamp 1680363874
transform 1 0 344 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_90
timestamp 1680363874
transform 1 0 352 0 -1 3170
box -8 -3 34 105
use INVX2  INVX2_231
timestamp 1680363874
transform 1 0 384 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3124
timestamp 1680363874
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1680363874
transform 1 0 408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1680363874
transform 1 0 416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1680363874
transform 1 0 424 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_5
timestamp 1680363874
transform -1 0 456 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3128
timestamp 1680363874
transform 1 0 456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1680363874
transform 1 0 464 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_232
timestamp 1680363874
transform 1 0 472 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3130
timestamp 1680363874
transform 1 0 488 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_233
timestamp 1680363874
transform -1 0 512 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3131
timestamp 1680363874
transform 1 0 512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1680363874
transform 1 0 520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1680363874
transform 1 0 528 0 -1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_27
timestamp 1680363874
transform -1 0 560 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3136
timestamp 1680363874
transform 1 0 560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1680363874
transform 1 0 568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1680363874
transform 1 0 576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1680363874
transform 1 0 584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1680363874
transform 1 0 592 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_93
timestamp 1680363874
transform 1 0 600 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3147
timestamp 1680363874
transform 1 0 632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1680363874
transform 1 0 640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1680363874
transform 1 0 648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1680363874
transform 1 0 656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1680363874
transform 1 0 664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1680363874
transform 1 0 672 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_94
timestamp 1680363874
transform 1 0 680 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3159
timestamp 1680363874
transform 1 0 712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1680363874
transform 1 0 720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1680363874
transform 1 0 728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1680363874
transform 1 0 736 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_236
timestamp 1680363874
transform -1 0 760 0 -1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_220
timestamp 1680363874
transform -1 0 856 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_237
timestamp 1680363874
transform -1 0 872 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3174
timestamp 1680363874
transform 1 0 872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1680363874
transform 1 0 880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1680363874
transform 1 0 888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1680363874
transform 1 0 896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1680363874
transform 1 0 904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1680363874
transform 1 0 912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1680363874
transform 1 0 920 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_238
timestamp 1680363874
transform 1 0 928 0 -1 3170
box -9 -3 26 105
use AND2X2  AND2X2_5
timestamp 1680363874
transform -1 0 976 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3192
timestamp 1680363874
transform 1 0 976 0 -1 3170
box -8 -3 16 105
use AND2X2  AND2X2_6
timestamp 1680363874
transform -1 0 1016 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3193
timestamp 1680363874
transform 1 0 1016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1680363874
transform 1 0 1024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1680363874
transform 1 0 1032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1680363874
transform 1 0 1040 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_189
timestamp 1680363874
transform 1 0 1048 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3201
timestamp 1680363874
transform 1 0 1088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1680363874
transform 1 0 1096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1680363874
transform 1 0 1104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1680363874
transform 1 0 1112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1680363874
transform 1 0 1120 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1680363874
transform 1 0 1128 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_241
timestamp 1680363874
transform -1 0 1240 0 -1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1680363874
transform 1 0 1240 0 -1 3170
box -8 -3 104 105
use NAND3X1  NAND3X1_0
timestamp 1680363874
transform 1 0 1336 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3228
timestamp 1680363874
transform 1 0 1368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1680363874
transform 1 0 1376 0 -1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1680363874
transform -1 0 1416 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3230
timestamp 1680363874
transform 1 0 1416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1680363874
transform 1 0 1424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1680363874
transform 1 0 1432 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_6
timestamp 1680363874
transform -1 0 1464 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3245
timestamp 1680363874
transform 1 0 1464 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3219
timestamp 1680363874
transform 1 0 1500 0 1 3075
box -3 -3 3 3
use BUFX2  BUFX2_7
timestamp 1680363874
transform -1 0 1496 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3246
timestamp 1680363874
transform 1 0 1496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1680363874
transform 1 0 1504 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1680363874
transform 1 0 1512 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3248
timestamp 1680363874
transform 1 0 1608 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1680363874
transform 1 0 1616 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3249
timestamp 1680363874
transform 1 0 1712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1680363874
transform 1 0 1720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1680363874
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_244
timestamp 1680363874
transform 1 0 1736 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3257
timestamp 1680363874
transform 1 0 1752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1680363874
transform 1 0 1760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1680363874
transform 1 0 1768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1680363874
transform 1 0 1776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1680363874
transform 1 0 1784 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_195
timestamp 1680363874
transform 1 0 1792 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3262
timestamp 1680363874
transform 1 0 1832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1680363874
transform 1 0 1840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1680363874
transform 1 0 1848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1680363874
transform 1 0 1856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1680363874
transform 1 0 1864 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_196
timestamp 1680363874
transform -1 0 1912 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3267
timestamp 1680363874
transform 1 0 1912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1680363874
transform 1 0 1920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1680363874
transform 1 0 1928 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_245
timestamp 1680363874
transform 1 0 1936 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3270
timestamp 1680363874
transform 1 0 1952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1680363874
transform 1 0 1960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1680363874
transform 1 0 1968 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_197
timestamp 1680363874
transform 1 0 1976 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3273
timestamp 1680363874
transform 1 0 2016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1680363874
transform 1 0 2024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1680363874
transform 1 0 2032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1680363874
transform 1 0 2040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1680363874
transform 1 0 2048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1680363874
transform 1 0 2056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1680363874
transform 1 0 2064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1680363874
transform 1 0 2072 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_199
timestamp 1680363874
transform 1 0 2080 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3285
timestamp 1680363874
transform 1 0 2120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1680363874
transform 1 0 2128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1680363874
transform 1 0 2136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1680363874
transform 1 0 2144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1680363874
transform 1 0 2152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1680363874
transform 1 0 2160 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_246
timestamp 1680363874
transform 1 0 2168 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3296
timestamp 1680363874
transform 1 0 2184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1680363874
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1680363874
transform 1 0 2200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1680363874
transform 1 0 2208 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3220
timestamp 1680363874
transform 1 0 2260 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_200
timestamp 1680363874
transform 1 0 2216 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3302
timestamp 1680363874
transform 1 0 2256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1680363874
transform 1 0 2264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1680363874
transform 1 0 2272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1680363874
transform 1 0 2280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1680363874
transform 1 0 2288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1680363874
transform 1 0 2296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1680363874
transform 1 0 2304 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3221
timestamp 1680363874
transform 1 0 2332 0 1 3075
box -3 -3 3 3
use BUFX2  BUFX2_9
timestamp 1680363874
transform 1 0 2312 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3313
timestamp 1680363874
transform 1 0 2336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1680363874
transform 1 0 2344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1680363874
transform 1 0 2352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1680363874
transform 1 0 2360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1680363874
transform 1 0 2368 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3222
timestamp 1680363874
transform 1 0 2388 0 1 3075
box -3 -3 3 3
use FILL  FILL_3320
timestamp 1680363874
transform 1 0 2376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1680363874
transform 1 0 2384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1680363874
transform 1 0 2392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1680363874
transform 1 0 2400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1680363874
transform 1 0 2408 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1680363874
transform 1 0 2416 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3335
timestamp 1680363874
transform 1 0 2512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1680363874
transform 1 0 2520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1680363874
transform 1 0 2528 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_248
timestamp 1680363874
transform 1 0 2536 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3338
timestamp 1680363874
transform 1 0 2552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1680363874
transform 1 0 2560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1680363874
transform 1 0 2568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1680363874
transform 1 0 2576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1680363874
transform 1 0 2584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1680363874
transform 1 0 2592 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_201
timestamp 1680363874
transform 1 0 2600 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3352
timestamp 1680363874
transform 1 0 2640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1680363874
transform 1 0 2648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1680363874
transform 1 0 2656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1680363874
transform 1 0 2664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1680363874
transform 1 0 2672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1680363874
transform 1 0 2680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1680363874
transform 1 0 2688 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1680363874
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_202
timestamp 1680363874
transform 1 0 2704 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3360
timestamp 1680363874
transform 1 0 2744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1680363874
transform 1 0 2752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1680363874
transform 1 0 2760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1680363874
transform 1 0 2768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1680363874
transform 1 0 2776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1680363874
transform 1 0 2784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1680363874
transform 1 0 2792 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_203
timestamp 1680363874
transform 1 0 2800 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3371
timestamp 1680363874
transform 1 0 2840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1680363874
transform 1 0 2848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1680363874
transform 1 0 2856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1680363874
transform 1 0 2864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1680363874
transform 1 0 2872 0 -1 3170
box -8 -3 16 105
use AND2X2  AND2X2_7
timestamp 1680363874
transform 1 0 2880 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3380
timestamp 1680363874
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1680363874
transform 1 0 2920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1680363874
transform 1 0 2928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1680363874
transform 1 0 2936 0 -1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1680363874
transform -1 0 2968 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3387
timestamp 1680363874
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1680363874
transform 1 0 2976 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_252
timestamp 1680363874
transform 1 0 2984 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3394
timestamp 1680363874
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1680363874
transform 1 0 3008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1680363874
transform 1 0 3016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1680363874
transform 1 0 3024 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_253
timestamp 1680363874
transform 1 0 3032 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3398
timestamp 1680363874
transform 1 0 3048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1680363874
transform 1 0 3056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1680363874
transform 1 0 3064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1680363874
transform 1 0 3072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1680363874
transform 1 0 3080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1680363874
transform 1 0 3088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1680363874
transform 1 0 3096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1680363874
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1680363874
transform 1 0 3112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1680363874
transform 1 0 3120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1680363874
transform 1 0 3128 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_128
timestamp 1680363874
transform 1 0 3136 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3418
timestamp 1680363874
transform 1 0 3176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1680363874
transform 1 0 3184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1680363874
transform 1 0 3192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1680363874
transform 1 0 3200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1680363874
transform 1 0 3208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1680363874
transform 1 0 3216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1680363874
transform 1 0 3224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1680363874
transform 1 0 3232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1680363874
transform 1 0 3240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1680363874
transform 1 0 3248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1680363874
transform 1 0 3256 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_129
timestamp 1680363874
transform 1 0 3264 0 -1 3170
box -8 -3 46 105
use M3_M2  M3_M2_3223
timestamp 1680363874
transform 1 0 3316 0 1 3075
box -3 -3 3 3
use FILL  FILL_3439
timestamp 1680363874
transform 1 0 3304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1680363874
transform 1 0 3312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1680363874
transform 1 0 3320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1680363874
transform 1 0 3328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1680363874
transform 1 0 3336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1680363874
transform 1 0 3344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1680363874
transform 1 0 3352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1680363874
transform 1 0 3360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1680363874
transform 1 0 3368 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_10
timestamp 1680363874
transform 1 0 3376 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3448
timestamp 1680363874
transform 1 0 3400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1680363874
transform 1 0 3408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1680363874
transform 1 0 3416 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_255
timestamp 1680363874
transform 1 0 3424 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3453
timestamp 1680363874
transform 1 0 3440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1680363874
transform 1 0 3448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1680363874
transform 1 0 3456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1680363874
transform 1 0 3464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1680363874
transform 1 0 3472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1680363874
transform 1 0 3480 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_130
timestamp 1680363874
transform 1 0 3488 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3464
timestamp 1680363874
transform 1 0 3528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1680363874
transform 1 0 3536 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1680363874
transform 1 0 3544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1680363874
transform 1 0 3552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1680363874
transform 1 0 3560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1680363874
transform 1 0 3568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1680363874
transform 1 0 3576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1680363874
transform 1 0 3584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1680363874
transform 1 0 3592 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_104
timestamp 1680363874
transform -1 0 3632 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3491
timestamp 1680363874
transform 1 0 3632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1680363874
transform 1 0 3640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1680363874
transform 1 0 3648 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_256
timestamp 1680363874
transform 1 0 3656 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3494
timestamp 1680363874
transform 1 0 3672 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_234
timestamp 1680363874
transform -1 0 3776 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3495
timestamp 1680363874
transform 1 0 3776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1680363874
transform 1 0 3784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1680363874
transform 1 0 3792 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_257
timestamp 1680363874
transform 1 0 3800 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3500
timestamp 1680363874
transform 1 0 3816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1680363874
transform 1 0 3824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1680363874
transform 1 0 3832 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_31
timestamp 1680363874
transform -1 0 3864 0 -1 3170
box -8 -3 32 105
use BUFX2  BUFX2_13
timestamp 1680363874
transform 1 0 3864 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3503
timestamp 1680363874
transform 1 0 3888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1680363874
transform 1 0 3896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1680363874
transform 1 0 3904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1680363874
transform 1 0 3912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1680363874
transform 1 0 3920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1680363874
transform 1 0 3928 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_14
timestamp 1680363874
transform 1 0 3936 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3515
timestamp 1680363874
transform 1 0 3960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1680363874
transform 1 0 3968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1680363874
transform 1 0 3976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1680363874
transform 1 0 3984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1680363874
transform 1 0 3992 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_131
timestamp 1680363874
transform -1 0 4040 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3527
timestamp 1680363874
transform 1 0 4040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1680363874
transform 1 0 4048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1680363874
transform 1 0 4056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1680363874
transform 1 0 4064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1680363874
transform 1 0 4072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1680363874
transform 1 0 4080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1680363874
transform 1 0 4088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1680363874
transform 1 0 4096 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_34
timestamp 1680363874
transform 1 0 4104 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3544
timestamp 1680363874
transform 1 0 4128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1680363874
transform 1 0 4136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1680363874
transform 1 0 4144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1680363874
transform 1 0 4152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1680363874
transform 1 0 4160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1680363874
transform 1 0 4168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1680363874
transform 1 0 4176 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_132
timestamp 1680363874
transform -1 0 4224 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3551
timestamp 1680363874
transform 1 0 4224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1680363874
transform 1 0 4232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1680363874
transform 1 0 4240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1680363874
transform 1 0 4248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1680363874
transform 1 0 4256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1680363874
transform 1 0 4264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1680363874
transform 1 0 4272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1680363874
transform 1 0 4280 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_206
timestamp 1680363874
transform 1 0 4288 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3569
timestamp 1680363874
transform 1 0 4328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1680363874
transform 1 0 4336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1680363874
transform 1 0 4344 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1680363874
transform 1 0 4352 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3595
timestamp 1680363874
transform 1 0 4448 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1680363874
transform -1 0 4552 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3596
timestamp 1680363874
transform 1 0 4552 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1680363874
transform 1 0 4560 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3597
timestamp 1680363874
transform 1 0 4656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1680363874
transform 1 0 4664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1680363874
transform 1 0 4672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1680363874
transform 1 0 4680 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_242
timestamp 1680363874
transform -1 0 4784 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3605
timestamp 1680363874
transform 1 0 4784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1680363874
transform 1 0 4792 0 -1 3170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_33
timestamp 1680363874
transform 1 0 4851 0 1 3070
box -10 -3 10 3
use M3_M2  M3_M2_3248
timestamp 1680363874
transform 1 0 68 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1680363874
transform 1 0 84 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1680363874
transform 1 0 108 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3635
timestamp 1680363874
transform 1 0 148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1680363874
transform 1 0 220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1680363874
transform 1 0 268 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3326
timestamp 1680363874
transform 1 0 268 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3784
timestamp 1680363874
transform 1 0 284 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1680363874
transform 1 0 316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1680363874
transform 1 0 324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1680363874
transform 1 0 332 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3368
timestamp 1680363874
transform 1 0 332 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1680363874
transform 1 0 444 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1680363874
transform 1 0 348 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3638
timestamp 1680363874
transform 1 0 348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1680363874
transform 1 0 364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1680363874
transform 1 0 372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1680363874
transform 1 0 356 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3327
timestamp 1680363874
transform 1 0 364 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1680363874
transform 1 0 436 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1680363874
transform 1 0 460 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3369
timestamp 1680363874
transform 1 0 356 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1680363874
transform 1 0 452 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3621
timestamp 1680363874
transform 1 0 492 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1680363874
transform 1 0 508 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3329
timestamp 1680363874
transform 1 0 508 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1680363874
transform 1 0 500 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3622
timestamp 1680363874
transform 1 0 524 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1680363874
transform 1 0 524 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3265
timestamp 1680363874
transform 1 0 540 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3641
timestamp 1680363874
transform 1 0 540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1680363874
transform 1 0 564 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3330
timestamp 1680363874
transform 1 0 572 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3729
timestamp 1680363874
transform 1 0 612 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3240
timestamp 1680363874
transform 1 0 644 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3623
timestamp 1680363874
transform 1 0 636 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3331
timestamp 1680363874
transform 1 0 636 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3624
timestamp 1680363874
transform 1 0 644 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3266
timestamp 1680363874
transform 1 0 652 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1680363874
transform 1 0 660 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3642
timestamp 1680363874
transform 1 0 700 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3289
timestamp 1680363874
transform 1 0 748 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3643
timestamp 1680363874
transform 1 0 756 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1680363874
transform 1 0 764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1680363874
transform 1 0 676 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3290
timestamp 1680363874
transform 1 0 772 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1680363874
transform 1 0 852 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3645
timestamp 1680363874
transform 1 0 852 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1680363874
transform 1 0 868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1680363874
transform 1 0 868 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3333
timestamp 1680363874
transform 1 0 868 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1680363874
transform 1 0 892 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3647
timestamp 1680363874
transform 1 0 892 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1680363874
transform 1 0 908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3269
timestamp 1680363874
transform 1 0 972 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3733
timestamp 1680363874
transform 1 0 964 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1680363874
transform 1 0 972 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3334
timestamp 1680363874
transform 1 0 964 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1680363874
transform 1 0 1004 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1680363874
transform 1 0 1036 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3648
timestamp 1680363874
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3335
timestamp 1680363874
transform 1 0 1020 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1680363874
transform 1 0 1012 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3649
timestamp 1680363874
transform 1 0 1076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1680363874
transform 1 0 1084 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3241
timestamp 1680363874
transform 1 0 1124 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3625
timestamp 1680363874
transform 1 0 1124 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1680363874
transform 1 0 1116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1680363874
transform 1 0 1124 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3336
timestamp 1680363874
transform 1 0 1124 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1680363874
transform 1 0 1108 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1680363874
transform 1 0 1164 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3736
timestamp 1680363874
transform 1 0 1164 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1680363874
transform 1 0 1172 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3337
timestamp 1680363874
transform 1 0 1172 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1680363874
transform 1 0 1212 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1680363874
transform 1 0 1204 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3652
timestamp 1680363874
transform 1 0 1212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1680363874
transform 1 0 1204 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3228
timestamp 1680363874
transform 1 0 1244 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3653
timestamp 1680363874
transform 1 0 1236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1680363874
transform 1 0 1268 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1680363874
transform 1 0 1260 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3272
timestamp 1680363874
transform 1 0 1268 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1680363874
transform 1 0 1260 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1680363874
transform 1 0 1268 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3627
timestamp 1680363874
transform 1 0 1292 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3242
timestamp 1680363874
transform 1 0 1324 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3617
timestamp 1680363874
transform 1 0 1324 0 1 3035
box -2 -2 2 2
use M3_M2  M3_M2_3250
timestamp 1680363874
transform 1 0 1340 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1680363874
transform 1 0 1356 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1680363874
transform 1 0 1332 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3654
timestamp 1680363874
transform 1 0 1332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1680363874
transform 1 0 1348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1680363874
transform 1 0 1324 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3339
timestamp 1680363874
transform 1 0 1316 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1680363874
transform 1 0 1348 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1680363874
transform 1 0 1340 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1680363874
transform 1 0 1372 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1680363874
transform 1 0 1364 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1680363874
transform 1 0 1396 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3628
timestamp 1680363874
transform 1 0 1388 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3292
timestamp 1680363874
transform 1 0 1380 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1680363874
transform 1 0 1412 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3618
timestamp 1680363874
transform 1 0 1428 0 1 3035
box -2 -2 2 2
use M3_M2  M3_M2_3274
timestamp 1680363874
transform 1 0 1420 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1680363874
transform 1 0 1444 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3629
timestamp 1680363874
transform 1 0 1436 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1680363874
transform 1 0 1404 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3293
timestamp 1680363874
transform 1 0 1412 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3657
timestamp 1680363874
transform 1 0 1420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1680363874
transform 1 0 1404 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3315
timestamp 1680363874
transform 1 0 1412 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3658
timestamp 1680363874
transform 1 0 1444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1680363874
transform 1 0 1444 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3375
timestamp 1680363874
transform 1 0 1444 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1680363874
transform 1 0 1508 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3659
timestamp 1680363874
transform 1 0 1492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1680363874
transform 1 0 1508 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3294
timestamp 1680363874
transform 1 0 1516 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3661
timestamp 1680363874
transform 1 0 1524 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3341
timestamp 1680363874
transform 1 0 1508 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1680363874
transform 1 0 1516 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1680363874
transform 1 0 1540 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3742
timestamp 1680363874
transform 1 0 1556 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3377
timestamp 1680363874
transform 1 0 1548 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1680363874
transform 1 0 1572 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3662
timestamp 1680363874
transform 1 0 1620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1680363874
transform 1 0 1572 0 1 3007
box -2 -2 2 2
use M3_M2  M3_M2_3378
timestamp 1680363874
transform 1 0 1620 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3663
timestamp 1680363874
transform 1 0 1668 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3316
timestamp 1680363874
transform 1 0 1668 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1680363874
transform 1 0 1668 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1680363874
transform 1 0 1684 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1680363874
transform 1 0 1700 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3664
timestamp 1680363874
transform 1 0 1748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1680363874
transform 1 0 1780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1680363874
transform 1 0 1820 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1680363874
transform 1 0 1700 0 1 3007
box -2 -2 2 2
use M3_M2  M3_M2_3343
timestamp 1680363874
transform 1 0 1724 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1680363874
transform 1 0 1692 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3743
timestamp 1680363874
transform 1 0 1796 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3344
timestamp 1680363874
transform 1 0 1796 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3667
timestamp 1680363874
transform 1 0 1900 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3244
timestamp 1680363874
transform 1 0 1980 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3668
timestamp 1680363874
transform 1 0 1972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1680363874
transform 1 0 1932 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3345
timestamp 1680363874
transform 1 0 1932 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3669
timestamp 1680363874
transform 1 0 2036 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3380
timestamp 1680363874
transform 1 0 2060 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3670
timestamp 1680363874
transform 1 0 2108 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3298
timestamp 1680363874
transform 1 0 2124 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1680363874
transform 1 0 2164 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3671
timestamp 1680363874
transform 1 0 2172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1680363874
transform 1 0 2084 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3346
timestamp 1680363874
transform 1 0 2084 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1680363874
transform 1 0 2100 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1680363874
transform 1 0 2212 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1680363874
transform 1 0 2268 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1680363874
transform 1 0 2228 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3619
timestamp 1680363874
transform 1 0 2316 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1680363874
transform 1 0 2252 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1680363874
transform 1 0 2308 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1680363874
transform 1 0 2228 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3318
timestamp 1680363874
transform 1 0 2252 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1680363874
transform 1 0 2228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1680363874
transform 1 0 2292 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3620
timestamp 1680363874
transform 1 0 2348 0 1 3035
box -2 -2 2 2
use M3_M2  M3_M2_3276
timestamp 1680363874
transform 1 0 2356 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3674
timestamp 1680363874
transform 1 0 2356 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3231
timestamp 1680363874
transform 1 0 2364 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3675
timestamp 1680363874
transform 1 0 2364 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3319
timestamp 1680363874
transform 1 0 2364 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3747
timestamp 1680363874
transform 1 0 2372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3232
timestamp 1680363874
transform 1 0 2388 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3676
timestamp 1680363874
transform 1 0 2404 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1680363874
transform 1 0 2444 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3253
timestamp 1680363874
transform 1 0 2468 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3677
timestamp 1680363874
transform 1 0 2468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1680363874
transform 1 0 2492 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3320
timestamp 1680363874
transform 1 0 2508 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1680363874
transform 1 0 2524 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1680363874
transform 1 0 2556 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1680363874
transform 1 0 2524 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3678
timestamp 1680363874
transform 1 0 2556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1680363874
transform 1 0 2524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1680363874
transform 1 0 2628 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3254
timestamp 1680363874
transform 1 0 2764 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1680363874
transform 1 0 2700 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3680
timestamp 1680363874
transform 1 0 2724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1680363874
transform 1 0 2700 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3349
timestamp 1680363874
transform 1 0 2700 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1680363874
transform 1 0 2724 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3681
timestamp 1680363874
transform 1 0 2788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1680363874
transform 1 0 2796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1680363874
transform 1 0 2812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1680363874
transform 1 0 2820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1680363874
transform 1 0 2868 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3351
timestamp 1680363874
transform 1 0 2876 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1680363874
transform 1 0 2892 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1680363874
transform 1 0 2908 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3753
timestamp 1680363874
transform 1 0 2900 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3256
timestamp 1680363874
transform 1 0 2932 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3630
timestamp 1680363874
transform 1 0 2932 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3234
timestamp 1680363874
transform 1 0 2948 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1680363874
transform 1 0 2964 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1680363874
transform 1 0 2972 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3631
timestamp 1680363874
transform 1 0 2972 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1680363874
transform 1 0 2948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1680363874
transform 1 0 2956 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3280
timestamp 1680363874
transform 1 0 2996 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1680363874
transform 1 0 3044 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3754
timestamp 1680363874
transform 1 0 3044 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3352
timestamp 1680363874
transform 1 0 3036 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1680363874
transform 1 0 3060 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3687
timestamp 1680363874
transform 1 0 3092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1680363874
transform 1 0 3060 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3353
timestamp 1680363874
transform 1 0 3060 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3688
timestamp 1680363874
transform 1 0 3180 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3301
timestamp 1680363874
transform 1 0 3212 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1680363874
transform 1 0 3260 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3632
timestamp 1680363874
transform 1 0 3260 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1680363874
transform 1 0 3244 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3354
timestamp 1680363874
transform 1 0 3244 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3690
timestamp 1680363874
transform 1 0 3284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1680363874
transform 1 0 3300 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3383
timestamp 1680363874
transform 1 0 3300 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3691
timestamp 1680363874
transform 1 0 3316 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3321
timestamp 1680363874
transform 1 0 3316 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1680363874
transform 1 0 3332 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3692
timestamp 1680363874
transform 1 0 3340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1680363874
transform 1 0 3332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1680363874
transform 1 0 3372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3355
timestamp 1680363874
transform 1 0 3364 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3693
timestamp 1680363874
transform 1 0 3460 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3302
timestamp 1680363874
transform 1 0 3492 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3759
timestamp 1680363874
transform 1 0 3428 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3322
timestamp 1680363874
transform 1 0 3468 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1680363874
transform 1 0 3428 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1680363874
transform 1 0 3476 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3694
timestamp 1680363874
transform 1 0 3516 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3235
timestamp 1680363874
transform 1 0 3532 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1680363874
transform 1 0 3548 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3695
timestamp 1680363874
transform 1 0 3548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1680363874
transform 1 0 3572 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1680363874
transform 1 0 3580 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3283
timestamp 1680363874
transform 1 0 3596 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3760
timestamp 1680363874
transform 1 0 3596 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3358
timestamp 1680363874
transform 1 0 3604 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1680363874
transform 1 0 3620 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1680363874
transform 1 0 3620 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3761
timestamp 1680363874
transform 1 0 3620 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1680363874
transform 1 0 3628 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3359
timestamp 1680363874
transform 1 0 3628 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3697
timestamp 1680363874
transform 1 0 3684 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1680363874
transform 1 0 3700 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3304
timestamp 1680363874
transform 1 0 3708 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1680363874
transform 1 0 3724 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3699
timestamp 1680363874
transform 1 0 3716 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1680363874
transform 1 0 3724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1680363874
transform 1 0 3692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1680363874
transform 1 0 3708 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3360
timestamp 1680363874
transform 1 0 3692 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1680363874
transform 1 0 3724 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1680363874
transform 1 0 3764 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3701
timestamp 1680363874
transform 1 0 3812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1680363874
transform 1 0 3844 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3323
timestamp 1680363874
transform 1 0 3868 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3766
timestamp 1680363874
transform 1 0 3876 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3247
timestamp 1680363874
transform 1 0 3932 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3702
timestamp 1680363874
transform 1 0 3940 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3384
timestamp 1680363874
transform 1 0 4060 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3767
timestamp 1680363874
transform 1 0 4076 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3238
timestamp 1680363874
transform 1 0 4108 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3703
timestamp 1680363874
transform 1 0 4116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1680363874
transform 1 0 4092 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3385
timestamp 1680363874
transform 1 0 4084 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1680363874
transform 1 0 4188 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3704
timestamp 1680363874
transform 1 0 4180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1680363874
transform 1 0 4188 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3227
timestamp 1680363874
transform 1 0 4204 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3769
timestamp 1680363874
transform 1 0 4212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1680363874
transform 1 0 4244 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3305
timestamp 1680363874
transform 1 0 4260 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3786
timestamp 1680363874
transform 1 0 4260 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3386
timestamp 1680363874
transform 1 0 4276 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3707
timestamp 1680363874
transform 1 0 4292 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3306
timestamp 1680363874
transform 1 0 4308 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3770
timestamp 1680363874
transform 1 0 4300 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1680363874
transform 1 0 4308 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3362
timestamp 1680363874
transform 1 0 4292 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1680363874
transform 1 0 4324 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3787
timestamp 1680363874
transform 1 0 4316 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3363
timestamp 1680363874
transform 1 0 4324 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1680363874
transform 1 0 4316 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3788
timestamp 1680363874
transform 1 0 4340 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3308
timestamp 1680363874
transform 1 0 4372 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3708
timestamp 1680363874
transform 1 0 4396 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3309
timestamp 1680363874
transform 1 0 4404 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1680363874
transform 1 0 4420 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3709
timestamp 1680363874
transform 1 0 4420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1680363874
transform 1 0 4380 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1680363874
transform 1 0 4388 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1680363874
transform 1 0 4404 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1680363874
transform 1 0 4412 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3364
timestamp 1680363874
transform 1 0 4380 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1680363874
transform 1 0 4388 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1680363874
transform 1 0 4436 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1680363874
transform 1 0 4452 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3710
timestamp 1680363874
transform 1 0 4508 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1680363874
transform 1 0 4556 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3324
timestamp 1680363874
transform 1 0 4548 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1680363874
transform 1 0 4580 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3712
timestamp 1680363874
transform 1 0 4588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1680363874
transform 1 0 4564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1680363874
transform 1 0 4580 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3366
timestamp 1680363874
transform 1 0 4564 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3778
timestamp 1680363874
transform 1 0 4604 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1680363874
transform 1 0 4612 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3389
timestamp 1680363874
transform 1 0 4612 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1680363874
transform 1 0 4660 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3713
timestamp 1680363874
transform 1 0 4628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1680363874
transform 1 0 4644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1680363874
transform 1 0 4660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1680363874
transform 1 0 4652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1680363874
transform 1 0 4660 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3367
timestamp 1680363874
transform 1 0 4652 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1680363874
transform 1 0 4660 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3716
timestamp 1680363874
transform 1 0 4684 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3311
timestamp 1680363874
transform 1 0 4692 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1680363874
transform 1 0 4732 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3717
timestamp 1680363874
transform 1 0 4700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1680363874
transform 1 0 4716 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3312
timestamp 1680363874
transform 1 0 4724 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3782
timestamp 1680363874
transform 1 0 4724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1680363874
transform 1 0 4732 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3288
timestamp 1680363874
transform 1 0 4756 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3719
timestamp 1680363874
transform 1 0 4756 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3262
timestamp 1680363874
transform 1 0 4764 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3634
timestamp 1680363874
transform 1 0 4764 0 1 3025
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_34
timestamp 1680363874
transform 1 0 48 0 1 2970
box -10 -3 10 3
use FILL  FILL_3607
timestamp 1680363874
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1680363874
transform 1 0 80 0 1 2970
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1680363874
transform 1 0 88 0 1 2970
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1680363874
transform 1 0 96 0 1 2970
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1680363874
transform 1 0 104 0 1 2970
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1680363874
transform 1 0 112 0 1 2970
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1680363874
transform 1 0 120 0 1 2970
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1680363874
transform 1 0 128 0 1 2970
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1680363874
transform 1 0 136 0 1 2970
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1680363874
transform 1 0 144 0 1 2970
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1680363874
transform 1 0 152 0 1 2970
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1680363874
transform 1 0 160 0 1 2970
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1680363874
transform 1 0 168 0 1 2970
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1680363874
transform 1 0 176 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1680363874
transform -1 0 280 0 1 2970
box -8 -3 104 105
use FILL  FILL_3621
timestamp 1680363874
transform 1 0 280 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_35
timestamp 1680363874
transform 1 0 288 0 1 2970
box -8 -3 32 105
use FILL  FILL_3628
timestamp 1680363874
transform 1 0 312 0 1 2970
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1680363874
transform 1 0 320 0 1 2970
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1680363874
transform 1 0 328 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_260
timestamp 1680363874
transform 1 0 336 0 1 2970
box -9 -3 26 105
use FAX1  FAX1_0
timestamp 1680363874
transform 1 0 352 0 1 2970
box -5 -3 126 105
use FILL  FILL_3635
timestamp 1680363874
transform 1 0 472 0 1 2970
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1680363874
transform 1 0 480 0 1 2970
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1680363874
transform 1 0 488 0 1 2970
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1680363874
transform 1 0 496 0 1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1680363874
transform -1 0 528 0 1 2970
box -8 -3 32 105
use FILL  FILL_3639
timestamp 1680363874
transform 1 0 528 0 1 2970
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1680363874
transform 1 0 536 0 1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1680363874
transform -1 0 568 0 1 2970
box -8 -3 32 105
use FILL  FILL_3641
timestamp 1680363874
transform 1 0 568 0 1 2970
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1680363874
transform 1 0 576 0 1 2970
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1680363874
transform 1 0 584 0 1 2970
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1680363874
transform 1 0 592 0 1 2970
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1680363874
transform 1 0 600 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_105
timestamp 1680363874
transform 1 0 608 0 1 2970
box -8 -3 34 105
use FILL  FILL_3661
timestamp 1680363874
transform 1 0 640 0 1 2970
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1680363874
transform 1 0 648 0 1 2970
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1680363874
transform 1 0 656 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1680363874
transform 1 0 664 0 1 2970
box -8 -3 104 105
use FILL  FILL_3664
timestamp 1680363874
transform 1 0 760 0 1 2970
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1680363874
transform 1 0 768 0 1 2970
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1680363874
transform 1 0 776 0 1 2970
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1680363874
transform 1 0 784 0 1 2970
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1680363874
transform 1 0 792 0 1 2970
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1680363874
transform 1 0 800 0 1 2970
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1680363874
transform 1 0 808 0 1 2970
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1680363874
transform 1 0 816 0 1 2970
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1680363874
transform 1 0 824 0 1 2970
box -8 -3 16 105
use AND2X2  AND2X2_9
timestamp 1680363874
transform -1 0 864 0 1 2970
box -8 -3 40 105
use FILL  FILL_3677
timestamp 1680363874
transform 1 0 864 0 1 2970
box -8 -3 16 105
use AND2X2  AND2X2_10
timestamp 1680363874
transform -1 0 904 0 1 2970
box -8 -3 40 105
use FILL  FILL_3678
timestamp 1680363874
transform 1 0 904 0 1 2970
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1680363874
transform 1 0 912 0 1 2970
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1680363874
transform 1 0 920 0 1 2970
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1680363874
transform 1 0 928 0 1 2970
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1680363874
transform 1 0 936 0 1 2970
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1680363874
transform 1 0 944 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_261
timestamp 1680363874
transform -1 0 968 0 1 2970
box -9 -3 26 105
use FILL  FILL_3695
timestamp 1680363874
transform 1 0 968 0 1 2970
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1680363874
transform 1 0 976 0 1 2970
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1680363874
transform 1 0 984 0 1 2970
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1680363874
transform 1 0 992 0 1 2970
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1680363874
transform 1 0 1000 0 1 2970
box -8 -3 16 105
use AND2X2  AND2X2_12
timestamp 1680363874
transform 1 0 1008 0 1 2970
box -8 -3 40 105
use FILL  FILL_3700
timestamp 1680363874
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1680363874
transform 1 0 1048 0 1 2970
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1680363874
transform 1 0 1056 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_263
timestamp 1680363874
transform 1 0 1064 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1680363874
transform -1 0 1096 0 1 2970
box -9 -3 26 105
use AND2X2  AND2X2_13
timestamp 1680363874
transform -1 0 1128 0 1 2970
box -8 -3 40 105
use FILL  FILL_3711
timestamp 1680363874
transform 1 0 1128 0 1 2970
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1680363874
transform 1 0 1136 0 1 2970
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1680363874
transform 1 0 1144 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_265
timestamp 1680363874
transform -1 0 1168 0 1 2970
box -9 -3 26 105
use FILL  FILL_3720
timestamp 1680363874
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1680363874
transform 1 0 1176 0 1 2970
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1680363874
transform 1 0 1184 0 1 2970
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1680363874
transform 1 0 1192 0 1 2970
box -8 -3 16 105
use AND2X2  AND2X2_15
timestamp 1680363874
transform 1 0 1200 0 1 2970
box -8 -3 40 105
use FILL  FILL_3724
timestamp 1680363874
transform 1 0 1232 0 1 2970
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1680363874
transform 1 0 1240 0 1 2970
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1680363874
transform 1 0 1248 0 1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_3
timestamp 1680363874
transform -1 0 1288 0 1 2970
box -8 -3 40 105
use FILL  FILL_3736
timestamp 1680363874
transform 1 0 1288 0 1 2970
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1680363874
transform 1 0 1296 0 1 2970
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1680363874
transform 1 0 1304 0 1 2970
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1680363874
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1680363874
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_134
timestamp 1680363874
transform 1 0 1328 0 1 2970
box -8 -3 46 105
use FILL  FILL_3747
timestamp 1680363874
transform 1 0 1368 0 1 2970
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1680363874
transform 1 0 1376 0 1 2970
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1680363874
transform 1 0 1384 0 1 2970
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1680363874
transform 1 0 1392 0 1 2970
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1680363874
transform 1 0 1400 0 1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1680363874
transform 1 0 1408 0 1 2970
box -8 -3 40 105
use FILL  FILL_3762
timestamp 1680363874
transform 1 0 1440 0 1 2970
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1680363874
transform 1 0 1448 0 1 2970
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1680363874
transform 1 0 1456 0 1 2970
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1680363874
transform 1 0 1464 0 1 2970
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1680363874
transform 1 0 1472 0 1 2970
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1680363874
transform 1 0 1480 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_135
timestamp 1680363874
transform 1 0 1488 0 1 2970
box -8 -3 46 105
use FILL  FILL_3776
timestamp 1680363874
transform 1 0 1528 0 1 2970
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1680363874
transform 1 0 1536 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3391
timestamp 1680363874
transform 1 0 1556 0 1 2975
box -3 -3 3 3
use FILL  FILL_3780
timestamp 1680363874
transform 1 0 1544 0 1 2970
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1680363874
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3392
timestamp 1680363874
transform 1 0 1580 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_248
timestamp 1680363874
transform 1 0 1560 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_267
timestamp 1680363874
transform 1 0 1656 0 1 2970
box -9 -3 26 105
use FILL  FILL_3783
timestamp 1680363874
transform 1 0 1672 0 1 2970
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1680363874
transform 1 0 1680 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_249
timestamp 1680363874
transform 1 0 1688 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1680363874
transform 1 0 1784 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_268
timestamp 1680363874
transform 1 0 1880 0 1 2970
box -9 -3 26 105
use FILL  FILL_3785
timestamp 1680363874
transform 1 0 1896 0 1 2970
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1680363874
transform 1 0 1904 0 1 2970
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1680363874
transform 1 0 1912 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1680363874
transform 1 0 1920 0 1 2970
box -8 -3 104 105
use FILL  FILL_3788
timestamp 1680363874
transform 1 0 2016 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_269
timestamp 1680363874
transform 1 0 2024 0 1 2970
box -9 -3 26 105
use FILL  FILL_3789
timestamp 1680363874
transform 1 0 2040 0 1 2970
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1680363874
transform 1 0 2048 0 1 2970
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1680363874
transform 1 0 2056 0 1 2970
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1680363874
transform 1 0 2064 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1680363874
transform 1 0 2072 0 1 2970
box -8 -3 104 105
use FILL  FILL_3813
timestamp 1680363874
transform 1 0 2168 0 1 2970
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1680363874
transform 1 0 2176 0 1 2970
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1680363874
transform 1 0 2184 0 1 2970
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1680363874
transform 1 0 2192 0 1 2970
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1680363874
transform 1 0 2200 0 1 2970
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1680363874
transform 1 0 2208 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1680363874
transform 1 0 2216 0 1 2970
box -8 -3 104 105
use FILL  FILL_3825
timestamp 1680363874
transform 1 0 2312 0 1 2970
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1680363874
transform 1 0 2320 0 1 2970
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1680363874
transform 1 0 2328 0 1 2970
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1680363874
transform 1 0 2336 0 1 2970
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1680363874
transform 1 0 2344 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_274
timestamp 1680363874
transform 1 0 2352 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1680363874
transform 1 0 2368 0 1 2970
box -9 -3 26 105
use FILL  FILL_3836
timestamp 1680363874
transform 1 0 2384 0 1 2970
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1680363874
transform 1 0 2392 0 1 2970
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1680363874
transform 1 0 2400 0 1 2970
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1680363874
transform 1 0 2408 0 1 2970
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1680363874
transform 1 0 2416 0 1 2970
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1680363874
transform 1 0 2424 0 1 2970
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1680363874
transform 1 0 2432 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3393
timestamp 1680363874
transform 1 0 2452 0 1 2975
box -3 -3 3 3
use FILL  FILL_3843
timestamp 1680363874
transform 1 0 2440 0 1 2970
box -8 -3 16 105
use AND2X2  AND2X2_16
timestamp 1680363874
transform -1 0 2480 0 1 2970
box -8 -3 40 105
use FILL  FILL_3844
timestamp 1680363874
transform 1 0 2480 0 1 2970
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1680363874
transform 1 0 2488 0 1 2970
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1680363874
transform 1 0 2496 0 1 2970
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1680363874
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1680363874
transform 1 0 2512 0 1 2970
box -8 -3 104 105
use FILL  FILL_3856
timestamp 1680363874
transform 1 0 2608 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_276
timestamp 1680363874
transform 1 0 2616 0 1 2970
box -9 -3 26 105
use FILL  FILL_3857
timestamp 1680363874
transform 1 0 2632 0 1 2970
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1680363874
transform 1 0 2640 0 1 2970
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1680363874
transform 1 0 2648 0 1 2970
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1680363874
transform 1 0 2656 0 1 2970
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1680363874
transform 1 0 2664 0 1 2970
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1680363874
transform 1 0 2672 0 1 2970
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1680363874
transform 1 0 2680 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1680363874
transform 1 0 2688 0 1 2970
box -8 -3 104 105
use FILL  FILL_3875
timestamp 1680363874
transform 1 0 2784 0 1 2970
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1680363874
transform 1 0 2792 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3394
timestamp 1680363874
transform 1 0 2820 0 1 2975
box -3 -3 3 3
use INVX2  INVX2_277
timestamp 1680363874
transform -1 0 2816 0 1 2970
box -9 -3 26 105
use FILL  FILL_3883
timestamp 1680363874
transform 1 0 2816 0 1 2970
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1680363874
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1680363874
transform 1 0 2832 0 1 2970
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1680363874
transform 1 0 2840 0 1 2970
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1680363874
transform 1 0 2848 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_106
timestamp 1680363874
transform 1 0 2856 0 1 2970
box -8 -3 34 105
use FILL  FILL_3894
timestamp 1680363874
transform 1 0 2888 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3395
timestamp 1680363874
transform 1 0 2908 0 1 2975
box -3 -3 3 3
use FILL  FILL_3895
timestamp 1680363874
transform 1 0 2896 0 1 2970
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1680363874
transform 1 0 2904 0 1 2970
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1680363874
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1680363874
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1680363874
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1680363874
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_108
timestamp 1680363874
transform 1 0 2944 0 1 2970
box -8 -3 34 105
use FILL  FILL_3905
timestamp 1680363874
transform 1 0 2976 0 1 2970
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1680363874
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1680363874
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1680363874
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1680363874
transform 1 0 3008 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3396
timestamp 1680363874
transform 1 0 3028 0 1 2975
box -3 -3 3 3
use FILL  FILL_3917
timestamp 1680363874
transform 1 0 3016 0 1 2970
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1680363874
transform 1 0 3024 0 1 2970
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1680363874
transform 1 0 3032 0 1 2970
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1680363874
transform 1 0 3040 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3397
timestamp 1680363874
transform 1 0 3148 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_259
timestamp 1680363874
transform 1 0 3048 0 1 2970
box -8 -3 104 105
use FILL  FILL_3923
timestamp 1680363874
transform 1 0 3144 0 1 2970
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1680363874
transform 1 0 3152 0 1 2970
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1680363874
transform 1 0 3160 0 1 2970
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1680363874
transform 1 0 3168 0 1 2970
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1680363874
transform 1 0 3176 0 1 2970
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1680363874
transform 1 0 3184 0 1 2970
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1680363874
transform 1 0 3192 0 1 2970
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1680363874
transform 1 0 3200 0 1 2970
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1680363874
transform 1 0 3208 0 1 2970
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1680363874
transform 1 0 3216 0 1 2970
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1680363874
transform 1 0 3224 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_110
timestamp 1680363874
transform 1 0 3232 0 1 2970
box -8 -3 34 105
use FILL  FILL_3955
timestamp 1680363874
transform 1 0 3264 0 1 2970
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1680363874
transform 1 0 3272 0 1 2970
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1680363874
transform 1 0 3280 0 1 2970
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1680363874
transform 1 0 3288 0 1 2970
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1680363874
transform 1 0 3296 0 1 2970
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1680363874
transform 1 0 3304 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3398
timestamp 1680363874
transform 1 0 3332 0 1 2975
box -3 -3 3 3
use BUFX2  BUFX2_24
timestamp 1680363874
transform 1 0 3312 0 1 2970
box -5 -3 28 105
use FILL  FILL_3961
timestamp 1680363874
transform 1 0 3336 0 1 2970
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1680363874
transform 1 0 3344 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_25
timestamp 1680363874
transform 1 0 3352 0 1 2970
box -5 -3 28 105
use FILL  FILL_3973
timestamp 1680363874
transform 1 0 3376 0 1 2970
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1680363874
transform 1 0 3384 0 1 2970
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1680363874
transform 1 0 3392 0 1 2970
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1680363874
transform 1 0 3400 0 1 2970
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1680363874
transform 1 0 3408 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1680363874
transform 1 0 3416 0 1 2970
box -8 -3 104 105
use FILL  FILL_3984
timestamp 1680363874
transform 1 0 3512 0 1 2970
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1680363874
transform 1 0 3520 0 1 2970
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1680363874
transform 1 0 3528 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_111
timestamp 1680363874
transform 1 0 3536 0 1 2970
box -8 -3 34 105
use FILL  FILL_3987
timestamp 1680363874
transform 1 0 3568 0 1 2970
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1680363874
transform 1 0 3576 0 1 2970
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1680363874
transform 1 0 3584 0 1 2970
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1680363874
transform 1 0 3592 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_281
timestamp 1680363874
transform -1 0 3616 0 1 2970
box -9 -3 26 105
use FILL  FILL_3991
timestamp 1680363874
transform 1 0 3616 0 1 2970
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1680363874
transform 1 0 3624 0 1 2970
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1680363874
transform 1 0 3632 0 1 2970
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1680363874
transform 1 0 3640 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3399
timestamp 1680363874
transform 1 0 3660 0 1 2975
box -3 -3 3 3
use FILL  FILL_4004
timestamp 1680363874
transform 1 0 3648 0 1 2970
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1680363874
transform 1 0 3656 0 1 2970
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1680363874
transform 1 0 3664 0 1 2970
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1680363874
transform 1 0 3672 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_138
timestamp 1680363874
transform -1 0 3720 0 1 2970
box -8 -3 46 105
use FILL  FILL_4008
timestamp 1680363874
transform 1 0 3720 0 1 2970
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1680363874
transform 1 0 3728 0 1 2970
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1680363874
transform 1 0 3736 0 1 2970
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1680363874
transform 1 0 3744 0 1 2970
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1680363874
transform 1 0 3752 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1680363874
transform -1 0 3856 0 1 2970
box -8 -3 104 105
use FILL  FILL_4020
timestamp 1680363874
transform 1 0 3856 0 1 2970
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1680363874
transform 1 0 3864 0 1 2970
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1680363874
transform 1 0 3872 0 1 2970
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1680363874
transform 1 0 3880 0 1 2970
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1680363874
transform 1 0 3888 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_28
timestamp 1680363874
transform -1 0 3920 0 1 2970
box -5 -3 28 105
use FILL  FILL_4025
timestamp 1680363874
transform 1 0 3920 0 1 2970
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1680363874
transform 1 0 3928 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_29
timestamp 1680363874
transform 1 0 3936 0 1 2970
box -5 -3 28 105
use FILL  FILL_4027
timestamp 1680363874
transform 1 0 3960 0 1 2970
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1680363874
transform 1 0 3968 0 1 2970
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1680363874
transform 1 0 3976 0 1 2970
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1680363874
transform 1 0 3984 0 1 2970
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1680363874
transform 1 0 3992 0 1 2970
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1680363874
transform 1 0 4000 0 1 2970
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1680363874
transform 1 0 4008 0 1 2970
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1680363874
transform 1 0 4016 0 1 2970
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1680363874
transform 1 0 4024 0 1 2970
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1680363874
transform 1 0 4032 0 1 2970
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1680363874
transform 1 0 4040 0 1 2970
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1680363874
transform 1 0 4048 0 1 2970
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1680363874
transform 1 0 4056 0 1 2970
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1680363874
transform 1 0 4064 0 1 2970
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1680363874
transform 1 0 4072 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1680363874
transform 1 0 4080 0 1 2970
box -8 -3 104 105
use FILL  FILL_4048
timestamp 1680363874
transform 1 0 4176 0 1 2970
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1680363874
transform 1 0 4184 0 1 2970
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1680363874
transform 1 0 4192 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_36
timestamp 1680363874
transform -1 0 4224 0 1 2970
box -8 -3 32 105
use FILL  FILL_4063
timestamp 1680363874
transform 1 0 4224 0 1 2970
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1680363874
transform 1 0 4232 0 1 2970
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1680363874
transform 1 0 4240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1680363874
transform 1 0 4248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1680363874
transform 1 0 4256 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_38
timestamp 1680363874
transform -1 0 4288 0 1 2970
box -8 -3 32 105
use FILL  FILL_4072
timestamp 1680363874
transform 1 0 4288 0 1 2970
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1680363874
transform 1 0 4296 0 1 2970
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1680363874
transform 1 0 4304 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_39
timestamp 1680363874
transform -1 0 4336 0 1 2970
box -8 -3 32 105
use FILL  FILL_4077
timestamp 1680363874
transform 1 0 4336 0 1 2970
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1680363874
transform 1 0 4344 0 1 2970
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1680363874
transform 1 0 4352 0 1 2970
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1680363874
transform 1 0 4360 0 1 2970
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1680363874
transform 1 0 4368 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_141
timestamp 1680363874
transform 1 0 4376 0 1 2970
box -8 -3 46 105
use FILL  FILL_4090
timestamp 1680363874
transform 1 0 4416 0 1 2970
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1680363874
transform 1 0 4424 0 1 2970
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1680363874
transform 1 0 4432 0 1 2970
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1680363874
transform 1 0 4440 0 1 2970
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1680363874
transform 1 0 4448 0 1 2970
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1680363874
transform 1 0 4456 0 1 2970
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1680363874
transform 1 0 4464 0 1 2970
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1680363874
transform 1 0 4472 0 1 2970
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1680363874
transform 1 0 4480 0 1 2970
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1680363874
transform 1 0 4488 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_284
timestamp 1680363874
transform 1 0 4496 0 1 2970
box -9 -3 26 105
use FILL  FILL_4104
timestamp 1680363874
transform 1 0 4512 0 1 2970
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1680363874
transform 1 0 4520 0 1 2970
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1680363874
transform 1 0 4528 0 1 2970
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1680363874
transform 1 0 4536 0 1 2970
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1680363874
transform 1 0 4544 0 1 2970
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1680363874
transform 1 0 4552 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_216
timestamp 1680363874
transform 1 0 4560 0 1 2970
box -8 -3 46 105
use FILL  FILL_4113
timestamp 1680363874
transform 1 0 4600 0 1 2970
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1680363874
transform 1 0 4608 0 1 2970
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1680363874
transform 1 0 4616 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_142
timestamp 1680363874
transform 1 0 4624 0 1 2970
box -8 -3 46 105
use FILL  FILL_4124
timestamp 1680363874
transform 1 0 4664 0 1 2970
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1680363874
transform 1 0 4672 0 1 2970
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1680363874
transform 1 0 4680 0 1 2970
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1680363874
transform 1 0 4688 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_144
timestamp 1680363874
transform 1 0 4696 0 1 2970
box -8 -3 46 105
use FILL  FILL_4131
timestamp 1680363874
transform 1 0 4736 0 1 2970
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1680363874
transform 1 0 4744 0 1 2970
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1680363874
transform 1 0 4752 0 1 2970
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1680363874
transform 1 0 4760 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_285
timestamp 1680363874
transform 1 0 4768 0 1 2970
box -9 -3 26 105
use FILL  FILL_4135
timestamp 1680363874
transform 1 0 4784 0 1 2970
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1680363874
transform 1 0 4792 0 1 2970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_35
timestamp 1680363874
transform 1 0 4827 0 1 2970
box -10 -3 10 3
use M3_M2  M3_M2_3418
timestamp 1680363874
transform 1 0 116 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3797
timestamp 1680363874
transform 1 0 84 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3461
timestamp 1680363874
transform 1 0 148 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1680363874
transform 1 0 180 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3798
timestamp 1680363874
transform 1 0 172 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3462
timestamp 1680363874
transform 1 0 188 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3877
timestamp 1680363874
transform 1 0 124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1680363874
transform 1 0 164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1680363874
transform 1 0 180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1680363874
transform 1 0 188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1680363874
transform 1 0 204 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3548
timestamp 1680363874
transform 1 0 100 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1680363874
transform 1 0 116 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1680363874
transform 1 0 180 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3971
timestamp 1680363874
transform 1 0 188 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1680363874
transform 1 0 220 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3412
timestamp 1680363874
transform 1 0 244 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3792
timestamp 1680363874
transform 1 0 244 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3420
timestamp 1680363874
transform 1 0 268 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3800
timestamp 1680363874
transform 1 0 260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1680363874
transform 1 0 292 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3463
timestamp 1680363874
transform 1 0 316 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1680363874
transform 1 0 340 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3802
timestamp 1680363874
transform 1 0 324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1680363874
transform 1 0 340 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1680363874
transform 1 0 316 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1680363874
transform 1 0 324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1680363874
transform 1 0 348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1680363874
transform 1 0 396 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3464
timestamp 1680363874
transform 1 0 460 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1680363874
transform 1 0 564 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3793
timestamp 1680363874
transform 1 0 484 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3488
timestamp 1680363874
transform 1 0 484 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3885
timestamp 1680363874
transform 1 0 572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1680363874
transform 1 0 580 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3421
timestamp 1680363874
transform 1 0 612 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1680363874
transform 1 0 676 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3805
timestamp 1680363874
transform 1 0 596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1680363874
transform 1 0 612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1680363874
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3400
timestamp 1680363874
transform 1 0 804 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1680363874
transform 1 0 796 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3807
timestamp 1680363874
transform 1 0 796 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1680363874
transform 1 0 708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1680363874
transform 1 0 716 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1680363874
transform 1 0 748 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3401
timestamp 1680363874
transform 1 0 836 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1680363874
transform 1 0 844 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3808
timestamp 1680363874
transform 1 0 860 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3415
timestamp 1680363874
transform 1 0 892 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1680363874
transform 1 0 884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1680363874
transform 1 0 900 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3809
timestamp 1680363874
transform 1 0 900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1680363874
transform 1 0 908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1680363874
transform 1 0 924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1680363874
transform 1 0 932 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3515
timestamp 1680363874
transform 1 0 924 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1680363874
transform 1 0 956 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1680363874
transform 1 0 956 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1680363874
transform 1 0 972 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3810
timestamp 1680363874
transform 1 0 980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1680363874
transform 1 0 996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1680363874
transform 1 0 988 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3490
timestamp 1680363874
transform 1 0 996 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3895
timestamp 1680363874
transform 1 0 1028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1680363874
transform 1 0 1036 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3516
timestamp 1680363874
transform 1 0 1028 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1680363874
transform 1 0 1084 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3812
timestamp 1680363874
transform 1 0 1084 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1680363874
transform 1 0 1084 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3428
timestamp 1680363874
transform 1 0 1124 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3813
timestamp 1680363874
transform 1 0 1116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1680363874
transform 1 0 1108 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3525
timestamp 1680363874
transform 1 0 1108 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1680363874
transform 1 0 1124 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3972
timestamp 1680363874
transform 1 0 1124 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3517
timestamp 1680363874
transform 1 0 1140 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1680363874
transform 1 0 1156 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3899
timestamp 1680363874
transform 1 0 1188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1680363874
transform 1 0 1196 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3527
timestamp 1680363874
transform 1 0 1188 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1680363874
transform 1 0 1212 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1680363874
transform 1 0 1260 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3518
timestamp 1680363874
transform 1 0 1260 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3980
timestamp 1680363874
transform 1 0 1260 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1680363874
transform 1 0 1268 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1680363874
transform 1 0 1284 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3528
timestamp 1680363874
transform 1 0 1284 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3901
timestamp 1680363874
transform 1 0 1412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1680363874
transform 1 0 1476 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3529
timestamp 1680363874
transform 1 0 1476 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3902
timestamp 1680363874
transform 1 0 1492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1680363874
transform 1 0 1508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1680363874
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3530
timestamp 1680363874
transform 1 0 1508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1680363874
transform 1 0 1556 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3815
timestamp 1680363874
transform 1 0 1548 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1680363874
transform 1 0 1556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1680363874
transform 1 0 1572 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3491
timestamp 1680363874
transform 1 0 1548 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1680363874
transform 1 0 1580 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3905
timestamp 1680363874
transform 1 0 1556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1680363874
transform 1 0 1564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1680363874
transform 1 0 1580 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3531
timestamp 1680363874
transform 1 0 1564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1680363874
transform 1 0 1596 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1680363874
transform 1 0 1620 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3818
timestamp 1680363874
transform 1 0 1620 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3432
timestamp 1680363874
transform 1 0 1644 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1680363874
transform 1 0 1636 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3819
timestamp 1680363874
transform 1 0 1644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1680363874
transform 1 0 1628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1680363874
transform 1 0 1636 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3402
timestamp 1680363874
transform 1 0 1676 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3820
timestamp 1680363874
transform 1 0 1692 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3403
timestamp 1680363874
transform 1 0 1716 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1680363874
transform 1 0 1724 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3875
timestamp 1680363874
transform 1 0 1708 0 1 2933
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1680363874
transform 1 0 1716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1680363874
transform 1 0 1684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1680363874
transform 1 0 1700 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3532
timestamp 1680363874
transform 1 0 1700 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1680363874
transform 1 0 1716 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1680363874
transform 1 0 1708 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1680363874
transform 1 0 1764 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3822
timestamp 1680363874
transform 1 0 1748 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1680363874
transform 1 0 1764 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3492
timestamp 1680363874
transform 1 0 1748 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3912
timestamp 1680363874
transform 1 0 1756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1680363874
transform 1 0 1772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1680363874
transform 1 0 1780 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3435
timestamp 1680363874
transform 1 0 1844 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1680363874
transform 1 0 1860 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3824
timestamp 1680363874
transform 1 0 1844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1680363874
transform 1 0 1884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1680363874
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1680363874
transform 1 0 1956 0 1 2933
box -2 -2 2 2
use M3_M2  M3_M2_3493
timestamp 1680363874
transform 1 0 1956 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3916
timestamp 1680363874
transform 1 0 1980 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1680363874
transform 1 0 2036 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3437
timestamp 1680363874
transform 1 0 2076 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3825
timestamp 1680363874
transform 1 0 2076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1680363874
transform 1 0 2060 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3494
timestamp 1680363874
transform 1 0 2068 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1680363874
transform 1 0 2092 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3826
timestamp 1680363874
transform 1 0 2092 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3438
timestamp 1680363874
transform 1 0 2108 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3919
timestamp 1680363874
transform 1 0 2100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1680363874
transform 1 0 2124 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3495
timestamp 1680363874
transform 1 0 2124 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3920
timestamp 1680363874
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1680363874
transform 1 0 2164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1680363874
transform 1 0 2188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1680363874
transform 1 0 2212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1680363874
transform 1 0 2220 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3469
timestamp 1680363874
transform 1 0 2260 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3922
timestamp 1680363874
transform 1 0 2260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1680363874
transform 1 0 2268 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3534
timestamp 1680363874
transform 1 0 2252 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1680363874
transform 1 0 2292 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1680363874
transform 1 0 2324 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3831
timestamp 1680363874
transform 1 0 2300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1680363874
transform 1 0 2308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1680363874
transform 1 0 2324 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3496
timestamp 1680363874
transform 1 0 2284 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1680363874
transform 1 0 2308 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3924
timestamp 1680363874
transform 1 0 2316 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3498
timestamp 1680363874
transform 1 0 2324 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1680363874
transform 1 0 2340 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3925
timestamp 1680363874
transform 1 0 2340 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3472
timestamp 1680363874
transform 1 0 2356 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3834
timestamp 1680363874
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3440
timestamp 1680363874
transform 1 0 2476 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3835
timestamp 1680363874
transform 1 0 2476 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3499
timestamp 1680363874
transform 1 0 2396 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3926
timestamp 1680363874
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3552
timestamp 1680363874
transform 1 0 2412 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1680363874
transform 1 0 2468 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1680363874
transform 1 0 2492 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3927
timestamp 1680363874
transform 1 0 2492 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3535
timestamp 1680363874
transform 1 0 2492 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1680363874
transform 1 0 2524 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3836
timestamp 1680363874
transform 1 0 2508 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3474
timestamp 1680363874
transform 1 0 2516 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3837
timestamp 1680363874
transform 1 0 2540 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3475
timestamp 1680363874
transform 1 0 2548 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3928
timestamp 1680363874
transform 1 0 2548 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1680363874
transform 1 0 2564 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3536
timestamp 1680363874
transform 1 0 2564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1680363874
transform 1 0 2580 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3838
timestamp 1680363874
transform 1 0 2580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1680363874
transform 1 0 2596 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3443
timestamp 1680363874
transform 1 0 2636 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3840
timestamp 1680363874
transform 1 0 2620 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3476
timestamp 1680363874
transform 1 0 2628 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3841
timestamp 1680363874
transform 1 0 2636 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1680363874
transform 1 0 2628 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3500
timestamp 1680363874
transform 1 0 2636 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3931
timestamp 1680363874
transform 1 0 2644 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3501
timestamp 1680363874
transform 1 0 2652 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1680363874
transform 1 0 2644 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1680363874
transform 1 0 2684 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3842
timestamp 1680363874
transform 1 0 2684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1680363874
transform 1 0 2700 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3477
timestamp 1680363874
transform 1 0 2708 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3844
timestamp 1680363874
transform 1 0 2716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1680363874
transform 1 0 2708 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3551
timestamp 1680363874
transform 1 0 2684 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1680363874
transform 1 0 2716 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3933
timestamp 1680363874
transform 1 0 2740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1680363874
transform 1 0 2772 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3478
timestamp 1680363874
transform 1 0 2780 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1680363874
transform 1 0 2796 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3846
timestamp 1680363874
transform 1 0 2788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1680363874
transform 1 0 2780 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3444
timestamp 1680363874
transform 1 0 2836 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3847
timestamp 1680363874
transform 1 0 2836 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3445
timestamp 1680363874
transform 1 0 2868 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3935
timestamp 1680363874
transform 1 0 2868 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3479
timestamp 1680363874
transform 1 0 2900 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3795
timestamp 1680363874
transform 1 0 2916 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1680363874
transform 1 0 2908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1680363874
transform 1 0 2916 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3538
timestamp 1680363874
transform 1 0 2916 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1680363874
transform 1 0 2932 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1680363874
transform 1 0 2948 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1680363874
transform 1 0 2932 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3936
timestamp 1680363874
transform 1 0 2932 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3447
timestamp 1680363874
transform 1 0 2956 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3977
timestamp 1680363874
transform 1 0 2948 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3539
timestamp 1680363874
transform 1 0 2948 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1680363874
transform 1 0 2972 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3849
timestamp 1680363874
transform 1 0 3012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1680363874
transform 1 0 3020 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3480
timestamp 1680363874
transform 1 0 3076 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3937
timestamp 1680363874
transform 1 0 3076 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1680363874
transform 1 0 3092 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3554
timestamp 1680363874
transform 1 0 3084 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1680363874
transform 1 0 3132 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3851
timestamp 1680363874
transform 1 0 3156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1680363874
transform 1 0 3252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1680363874
transform 1 0 3268 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3448
timestamp 1680363874
transform 1 0 3292 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1680363874
transform 1 0 3284 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3853
timestamp 1680363874
transform 1 0 3300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1680363874
transform 1 0 3292 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3503
timestamp 1680363874
transform 1 0 3300 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1680363874
transform 1 0 3316 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3854
timestamp 1680363874
transform 1 0 3316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1680363874
transform 1 0 3308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1680363874
transform 1 0 3324 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3504
timestamp 1680363874
transform 1 0 3356 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3942
timestamp 1680363874
transform 1 0 3380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1680363874
transform 1 0 3396 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1680363874
transform 1 0 3420 0 1 2955
box -2 -2 2 2
use M3_M2  M3_M2_3450
timestamp 1680363874
transform 1 0 3460 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3855
timestamp 1680363874
transform 1 0 3460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1680363874
transform 1 0 3452 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3451
timestamp 1680363874
transform 1 0 3476 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3944
timestamp 1680363874
transform 1 0 3476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1680363874
transform 1 0 3484 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3409
timestamp 1680363874
transform 1 0 3572 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1680363874
transform 1 0 3588 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3856
timestamp 1680363874
transform 1 0 3588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1680363874
transform 1 0 3556 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3505
timestamp 1680363874
transform 1 0 3588 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3857
timestamp 1680363874
transform 1 0 3620 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3453
timestamp 1680363874
transform 1 0 3652 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3858
timestamp 1680363874
transform 1 0 3676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1680363874
transform 1 0 3636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1680363874
transform 1 0 3652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1680363874
transform 1 0 3668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1680363874
transform 1 0 3684 0 1 2955
box -2 -2 2 2
use M3_M2  M3_M2_3540
timestamp 1680363874
transform 1 0 3676 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1680363874
transform 1 0 3700 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3859
timestamp 1680363874
transform 1 0 3700 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3482
timestamp 1680363874
transform 1 0 3748 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1680363874
transform 1 0 3788 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3860
timestamp 1680363874
transform 1 0 3836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1680363874
transform 1 0 3748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1680363874
transform 1 0 3756 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3506
timestamp 1680363874
transform 1 0 3772 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3952
timestamp 1680363874
transform 1 0 3788 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3507
timestamp 1680363874
transform 1 0 3836 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1680363874
transform 1 0 3756 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1680363874
transform 1 0 3844 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1680363874
transform 1 0 3948 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1680363874
transform 1 0 3868 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3861
timestamp 1680363874
transform 1 0 3948 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1680363874
transform 1 0 3860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1680363874
transform 1 0 3916 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3485
timestamp 1680363874
transform 1 0 3964 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3955
timestamp 1680363874
transform 1 0 3964 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3410
timestamp 1680363874
transform 1 0 3980 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1680363874
transform 1 0 4044 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1680363874
transform 1 0 4052 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3862
timestamp 1680363874
transform 1 0 4052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1680363874
transform 1 0 4028 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3457
timestamp 1680363874
transform 1 0 4076 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1680363874
transform 1 0 4092 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3863
timestamp 1680363874
transform 1 0 4092 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3508
timestamp 1680363874
transform 1 0 4092 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3957
timestamp 1680363874
transform 1 0 4116 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3509
timestamp 1680363874
transform 1 0 4140 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3796
timestamp 1680363874
transform 1 0 4204 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3486
timestamp 1680363874
transform 1 0 4204 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3864
timestamp 1680363874
transform 1 0 4236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1680363874
transform 1 0 4236 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3543
timestamp 1680363874
transform 1 0 4244 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3865
timestamp 1680363874
transform 1 0 4252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1680363874
transform 1 0 4292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1680363874
transform 1 0 4260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1680363874
transform 1 0 4276 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1680363874
transform 1 0 4276 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3961
timestamp 1680363874
transform 1 0 4308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1680363874
transform 1 0 4372 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3544
timestamp 1680363874
transform 1 0 4364 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1680363874
transform 1 0 4380 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3868
timestamp 1680363874
transform 1 0 4388 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1680363874
transform 1 0 4380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1680363874
transform 1 0 4396 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3520
timestamp 1680363874
transform 1 0 4380 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1680363874
transform 1 0 4396 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3964
timestamp 1680363874
transform 1 0 4412 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3458
timestamp 1680363874
transform 1 0 4444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1680363874
transform 1 0 4532 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3869
timestamp 1680363874
transform 1 0 4532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1680363874
transform 1 0 4508 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3521
timestamp 1680363874
transform 1 0 4532 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1680363874
transform 1 0 4556 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1680363874
transform 1 0 4572 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1680363874
transform 1 0 4588 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1680363874
transform 1 0 4604 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3979
timestamp 1680363874
transform 1 0 4604 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1680363874
transform 1 0 4628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1680363874
transform 1 0 4636 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1680363874
transform 1 0 4652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1680363874
transform 1 0 4660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1680363874
transform 1 0 4644 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3511
timestamp 1680363874
transform 1 0 4652 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3967
timestamp 1680363874
transform 1 0 4660 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3460
timestamp 1680363874
transform 1 0 4788 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3874
timestamp 1680363874
transform 1 0 4788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1680363874
transform 1 0 4700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1680363874
transform 1 0 4708 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3512
timestamp 1680363874
transform 1 0 4716 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3970
timestamp 1680363874
transform 1 0 4756 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3523
timestamp 1680363874
transform 1 0 4700 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1680363874
transform 1 0 4756 0 1 2915
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_36
timestamp 1680363874
transform 1 0 24 0 1 2870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_244
timestamp 1680363874
transform 1 0 72 0 -1 2970
box -8 -3 104 105
use NAND2X1  NAND2X1_32
timestamp 1680363874
transform 1 0 168 0 -1 2970
box -8 -3 32 105
use INVX2  INVX2_259
timestamp 1680363874
transform -1 0 208 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3622
timestamp 1680363874
transform 1 0 208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1680363874
transform 1 0 216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1680363874
transform 1 0 224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1680363874
transform 1 0 232 0 -1 2970
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1680363874
transform -1 0 272 0 -1 2970
box -7 -3 39 105
use FILL  FILL_3626
timestamp 1680363874
transform 1 0 272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1680363874
transform 1 0 280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1680363874
transform 1 0 288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1680363874
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1680363874
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1680363874
transform 1 0 312 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_208
timestamp 1680363874
transform 1 0 320 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3645
timestamp 1680363874
transform 1 0 360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1680363874
transform 1 0 368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1680363874
transform 1 0 376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1680363874
transform 1 0 384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1680363874
transform 1 0 392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1680363874
transform 1 0 400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1680363874
transform 1 0 408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1680363874
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1680363874
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1680363874
transform 1 0 432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1680363874
transform 1 0 440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1680363874
transform 1 0 448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1680363874
transform 1 0 456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1680363874
transform 1 0 464 0 -1 2970
box -8 -3 16 105
use FAX1  FAX1_1
timestamp 1680363874
transform -1 0 592 0 -1 2970
box -5 -3 126 105
use FILL  FILL_3659
timestamp 1680363874
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1680363874
transform 1 0 600 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3671
timestamp 1680363874
transform 1 0 696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1680363874
transform 1 0 704 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3556
timestamp 1680363874
transform 1 0 788 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1680363874
transform 1 0 812 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_247
timestamp 1680363874
transform -1 0 808 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3673
timestamp 1680363874
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1680363874
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1680363874
transform 1 0 824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1680363874
transform 1 0 832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1680363874
transform 1 0 840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1680363874
transform 1 0 848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1680363874
transform 1 0 856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1680363874
transform 1 0 864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1680363874
transform 1 0 872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1680363874
transform 1 0 880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1680363874
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1680363874
transform 1 0 896 0 -1 2970
box -8 -3 40 105
use FILL  FILL_3691
timestamp 1680363874
transform 1 0 928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1680363874
transform 1 0 936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1680363874
transform 1 0 944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1680363874
transform 1 0 952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1680363874
transform 1 0 960 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_133
timestamp 1680363874
transform 1 0 968 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3705
timestamp 1680363874
transform 1 0 1008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1680363874
transform 1 0 1016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1680363874
transform 1 0 1024 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_262
timestamp 1680363874
transform -1 0 1048 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3708
timestamp 1680363874
transform 1 0 1048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1680363874
transform 1 0 1056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1680363874
transform 1 0 1064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1680363874
transform 1 0 1072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1680363874
transform 1 0 1080 0 -1 2970
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1680363874
transform -1 0 1120 0 -1 2970
box -8 -3 40 105
use FILL  FILL_3715
timestamp 1680363874
transform 1 0 1120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1680363874
transform 1 0 1128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1680363874
transform 1 0 1136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1680363874
transform 1 0 1144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1680363874
transform 1 0 1152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1680363874
transform 1 0 1160 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1680363874
transform -1 0 1200 0 -1 2970
box -8 -3 40 105
use FILL  FILL_3728
timestamp 1680363874
transform 1 0 1200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1680363874
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1680363874
transform 1 0 1216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1680363874
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1680363874
transform 1 0 1232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1680363874
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1680363874
transform 1 0 1248 0 -1 2970
box -8 -3 40 105
use FILL  FILL_3737
timestamp 1680363874
transform 1 0 1280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1680363874
transform 1 0 1288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1680363874
transform 1 0 1296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1680363874
transform 1 0 1304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1680363874
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1680363874
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1680363874
transform 1 0 1328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1680363874
transform 1 0 1336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1680363874
transform 1 0 1344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1680363874
transform 1 0 1352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1680363874
transform 1 0 1360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1680363874
transform 1 0 1368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1680363874
transform 1 0 1376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1680363874
transform 1 0 1384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1680363874
transform 1 0 1392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1680363874
transform 1 0 1400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1680363874
transform 1 0 1408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1680363874
transform 1 0 1416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1680363874
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1680363874
transform 1 0 1432 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_266
timestamp 1680363874
transform -1 0 1456 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3769
timestamp 1680363874
transform 1 0 1456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1680363874
transform 1 0 1464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1680363874
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1680363874
transform 1 0 1480 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_136
timestamp 1680363874
transform 1 0 1488 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3777
timestamp 1680363874
transform 1 0 1528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1680363874
transform 1 0 1536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1680363874
transform 1 0 1544 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_209
timestamp 1680363874
transform 1 0 1552 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3790
timestamp 1680363874
transform 1 0 1592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1680363874
transform 1 0 1600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1680363874
transform 1 0 1608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1680363874
transform 1 0 1616 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_270
timestamp 1680363874
transform 1 0 1624 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3794
timestamp 1680363874
transform 1 0 1640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1680363874
transform 1 0 1648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1680363874
transform 1 0 1656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1680363874
transform 1 0 1664 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_210
timestamp 1680363874
transform -1 0 1712 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3798
timestamp 1680363874
transform 1 0 1712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1680363874
transform 1 0 1720 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_211
timestamp 1680363874
transform 1 0 1728 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3800
timestamp 1680363874
transform 1 0 1768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1680363874
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1680363874
transform 1 0 1784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1680363874
transform 1 0 1792 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_271
timestamp 1680363874
transform 1 0 1800 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3804
timestamp 1680363874
transform 1 0 1816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1680363874
transform 1 0 1824 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1680363874
transform 1 0 1832 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3806
timestamp 1680363874
transform 1 0 1928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1680363874
transform 1 0 1936 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_253
timestamp 1680363874
transform 1 0 1944 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3808
timestamp 1680363874
transform 1 0 2040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1680363874
transform 1 0 2048 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_15
timestamp 1680363874
transform 1 0 2056 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3814
timestamp 1680363874
transform 1 0 2080 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_272
timestamp 1680363874
transform 1 0 2088 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3815
timestamp 1680363874
transform 1 0 2104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1680363874
transform 1 0 2112 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_16
timestamp 1680363874
transform -1 0 2144 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1680363874
transform 1 0 2144 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3817
timestamp 1680363874
transform 1 0 2168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1680363874
transform 1 0 2176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1680363874
transform 1 0 2184 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_18
timestamp 1680363874
transform 1 0 2192 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3830
timestamp 1680363874
transform 1 0 2216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1680363874
transform 1 0 2224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1680363874
transform 1 0 2232 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3558
timestamp 1680363874
transform 1 0 2260 0 1 2875
box -3 -3 3 3
use BUFX2  BUFX2_19
timestamp 1680363874
transform -1 0 2264 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3833
timestamp 1680363874
transform 1 0 2264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1680363874
transform 1 0 2272 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_20
timestamp 1680363874
transform 1 0 2280 0 -1 2970
box -5 -3 28 105
use INVX2  INVX2_273
timestamp 1680363874
transform 1 0 2304 0 -1 2970
box -9 -3 26 105
use BUFX2  BUFX2_21
timestamp 1680363874
transform -1 0 2344 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3835
timestamp 1680363874
transform 1 0 2344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1680363874
transform 1 0 2352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1680363874
transform 1 0 2360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1680363874
transform 1 0 2368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1680363874
transform 1 0 2376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1680363874
transform 1 0 2384 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1680363874
transform -1 0 2488 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3851
timestamp 1680363874
transform 1 0 2488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1680363874
transform 1 0 2496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1680363874
transform 1 0 2504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1680363874
transform 1 0 2512 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_212
timestamp 1680363874
transform 1 0 2520 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3860
timestamp 1680363874
transform 1 0 2560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1680363874
transform 1 0 2568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1680363874
transform 1 0 2576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1680363874
transform 1 0 2584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1680363874
transform 1 0 2592 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_213
timestamp 1680363874
transform 1 0 2600 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3865
timestamp 1680363874
transform 1 0 2640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1680363874
transform 1 0 2648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1680363874
transform 1 0 2656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1680363874
transform 1 0 2664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1680363874
transform 1 0 2672 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_214
timestamp 1680363874
transform 1 0 2680 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3876
timestamp 1680363874
transform 1 0 2720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1680363874
transform 1 0 2728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1680363874
transform 1 0 2736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1680363874
transform 1 0 2744 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_22
timestamp 1680363874
transform 1 0 2752 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3880
timestamp 1680363874
transform 1 0 2776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1680363874
transform 1 0 2784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1680363874
transform 1 0 2792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1680363874
transform 1 0 2800 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_278
timestamp 1680363874
transform 1 0 2808 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3887
timestamp 1680363874
transform 1 0 2824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1680363874
transform 1 0 2832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1680363874
transform 1 0 2840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1680363874
transform 1 0 2848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1680363874
transform 1 0 2856 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_107
timestamp 1680363874
transform 1 0 2864 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3897
timestamp 1680363874
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1680363874
transform 1 0 2904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1680363874
transform 1 0 2912 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_109
timestamp 1680363874
transform 1 0 2920 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3906
timestamp 1680363874
transform 1 0 2952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1680363874
transform 1 0 2960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1680363874
transform 1 0 2968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1680363874
transform 1 0 2976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1680363874
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1680363874
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1680363874
transform 1 0 3000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1680363874
transform 1 0 3008 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_23
timestamp 1680363874
transform -1 0 3040 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3922
timestamp 1680363874
transform 1 0 3040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1680363874
transform 1 0 3048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1680363874
transform 1 0 3056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1680363874
transform 1 0 3064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1680363874
transform 1 0 3072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1680363874
transform 1 0 3080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1680363874
transform 1 0 3088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1680363874
transform 1 0 3096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1680363874
transform 1 0 3104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1680363874
transform 1 0 3112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1680363874
transform 1 0 3120 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_279
timestamp 1680363874
transform -1 0 3144 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3934
timestamp 1680363874
transform 1 0 3144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1680363874
transform 1 0 3152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1680363874
transform 1 0 3160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1680363874
transform 1 0 3168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1680363874
transform 1 0 3176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1680363874
transform 1 0 3184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1680363874
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1680363874
transform 1 0 3200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1680363874
transform 1 0 3208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1680363874
transform 1 0 3216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1680363874
transform 1 0 3224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1680363874
transform 1 0 3232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1680363874
transform 1 0 3240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1680363874
transform 1 0 3248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1680363874
transform 1 0 3256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1680363874
transform 1 0 3264 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_137
timestamp 1680363874
transform -1 0 3312 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3967
timestamp 1680363874
transform 1 0 3312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1680363874
transform 1 0 3320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1680363874
transform 1 0 3328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1680363874
transform 1 0 3336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1680363874
transform 1 0 3344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1680363874
transform 1 0 3352 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3559
timestamp 1680363874
transform 1 0 3380 0 1 2875
box -3 -3 3 3
use INVX2  INVX2_280
timestamp 1680363874
transform 1 0 3360 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3975
timestamp 1680363874
transform 1 0 3376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1680363874
transform 1 0 3384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1680363874
transform 1 0 3392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1680363874
transform 1 0 3400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1680363874
transform 1 0 3408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1680363874
transform 1 0 3416 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_26
timestamp 1680363874
transform 1 0 3424 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3993
timestamp 1680363874
transform 1 0 3448 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_27
timestamp 1680363874
transform -1 0 3480 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3994
timestamp 1680363874
transform 1 0 3480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1680363874
transform 1 0 3488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1680363874
transform 1 0 3496 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1680363874
transform -1 0 3600 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3997
timestamp 1680363874
transform 1 0 3600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1680363874
transform 1 0 3608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1680363874
transform 1 0 3616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1680363874
transform 1 0 3624 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_139
timestamp 1680363874
transform 1 0 3632 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4011
timestamp 1680363874
transform 1 0 3672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1680363874
transform 1 0 3680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1680363874
transform 1 0 3688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1680363874
transform 1 0 3696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1680363874
transform 1 0 3704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1680363874
transform 1 0 3712 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_282
timestamp 1680363874
transform 1 0 3720 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4017
timestamp 1680363874
transform 1 0 3736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1680363874
transform 1 0 3744 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_263
timestamp 1680363874
transform -1 0 3848 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4042
timestamp 1680363874
transform 1 0 3848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1680363874
transform 1 0 3856 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1680363874
transform -1 0 3960 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4044
timestamp 1680363874
transform 1 0 3960 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1680363874
transform -1 0 4064 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4045
timestamp 1680363874
transform 1 0 4064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1680363874
transform 1 0 4072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1680363874
transform 1 0 4080 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_283
timestamp 1680363874
transform 1 0 4088 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4050
timestamp 1680363874
transform 1 0 4104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1680363874
transform 1 0 4112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1680363874
transform 1 0 4120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1680363874
transform 1 0 4128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1680363874
transform 1 0 4136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1680363874
transform 1 0 4144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1680363874
transform 1 0 4152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1680363874
transform 1 0 4160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1680363874
transform 1 0 4168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1680363874
transform 1 0 4176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1680363874
transform 1 0 4184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1680363874
transform 1 0 4192 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_37
timestamp 1680363874
transform 1 0 4200 0 -1 2970
box -8 -3 32 105
use FILL  FILL_4065
timestamp 1680363874
transform 1 0 4224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1680363874
transform 1 0 4232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1680363874
transform 1 0 4240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1680363874
transform 1 0 4248 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_140
timestamp 1680363874
transform -1 0 4296 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4075
timestamp 1680363874
transform 1 0 4296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1680363874
transform 1 0 4304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1680363874
transform 1 0 4312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1680363874
transform 1 0 4320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1680363874
transform 1 0 4328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1680363874
transform 1 0 4336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1680363874
transform 1 0 4344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1680363874
transform 1 0 4352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1680363874
transform 1 0 4360 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_215
timestamp 1680363874
transform 1 0 4368 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4091
timestamp 1680363874
transform 1 0 4408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1680363874
transform 1 0 4416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1680363874
transform 1 0 4424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1680363874
transform 1 0 4432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1680363874
transform 1 0 4440 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_267
timestamp 1680363874
transform -1 0 4544 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4110
timestamp 1680363874
transform 1 0 4544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1680363874
transform 1 0 4552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1680363874
transform 1 0 4560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1680363874
transform 1 0 4568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1680363874
transform 1 0 4576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1680363874
transform 1 0 4584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1680363874
transform 1 0 4592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1680363874
transform 1 0 4600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1680363874
transform 1 0 4608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1680363874
transform 1 0 4616 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_143
timestamp 1680363874
transform 1 0 4624 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4125
timestamp 1680363874
transform 1 0 4664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1680363874
transform 1 0 4672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1680363874
transform 1 0 4680 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_286
timestamp 1680363874
transform 1 0 4688 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1680363874
transform -1 0 4800 0 -1 2970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_37
timestamp 1680363874
transform 1 0 4851 0 1 2870
box -10 -3 10 3
use M2_M1  M2_M1_3991
timestamp 1680363874
transform 1 0 100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1680363874
transform 1 0 124 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3739
timestamp 1680363874
transform 1 0 124 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4205
timestamp 1680363874
transform 1 0 156 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3576
timestamp 1680363874
transform 1 0 188 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3992
timestamp 1680363874
transform 1 0 180 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3671
timestamp 1680363874
transform 1 0 180 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3993
timestamp 1680363874
transform 1 0 204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1680363874
transform 1 0 188 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3740
timestamp 1680363874
transform 1 0 196 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1680363874
transform 1 0 228 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1680363874
transform 1 0 260 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1680363874
transform 1 0 260 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1680363874
transform 1 0 276 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1680363874
transform 1 0 252 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3994
timestamp 1680363874
transform 1 0 260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1680363874
transform 1 0 276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1680363874
transform 1 0 252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1680363874
transform 1 0 244 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3672
timestamp 1680363874
transform 1 0 260 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4105
timestamp 1680363874
transform 1 0 268 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3611
timestamp 1680363874
transform 1 0 300 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3996
timestamp 1680363874
transform 1 0 300 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3702
timestamp 1680363874
transform 1 0 292 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1680363874
transform 1 0 324 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1680363874
transform 1 0 316 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4106
timestamp 1680363874
transform 1 0 316 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3648
timestamp 1680363874
transform 1 0 332 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4107
timestamp 1680363874
transform 1 0 332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1680363874
transform 1 0 396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1680363874
transform 1 0 412 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3741
timestamp 1680363874
transform 1 0 412 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1680363874
transform 1 0 444 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3998
timestamp 1680363874
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1680363874
transform 1 0 444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1680363874
transform 1 0 444 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3742
timestamp 1680363874
transform 1 0 444 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4108
timestamp 1680363874
transform 1 0 492 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1680363874
transform 1 0 508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1680363874
transform 1 0 524 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1680363874
transform 1 0 532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1680363874
transform 1 0 564 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3614
timestamp 1680363874
transform 1 0 588 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4001
timestamp 1680363874
transform 1 0 588 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3673
timestamp 1680363874
transform 1 0 572 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1680363874
transform 1 0 596 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1680363874
transform 1 0 596 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1680363874
transform 1 0 636 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1680363874
transform 1 0 652 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3982
timestamp 1680363874
transform 1 0 660 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1680363874
transform 1 0 652 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1680363874
transform 1 0 660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1680363874
transform 1 0 668 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3592
timestamp 1680363874
transform 1 0 692 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4002
timestamp 1680363874
transform 1 0 684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1680363874
transform 1 0 692 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3675
timestamp 1680363874
transform 1 0 684 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1680363874
transform 1 0 700 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1680363874
transform 1 0 740 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4004
timestamp 1680363874
transform 1 0 740 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3677
timestamp 1680363874
transform 1 0 732 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4112
timestamp 1680363874
transform 1 0 748 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3703
timestamp 1680363874
transform 1 0 740 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4005
timestamp 1680363874
transform 1 0 780 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3678
timestamp 1680363874
transform 1 0 780 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1680363874
transform 1 0 804 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4006
timestamp 1680363874
transform 1 0 812 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3650
timestamp 1680363874
transform 1 0 820 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4113
timestamp 1680363874
transform 1 0 796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1680363874
transform 1 0 804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1680363874
transform 1 0 820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1680363874
transform 1 0 828 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3617
timestamp 1680363874
transform 1 0 844 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4007
timestamp 1680363874
transform 1 0 844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1680363874
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3744
timestamp 1680363874
transform 1 0 876 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1680363874
transform 1 0 916 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4008
timestamp 1680363874
transform 1 0 908 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1680363874
transform 1 0 916 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3679
timestamp 1680363874
transform 1 0 916 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1680363874
transform 1 0 916 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4010
timestamp 1680363874
transform 1 0 932 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1680363874
transform 1 0 948 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3651
timestamp 1680363874
transform 1 0 964 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4118
timestamp 1680363874
transform 1 0 956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1680363874
transform 1 0 964 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3705
timestamp 1680363874
transform 1 0 964 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4012
timestamp 1680363874
transform 1 0 980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1680363874
transform 1 0 1084 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1680363874
transform 1 0 1092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1680363874
transform 1 0 1100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1680363874
transform 1 0 1140 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3564
timestamp 1680363874
transform 1 0 1260 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4017
timestamp 1680363874
transform 1 0 1220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1680363874
transform 1 0 1100 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1680363874
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1680363874
transform 1 0 1156 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1680363874
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1680363874
transform 1 0 996 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3706
timestamp 1680363874
transform 1 0 1044 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1680363874
transform 1 0 1100 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1680363874
transform 1 0 996 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1680363874
transform 1 0 1124 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1680363874
transform 1 0 1220 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1680363874
transform 1 0 1196 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1680363874
transform 1 0 1284 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4124
timestamp 1680363874
transform 1 0 1284 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3565
timestamp 1680363874
transform 1 0 1308 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1680363874
transform 1 0 1300 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1680363874
transform 1 0 1324 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4018
timestamp 1680363874
transform 1 0 1300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1680363874
transform 1 0 1308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1680363874
transform 1 0 1324 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3681
timestamp 1680363874
transform 1 0 1308 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4125
timestamp 1680363874
transform 1 0 1316 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3566
timestamp 1680363874
transform 1 0 1340 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4021
timestamp 1680363874
transform 1 0 1340 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3578
timestamp 1680363874
transform 1 0 1348 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1680363874
transform 1 0 1380 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_4022
timestamp 1680363874
transform 1 0 1404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1680363874
transform 1 0 1372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1680363874
transform 1 0 1380 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1680363874
transform 1 0 1396 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1680363874
transform 1 0 1412 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3708
timestamp 1680363874
transform 1 0 1372 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1680363874
transform 1 0 1412 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1680363874
transform 1 0 1580 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1680363874
transform 1 0 1556 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_4023
timestamp 1680363874
transform 1 0 1572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1680363874
transform 1 0 1540 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3682
timestamp 1680363874
transform 1 0 1572 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1680363874
transform 1 0 1612 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1680363874
transform 1 0 1612 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1680363874
transform 1 0 1540 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4024
timestamp 1680363874
transform 1 0 1628 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3749
timestamp 1680363874
transform 1 0 1636 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4131
timestamp 1680363874
transform 1 0 1660 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3561
timestamp 1680363874
transform 1 0 1716 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1680363874
transform 1 0 1708 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1680363874
transform 1 0 1700 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4025
timestamp 1680363874
transform 1 0 1692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1680363874
transform 1 0 1708 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3652
timestamp 1680363874
transform 1 0 1716 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4132
timestamp 1680363874
transform 1 0 1700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1680363874
transform 1 0 1724 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3622
timestamp 1680363874
transform 1 0 1732 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4027
timestamp 1680363874
transform 1 0 1732 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3711
timestamp 1680363874
transform 1 0 1724 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1680363874
transform 1 0 1748 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4134
timestamp 1680363874
transform 1 0 1756 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1680363874
transform 1 0 1756 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1680363874
transform 1 0 1876 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1680363874
transform 1 0 1908 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4028
timestamp 1680363874
transform 1 0 1772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1680363874
transform 1 0 1828 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3653
timestamp 1680363874
transform 1 0 1868 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4030
timestamp 1680363874
transform 1 0 1876 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1680363874
transform 1 0 1892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1680363874
transform 1 0 1908 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1680363874
transform 1 0 1852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1680363874
transform 1 0 1868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1680363874
transform 1 0 1884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1680363874
transform 1 0 1900 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3750
timestamp 1680363874
transform 1 0 1900 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4139
timestamp 1680363874
transform 1 0 1924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1680363874
transform 1 0 1932 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3713
timestamp 1680363874
transform 1 0 1932 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1680363874
transform 1 0 1972 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1680363874
transform 1 0 1956 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1680363874
transform 1 0 1980 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4033
timestamp 1680363874
transform 1 0 1956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1680363874
transform 1 0 1972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1680363874
transform 1 0 1980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1680363874
transform 1 0 1964 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1680363874
transform 1 0 1980 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3751
timestamp 1680363874
transform 1 0 1980 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4143
timestamp 1680363874
transform 1 0 2036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1680363874
transform 1 0 2044 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3627
timestamp 1680363874
transform 1 0 2060 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4036
timestamp 1680363874
transform 1 0 2060 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3714
timestamp 1680363874
transform 1 0 2052 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4145
timestamp 1680363874
transform 1 0 2084 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3568
timestamp 1680363874
transform 1 0 2100 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1680363874
transform 1 0 2100 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4037
timestamp 1680363874
transform 1 0 2100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1680363874
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3715
timestamp 1680363874
transform 1 0 2124 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1680363874
transform 1 0 2156 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4039
timestamp 1680363874
transform 1 0 2164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1680363874
transform 1 0 2148 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3685
timestamp 1680363874
transform 1 0 2156 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1680363874
transform 1 0 2180 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4147
timestamp 1680363874
transform 1 0 2188 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3716
timestamp 1680363874
transform 1 0 2180 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1680363874
transform 1 0 2212 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4040
timestamp 1680363874
transform 1 0 2220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1680363874
transform 1 0 2212 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3687
timestamp 1680363874
transform 1 0 2220 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1680363874
transform 1 0 2268 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4041
timestamp 1680363874
transform 1 0 2244 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1680363874
transform 1 0 2252 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3656
timestamp 1680363874
transform 1 0 2260 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4043
timestamp 1680363874
transform 1 0 2276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1680363874
transform 1 0 2268 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3630
timestamp 1680363874
transform 1 0 2300 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4044
timestamp 1680363874
transform 1 0 2300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1680363874
transform 1 0 2292 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3631
timestamp 1680363874
transform 1 0 2348 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4151
timestamp 1680363874
transform 1 0 2332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1680363874
transform 1 0 2340 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3596
timestamp 1680363874
transform 1 0 2380 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1680363874
transform 1 0 2380 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4045
timestamp 1680363874
transform 1 0 2380 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3562
timestamp 1680363874
transform 1 0 2396 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_4046
timestamp 1680363874
transform 1 0 2396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1680363874
transform 1 0 2396 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3752
timestamp 1680363874
transform 1 0 2396 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1680363874
transform 1 0 2412 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1680363874
transform 1 0 2404 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4154
timestamp 1680363874
transform 1 0 2412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1680363874
transform 1 0 2420 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3633
timestamp 1680363874
transform 1 0 2436 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4048
timestamp 1680363874
transform 1 0 2436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1680363874
transform 1 0 2452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1680363874
transform 1 0 2444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1680363874
transform 1 0 2468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1680363874
transform 1 0 2468 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3634
timestamp 1680363874
transform 1 0 2492 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4157
timestamp 1680363874
transform 1 0 2484 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3717
timestamp 1680363874
transform 1 0 2524 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4051
timestamp 1680363874
transform 1 0 2540 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3570
timestamp 1680363874
transform 1 0 2596 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1680363874
transform 1 0 2620 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1680363874
transform 1 0 2556 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4052
timestamp 1680363874
transform 1 0 2596 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3658
timestamp 1680363874
transform 1 0 2628 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4158
timestamp 1680363874
transform 1 0 2628 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3718
timestamp 1680363874
transform 1 0 2628 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4053
timestamp 1680363874
transform 1 0 2644 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3598
timestamp 1680363874
transform 1 0 2660 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4159
timestamp 1680363874
transform 1 0 2660 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3719
timestamp 1680363874
transform 1 0 2652 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1680363874
transform 1 0 2676 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1680363874
transform 1 0 2692 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4054
timestamp 1680363874
transform 1 0 2692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1680363874
transform 1 0 2708 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3688
timestamp 1680363874
transform 1 0 2692 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4056
timestamp 1680363874
transform 1 0 2724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1680363874
transform 1 0 2700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1680363874
transform 1 0 2716 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3720
timestamp 1680363874
transform 1 0 2716 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4162
timestamp 1680363874
transform 1 0 2772 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3599
timestamp 1680363874
transform 1 0 2812 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1680363874
transform 1 0 2820 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1680363874
transform 1 0 2836 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4057
timestamp 1680363874
transform 1 0 2812 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1680363874
transform 1 0 2820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1680363874
transform 1 0 2836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1680363874
transform 1 0 2812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1680363874
transform 1 0 2828 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3689
timestamp 1680363874
transform 1 0 2836 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4165
timestamp 1680363874
transform 1 0 2844 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3721
timestamp 1680363874
transform 1 0 2820 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1680363874
transform 1 0 2844 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1680363874
transform 1 0 2884 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4166
timestamp 1680363874
transform 1 0 2884 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3580
timestamp 1680363874
transform 1 0 2900 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1680363874
transform 1 0 2908 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4060
timestamp 1680363874
transform 1 0 2900 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3581
timestamp 1680363874
transform 1 0 2932 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_4061
timestamp 1680363874
transform 1 0 2932 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3582
timestamp 1680363874
transform 1 0 2948 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3983
timestamp 1680363874
transform 1 0 2948 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_3638
timestamp 1680363874
transform 1 0 2948 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4167
timestamp 1680363874
transform 1 0 2948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1680363874
transform 1 0 2972 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3573
timestamp 1680363874
transform 1 0 2988 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4062
timestamp 1680363874
transform 1 0 2988 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3574
timestamp 1680363874
transform 1 0 3012 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1680363874
transform 1 0 3012 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3986
timestamp 1680363874
transform 1 0 3012 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3601
timestamp 1680363874
transform 1 0 3028 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4063
timestamp 1680363874
transform 1 0 3028 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3753
timestamp 1680363874
transform 1 0 3028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1680363874
transform 1 0 3044 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4168
timestamp 1680363874
transform 1 0 3044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1680363874
transform 1 0 3100 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3690
timestamp 1680363874
transform 1 0 3100 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4169
timestamp 1680363874
transform 1 0 3148 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3723
timestamp 1680363874
transform 1 0 3148 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1680363874
transform 1 0 3172 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3987
timestamp 1680363874
transform 1 0 3172 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3724
timestamp 1680363874
transform 1 0 3180 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4065
timestamp 1680363874
transform 1 0 3204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1680363874
transform 1 0 3220 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3691
timestamp 1680363874
transform 1 0 3220 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1680363874
transform 1 0 3244 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1680363874
transform 1 0 3308 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1680363874
transform 1 0 3348 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4067
timestamp 1680363874
transform 1 0 3268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1680363874
transform 1 0 3324 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3692
timestamp 1680363874
transform 1 0 3260 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4170
timestamp 1680363874
transform 1 0 3348 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3726
timestamp 1680363874
transform 1 0 3348 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3988
timestamp 1680363874
transform 1 0 3364 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3640
timestamp 1680363874
transform 1 0 3372 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1680363874
transform 1 0 3364 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4171
timestamp 1680363874
transform 1 0 3364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1680363874
transform 1 0 3388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1680363874
transform 1 0 3396 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3727
timestamp 1680363874
transform 1 0 3396 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4069
timestamp 1680363874
transform 1 0 3420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1680363874
transform 1 0 3436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1680363874
transform 1 0 3484 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1680363874
transform 1 0 3508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1680363874
transform 1 0 3556 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3602
timestamp 1680363874
transform 1 0 3580 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3989
timestamp 1680363874
transform 1 0 3596 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3662
timestamp 1680363874
transform 1 0 3588 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4177
timestamp 1680363874
transform 1 0 3636 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3603
timestamp 1680363874
transform 1 0 3660 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1680363874
transform 1 0 3652 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1680363874
transform 1 0 3668 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4071
timestamp 1680363874
transform 1 0 3660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1680363874
transform 1 0 3668 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3693
timestamp 1680363874
transform 1 0 3660 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1680363874
transform 1 0 3644 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4178
timestamp 1680363874
transform 1 0 3676 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3728
timestamp 1680363874
transform 1 0 3668 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4212
timestamp 1680363874
transform 1 0 3732 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1680363874
transform 1 0 3748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1680363874
transform 1 0 3764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1680363874
transform 1 0 3796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1680363874
transform 1 0 3812 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3663
timestamp 1680363874
transform 1 0 3820 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1680363874
transform 1 0 3836 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4075
timestamp 1680363874
transform 1 0 3836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1680363874
transform 1 0 3796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1680363874
transform 1 0 3804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1680363874
transform 1 0 3820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1680363874
transform 1 0 3828 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3729
timestamp 1680363874
transform 1 0 3804 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1680363874
transform 1 0 3860 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3990
timestamp 1680363874
transform 1 0 3908 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1680363874
transform 1 0 3892 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3694
timestamp 1680363874
transform 1 0 3900 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1680363874
transform 1 0 3892 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4076
timestamp 1680363874
transform 1 0 3916 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1680363874
transform 1 0 3932 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3665
timestamp 1680363874
transform 1 0 3964 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1680363874
transform 1 0 3996 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4078
timestamp 1680363874
transform 1 0 3996 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3666
timestamp 1680363874
transform 1 0 4004 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4186
timestamp 1680363874
transform 1 0 3988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1680363874
transform 1 0 4004 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3731
timestamp 1680363874
transform 1 0 3988 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1680363874
transform 1 0 4020 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4079
timestamp 1680363874
transform 1 0 4020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1680363874
transform 1 0 4028 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3695
timestamp 1680363874
transform 1 0 4028 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1680363874
transform 1 0 4036 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4188
timestamp 1680363874
transform 1 0 4036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1680363874
transform 1 0 4076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1680363874
transform 1 0 4060 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3696
timestamp 1680363874
transform 1 0 4068 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1680363874
transform 1 0 4060 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1680363874
transform 1 0 4076 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1680363874
transform 1 0 4156 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1680363874
transform 1 0 4132 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1680363874
transform 1 0 4132 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4082
timestamp 1680363874
transform 1 0 4140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1680363874
transform 1 0 4156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1680363874
transform 1 0 4132 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3697
timestamp 1680363874
transform 1 0 4140 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4191
timestamp 1680363874
transform 1 0 4148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1680363874
transform 1 0 4164 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1680363874
transform 1 0 4180 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3756
timestamp 1680363874
transform 1 0 4180 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4084
timestamp 1680363874
transform 1 0 4204 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3733
timestamp 1680363874
transform 1 0 4212 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1680363874
transform 1 0 4260 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_4085
timestamp 1680363874
transform 1 0 4244 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1680363874
transform 1 0 4260 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3734
timestamp 1680363874
transform 1 0 4228 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1680363874
transform 1 0 4260 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4193
timestamp 1680363874
transform 1 0 4268 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1680363874
transform 1 0 4300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1680363874
transform 1 0 4292 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3607
timestamp 1680363874
transform 1 0 4332 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4088
timestamp 1680363874
transform 1 0 4332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1680363874
transform 1 0 4340 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3585
timestamp 1680363874
transform 1 0 4420 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1680363874
transform 1 0 4404 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4090
timestamp 1680363874
transform 1 0 4404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1680363874
transform 1 0 4420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1680363874
transform 1 0 4396 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3757
timestamp 1680363874
transform 1 0 4396 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1680363874
transform 1 0 4428 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4092
timestamp 1680363874
transform 1 0 4436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1680363874
transform 1 0 4412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1680363874
transform 1 0 4428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1680363874
transform 1 0 4436 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3735
timestamp 1680363874
transform 1 0 4412 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1680363874
transform 1 0 4452 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1680363874
transform 1 0 4444 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4093
timestamp 1680363874
transform 1 0 4476 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3699
timestamp 1680363874
transform 1 0 4468 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4094
timestamp 1680363874
transform 1 0 4508 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3700
timestamp 1680363874
transform 1 0 4508 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4095
timestamp 1680363874
transform 1 0 4532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1680363874
transform 1 0 4572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1680363874
transform 1 0 4548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1680363874
transform 1 0 4564 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3758
timestamp 1680363874
transform 1 0 4564 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1680363874
transform 1 0 4628 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1680363874
transform 1 0 4660 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4097
timestamp 1680363874
transform 1 0 4628 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3670
timestamp 1680363874
transform 1 0 4636 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4098
timestamp 1680363874
transform 1 0 4644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1680363874
transform 1 0 4660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1680363874
transform 1 0 4628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1680363874
transform 1 0 4636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1680363874
transform 1 0 4652 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1680363874
transform 1 0 4628 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1680363874
transform 1 0 4652 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1680363874
transform 1 0 4684 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1680363874
transform 1 0 4716 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1680363874
transform 1 0 4868 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4100
timestamp 1680363874
transform 1 0 4764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1680363874
transform 1 0 4804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1680363874
transform 1 0 4868 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1680363874
transform 1 0 4788 0 1 2805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_38
timestamp 1680363874
transform 1 0 48 0 1 2770
box -10 -3 10 3
use FILL  FILL_4137
timestamp 1680363874
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1680363874
transform 1 0 80 0 1 2770
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1680363874
transform 1 0 88 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_40
timestamp 1680363874
transform -1 0 120 0 1 2770
box -8 -3 32 105
use FILL  FILL_4142
timestamp 1680363874
transform 1 0 120 0 1 2770
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1680363874
transform 1 0 128 0 1 2770
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1680363874
transform 1 0 136 0 1 2770
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1680363874
transform 1 0 144 0 1 2770
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1680363874
transform 1 0 152 0 1 2770
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1680363874
transform 1 0 160 0 1 2770
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1680363874
transform 1 0 168 0 1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1680363874
transform 1 0 176 0 1 2770
box -7 -3 39 105
use FILL  FILL_4154
timestamp 1680363874
transform 1 0 208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1680363874
transform 1 0 216 0 1 2770
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1680363874
transform 1 0 224 0 1 2770
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1680363874
transform 1 0 232 0 1 2770
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1680363874
transform 1 0 240 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_217
timestamp 1680363874
transform 1 0 248 0 1 2770
box -8 -3 46 105
use FILL  FILL_4165
timestamp 1680363874
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1680363874
transform 1 0 296 0 1 2770
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1680363874
transform 1 0 304 0 1 2770
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1680363874
transform 1 0 312 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_288
timestamp 1680363874
transform -1 0 336 0 1 2770
box -9 -3 26 105
use FILL  FILL_4177
timestamp 1680363874
transform 1 0 336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1680363874
transform 1 0 344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1680363874
transform 1 0 352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1680363874
transform 1 0 360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1680363874
transform 1 0 368 0 1 2770
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1680363874
transform 1 0 376 0 1 2770
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1680363874
transform 1 0 384 0 1 2770
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1680363874
transform 1 0 392 0 1 2770
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1680363874
transform 1 0 400 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3759
timestamp 1680363874
transform 1 0 444 0 1 2775
box -3 -3 3 3
use AOI21X1  AOI21X1_2
timestamp 1680363874
transform -1 0 440 0 1 2770
box -7 -3 39 105
use FILL  FILL_4186
timestamp 1680363874
transform 1 0 440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1680363874
transform 1 0 448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1680363874
transform 1 0 456 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3760
timestamp 1680363874
transform 1 0 476 0 1 2775
box -3 -3 3 3
use FILL  FILL_4189
timestamp 1680363874
transform 1 0 464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1680363874
transform 1 0 472 0 1 2770
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1680363874
transform 1 0 480 0 1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1680363874
transform -1 0 520 0 1 2770
box -7 -3 39 105
use FILL  FILL_4192
timestamp 1680363874
transform 1 0 520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1680363874
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1680363874
transform 1 0 536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1680363874
transform 1 0 544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1680363874
transform 1 0 552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1680363874
transform 1 0 560 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1680363874
transform -1 0 600 0 1 2770
box -8 -3 40 105
use FILL  FILL_4198
timestamp 1680363874
transform 1 0 600 0 1 2770
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1680363874
transform 1 0 608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1680363874
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1680363874
transform 1 0 624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1680363874
transform 1 0 632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1680363874
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1680363874
transform 1 0 648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1680363874
transform 1 0 656 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_42
timestamp 1680363874
transform 1 0 664 0 1 2770
box -8 -3 32 105
use FILL  FILL_4206
timestamp 1680363874
transform 1 0 688 0 1 2770
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1680363874
transform 1 0 696 0 1 2770
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1680363874
transform 1 0 704 0 1 2770
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1680363874
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1680363874
transform 1 0 720 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_289
timestamp 1680363874
transform -1 0 744 0 1 2770
box -9 -3 26 105
use FILL  FILL_4211
timestamp 1680363874
transform 1 0 744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1680363874
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1680363874
transform 1 0 760 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_290
timestamp 1680363874
transform -1 0 784 0 1 2770
box -9 -3 26 105
use FILL  FILL_4225
timestamp 1680363874
transform 1 0 784 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_145
timestamp 1680363874
transform 1 0 792 0 1 2770
box -8 -3 46 105
use FILL  FILL_4226
timestamp 1680363874
transform 1 0 832 0 1 2770
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1680363874
transform 1 0 840 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_291
timestamp 1680363874
transform -1 0 864 0 1 2770
box -9 -3 26 105
use FILL  FILL_4228
timestamp 1680363874
transform 1 0 864 0 1 2770
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1680363874
transform 1 0 872 0 1 2770
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1680363874
transform 1 0 880 0 1 2770
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1680363874
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1680363874
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1680363874
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1680363874
transform 1 0 912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1680363874
transform 1 0 920 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_146
timestamp 1680363874
transform 1 0 928 0 1 2770
box -8 -3 46 105
use FILL  FILL_4236
timestamp 1680363874
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1680363874
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1680363874
transform -1 0 1104 0 1 2770
box -5 -3 126 105
use XOR2X1  XOR2X1_0
timestamp 1680363874
transform 1 0 1104 0 1 2770
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1680363874
transform 1 0 1160 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_292
timestamp 1680363874
transform 1 0 1256 0 1 2770
box -9 -3 26 105
use FILL  FILL_4238
timestamp 1680363874
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1680363874
transform 1 0 1280 0 1 2770
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1680363874
transform 1 0 1288 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_218
timestamp 1680363874
transform 1 0 1296 0 1 2770
box -8 -3 46 105
use FILL  FILL_4272
timestamp 1680363874
transform 1 0 1336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1680363874
transform 1 0 1344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1680363874
transform 1 0 1352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1680363874
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1680363874
transform 1 0 1368 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_219
timestamp 1680363874
transform 1 0 1376 0 1 2770
box -8 -3 46 105
use FILL  FILL_4277
timestamp 1680363874
transform 1 0 1416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1680363874
transform 1 0 1424 0 1 2770
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1680363874
transform 1 0 1432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1680363874
transform 1 0 1440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1680363874
transform 1 0 1448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1680363874
transform 1 0 1456 0 1 2770
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1680363874
transform 1 0 1464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1680363874
transform 1 0 1472 0 1 2770
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1680363874
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1680363874
transform 1 0 1488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1680363874
transform 1 0 1496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1680363874
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1680363874
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3761
timestamp 1680363874
transform 1 0 1532 0 1 2775
box -3 -3 3 3
use FILL  FILL_4300
timestamp 1680363874
transform 1 0 1520 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_272
timestamp 1680363874
transform 1 0 1528 0 1 2770
box -8 -3 104 105
use FILL  FILL_4302
timestamp 1680363874
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1680363874
transform 1 0 1632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1680363874
transform 1 0 1640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1680363874
transform 1 0 1648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1680363874
transform 1 0 1656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1680363874
transform 1 0 1664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1680363874
transform 1 0 1672 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_221
timestamp 1680363874
transform 1 0 1680 0 1 2770
box -8 -3 46 105
use FILL  FILL_4309
timestamp 1680363874
transform 1 0 1720 0 1 2770
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1680363874
transform 1 0 1728 0 1 2770
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1680363874
transform 1 0 1736 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_294
timestamp 1680363874
transform -1 0 1760 0 1 2770
box -9 -3 26 105
use FILL  FILL_4325
timestamp 1680363874
transform 1 0 1760 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1680363874
transform -1 0 1864 0 1 2770
box -8 -3 104 105
use OAI22X1  OAI22X1_222
timestamp 1680363874
transform -1 0 1904 0 1 2770
box -8 -3 46 105
use INVX2  INVX2_295
timestamp 1680363874
transform -1 0 1920 0 1 2770
box -9 -3 26 105
use FILL  FILL_4326
timestamp 1680363874
transform 1 0 1920 0 1 2770
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1680363874
transform 1 0 1928 0 1 2770
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1680363874
transform 1 0 1936 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3762
timestamp 1680363874
transform 1 0 1964 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_224
timestamp 1680363874
transform -1 0 1984 0 1 2770
box -8 -3 46 105
use FILL  FILL_4345
timestamp 1680363874
transform 1 0 1984 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_298
timestamp 1680363874
transform -1 0 2008 0 1 2770
box -9 -3 26 105
use FILL  FILL_4346
timestamp 1680363874
transform 1 0 2008 0 1 2770
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1680363874
transform 1 0 2016 0 1 2770
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1680363874
transform 1 0 2024 0 1 2770
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1680363874
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_30
timestamp 1680363874
transform -1 0 2064 0 1 2770
box -5 -3 28 105
use FILL  FILL_4356
timestamp 1680363874
transform 1 0 2064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1680363874
transform 1 0 2072 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_31
timestamp 1680363874
transform -1 0 2104 0 1 2770
box -5 -3 28 105
use FILL  FILL_4358
timestamp 1680363874
transform 1 0 2104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1680363874
transform 1 0 2112 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_32
timestamp 1680363874
transform -1 0 2144 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1680363874
transform -1 0 2168 0 1 2770
box -5 -3 28 105
use FILL  FILL_4360
timestamp 1680363874
transform 1 0 2168 0 1 2770
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1680363874
transform 1 0 2176 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_34
timestamp 1680363874
transform -1 0 2208 0 1 2770
box -5 -3 28 105
use FILL  FILL_4362
timestamp 1680363874
transform 1 0 2208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1680363874
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_35
timestamp 1680363874
transform -1 0 2248 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1680363874
transform 1 0 2248 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1680363874
transform 1 0 2272 0 1 2770
box -5 -3 28 105
use FILL  FILL_4370
timestamp 1680363874
transform 1 0 2296 0 1 2770
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1680363874
transform 1 0 2304 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_38
timestamp 1680363874
transform 1 0 2312 0 1 2770
box -5 -3 28 105
use FILL  FILL_4372
timestamp 1680363874
transform 1 0 2336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1680363874
transform 1 0 2344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1680363874
transform 1 0 2352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1680363874
transform 1 0 2360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1680363874
transform 1 0 2368 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_302
timestamp 1680363874
transform -1 0 2392 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1680363874
transform 1 0 2392 0 1 2770
box -9 -3 26 105
use FILL  FILL_4389
timestamp 1680363874
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1680363874
transform 1 0 2416 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_226
timestamp 1680363874
transform 1 0 2424 0 1 2770
box -8 -3 46 105
use FILL  FILL_4393
timestamp 1680363874
transform 1 0 2464 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_305
timestamp 1680363874
transform -1 0 2488 0 1 2770
box -9 -3 26 105
use FILL  FILL_4394
timestamp 1680363874
transform 1 0 2488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1680363874
transform 1 0 2496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1680363874
transform 1 0 2504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1680363874
transform 1 0 2512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1680363874
transform 1 0 2520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1680363874
transform 1 0 2528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1680363874
transform 1 0 2536 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1680363874
transform -1 0 2640 0 1 2770
box -8 -3 104 105
use FILL  FILL_4410
timestamp 1680363874
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1680363874
transform 1 0 2648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1680363874
transform 1 0 2656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1680363874
transform 1 0 2664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1680363874
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_229
timestamp 1680363874
transform 1 0 2680 0 1 2770
box -8 -3 46 105
use FILL  FILL_4424
timestamp 1680363874
transform 1 0 2720 0 1 2770
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1680363874
transform 1 0 2728 0 1 2770
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1680363874
transform 1 0 2736 0 1 2770
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1680363874
transform 1 0 2744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1680363874
transform 1 0 2752 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_308
timestamp 1680363874
transform -1 0 2776 0 1 2770
box -9 -3 26 105
use FILL  FILL_4429
timestamp 1680363874
transform 1 0 2776 0 1 2770
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1680363874
transform 1 0 2784 0 1 2770
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1680363874
transform 1 0 2792 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3763
timestamp 1680363874
transform 1 0 2812 0 1 2775
box -3 -3 3 3
use FILL  FILL_4435
timestamp 1680363874
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3764
timestamp 1680363874
transform 1 0 2852 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_230
timestamp 1680363874
transform 1 0 2808 0 1 2770
box -8 -3 46 105
use FILL  FILL_4437
timestamp 1680363874
transform 1 0 2848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1680363874
transform 1 0 2856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1680363874
transform 1 0 2864 0 1 2770
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1680363874
transform 1 0 2872 0 1 2770
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1680363874
transform 1 0 2880 0 1 2770
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1680363874
transform 1 0 2888 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_112
timestamp 1680363874
transform 1 0 2896 0 1 2770
box -8 -3 34 105
use FILL  FILL_4449
timestamp 1680363874
transform 1 0 2928 0 1 2770
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1680363874
transform 1 0 2936 0 1 2770
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1680363874
transform 1 0 2944 0 1 2770
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1680363874
transform 1 0 2952 0 1 2770
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1680363874
transform 1 0 2960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1680363874
transform 1 0 2968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1680363874
transform 1 0 2976 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1680363874
transform 1 0 2984 0 1 2770
box -8 -3 34 105
use FILL  FILL_4464
timestamp 1680363874
transform 1 0 3016 0 1 2770
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1680363874
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1680363874
transform 1 0 3032 0 1 2770
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1680363874
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_309
timestamp 1680363874
transform -1 0 3064 0 1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_278
timestamp 1680363874
transform -1 0 3160 0 1 2770
box -8 -3 104 105
use FILL  FILL_4471
timestamp 1680363874
transform 1 0 3160 0 1 2770
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1680363874
transform 1 0 3168 0 1 2770
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1680363874
transform 1 0 3176 0 1 2770
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1680363874
transform 1 0 3184 0 1 2770
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1680363874
transform 1 0 3192 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3765
timestamp 1680363874
transform 1 0 3236 0 1 2775
box -3 -3 3 3
use OAI21X1  OAI21X1_116
timestamp 1680363874
transform -1 0 3232 0 1 2770
box -8 -3 34 105
use FILL  FILL_4476
timestamp 1680363874
transform 1 0 3232 0 1 2770
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1680363874
transform 1 0 3240 0 1 2770
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1680363874
transform 1 0 3248 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3766
timestamp 1680363874
transform 1 0 3268 0 1 2775
box -3 -3 3 3
use FILL  FILL_4479
timestamp 1680363874
transform 1 0 3256 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3767
timestamp 1680363874
transform 1 0 3356 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_279
timestamp 1680363874
transform -1 0 3360 0 1 2770
box -8 -3 104 105
use FILL  FILL_4480
timestamp 1680363874
transform 1 0 3360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1680363874
transform 1 0 3368 0 1 2770
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1680363874
transform 1 0 3376 0 1 2770
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1680363874
transform 1 0 3384 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3768
timestamp 1680363874
transform 1 0 3404 0 1 2775
box -3 -3 3 3
use FILL  FILL_4514
timestamp 1680363874
transform 1 0 3392 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_117
timestamp 1680363874
transform -1 0 3432 0 1 2770
box -8 -3 34 105
use FILL  FILL_4515
timestamp 1680363874
transform 1 0 3432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1680363874
transform 1 0 3440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1680363874
transform 1 0 3448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1680363874
transform 1 0 3456 0 1 2770
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1680363874
transform 1 0 3464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1680363874
transform 1 0 3472 0 1 2770
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1680363874
transform 1 0 3480 0 1 2770
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1680363874
transform 1 0 3488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1680363874
transform 1 0 3496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1680363874
transform 1 0 3504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1680363874
transform 1 0 3512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1680363874
transform 1 0 3520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1680363874
transform 1 0 3528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1680363874
transform 1 0 3536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1680363874
transform 1 0 3544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1680363874
transform 1 0 3552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1680363874
transform 1 0 3560 0 1 2770
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1680363874
transform 1 0 3568 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_311
timestamp 1680363874
transform 1 0 3576 0 1 2770
box -9 -3 26 105
use FILL  FILL_4551
timestamp 1680363874
transform 1 0 3592 0 1 2770
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1680363874
transform 1 0 3600 0 1 2770
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1680363874
transform 1 0 3608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1680363874
transform 1 0 3616 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3769
timestamp 1680363874
transform 1 0 3636 0 1 2775
box -3 -3 3 3
use FILL  FILL_4559
timestamp 1680363874
transform 1 0 3624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1680363874
transform 1 0 3632 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_118
timestamp 1680363874
transform -1 0 3672 0 1 2770
box -8 -3 34 105
use FILL  FILL_4561
timestamp 1680363874
transform 1 0 3672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1680363874
transform 1 0 3680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1680363874
transform 1 0 3688 0 1 2770
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1680363874
transform 1 0 3696 0 1 2770
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1680363874
transform 1 0 3704 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_43
timestamp 1680363874
transform -1 0 3736 0 1 2770
box -8 -3 32 105
use FILL  FILL_4570
timestamp 1680363874
transform 1 0 3736 0 1 2770
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1680363874
transform 1 0 3744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1680363874
transform 1 0 3752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1680363874
transform 1 0 3760 0 1 2770
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1680363874
transform 1 0 3768 0 1 2770
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1680363874
transform 1 0 3776 0 1 2770
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1680363874
transform 1 0 3784 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_150
timestamp 1680363874
transform 1 0 3792 0 1 2770
box -8 -3 46 105
use FILL  FILL_4579
timestamp 1680363874
transform 1 0 3832 0 1 2770
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1680363874
transform 1 0 3840 0 1 2770
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1680363874
transform 1 0 3848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1680363874
transform 1 0 3856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1680363874
transform 1 0 3864 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_312
timestamp 1680363874
transform 1 0 3872 0 1 2770
box -9 -3 26 105
use FILL  FILL_4590
timestamp 1680363874
transform 1 0 3888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1680363874
transform 1 0 3896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1680363874
transform 1 0 3904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1680363874
transform 1 0 3912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1680363874
transform 1 0 3920 0 1 2770
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1680363874
transform 1 0 3928 0 1 2770
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1680363874
transform 1 0 3936 0 1 2770
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1680363874
transform 1 0 3944 0 1 2770
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1680363874
transform 1 0 3952 0 1 2770
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1680363874
transform 1 0 3960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1680363874
transform 1 0 3968 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_151
timestamp 1680363874
transform 1 0 3976 0 1 2770
box -8 -3 46 105
use FILL  FILL_4601
timestamp 1680363874
transform 1 0 4016 0 1 2770
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1680363874
transform 1 0 4024 0 1 2770
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1680363874
transform 1 0 4032 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_313
timestamp 1680363874
transform 1 0 4040 0 1 2770
box -9 -3 26 105
use FILL  FILL_4604
timestamp 1680363874
transform 1 0 4056 0 1 2770
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1680363874
transform 1 0 4064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1680363874
transform 1 0 4072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1680363874
transform 1 0 4080 0 1 2770
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1680363874
transform 1 0 4088 0 1 2770
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1680363874
transform 1 0 4096 0 1 2770
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1680363874
transform 1 0 4104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1680363874
transform 1 0 4112 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_152
timestamp 1680363874
transform 1 0 4120 0 1 2770
box -8 -3 46 105
use FILL  FILL_4618
timestamp 1680363874
transform 1 0 4160 0 1 2770
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1680363874
transform 1 0 4168 0 1 2770
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1680363874
transform 1 0 4176 0 1 2770
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1680363874
transform 1 0 4184 0 1 2770
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1680363874
transform 1 0 4192 0 1 2770
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1680363874
transform 1 0 4200 0 1 2770
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1680363874
transform 1 0 4208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1680363874
transform 1 0 4216 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_154
timestamp 1680363874
transform 1 0 4224 0 1 2770
box -8 -3 46 105
use FILL  FILL_4629
timestamp 1680363874
transform 1 0 4264 0 1 2770
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1680363874
transform 1 0 4272 0 1 2770
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1680363874
transform 1 0 4280 0 1 2770
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1680363874
transform 1 0 4288 0 1 2770
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1680363874
transform 1 0 4296 0 1 2770
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1680363874
transform 1 0 4304 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_45
timestamp 1680363874
transform -1 0 4336 0 1 2770
box -8 -3 32 105
use FILL  FILL_4638
timestamp 1680363874
transform 1 0 4336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1680363874
transform 1 0 4344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1680363874
transform 1 0 4352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1680363874
transform 1 0 4360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1680363874
transform 1 0 4368 0 1 2770
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1680363874
transform 1 0 4376 0 1 2770
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1680363874
transform 1 0 4384 0 1 2770
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1680363874
transform 1 0 4392 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3770
timestamp 1680363874
transform 1 0 4444 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_155
timestamp 1680363874
transform -1 0 4440 0 1 2770
box -8 -3 46 105
use FILL  FILL_4646
timestamp 1680363874
transform 1 0 4440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1680363874
transform 1 0 4448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1680363874
transform 1 0 4456 0 1 2770
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1680363874
transform 1 0 4464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1680363874
transform 1 0 4472 0 1 2770
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1680363874
transform 1 0 4480 0 1 2770
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1680363874
transform 1 0 4488 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_317
timestamp 1680363874
transform 1 0 4496 0 1 2770
box -9 -3 26 105
use FILL  FILL_4659
timestamp 1680363874
transform 1 0 4512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1680363874
transform 1 0 4520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1680363874
transform 1 0 4528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1680363874
transform 1 0 4536 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_231
timestamp 1680363874
transform 1 0 4544 0 1 2770
box -8 -3 46 105
use FILL  FILL_4663
timestamp 1680363874
transform 1 0 4584 0 1 2770
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1680363874
transform 1 0 4592 0 1 2770
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1680363874
transform 1 0 4600 0 1 2770
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1680363874
transform 1 0 4608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1680363874
transform 1 0 4616 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_156
timestamp 1680363874
transform 1 0 4624 0 1 2770
box -8 -3 46 105
use FILL  FILL_4671
timestamp 1680363874
transform 1 0 4664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1680363874
transform 1 0 4672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1680363874
transform 1 0 4680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1680363874
transform 1 0 4688 0 1 2770
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1680363874
transform 1 0 4696 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3771
timestamp 1680363874
transform 1 0 4756 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1680363874
transform 1 0 4780 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_287
timestamp 1680363874
transform -1 0 4800 0 1 2770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_39
timestamp 1680363874
transform 1 0 4827 0 1 2770
box -10 -3 10 3
use M3_M2  M3_M2_3805
timestamp 1680363874
transform 1 0 92 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4229
timestamp 1680363874
transform 1 0 92 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3806
timestamp 1680363874
transform 1 0 132 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4383
timestamp 1680363874
transform 1 0 140 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1680363874
transform 1 0 156 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1680363874
transform 1 0 172 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1680363874
transform 1 0 172 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3905
timestamp 1680363874
transform 1 0 188 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4230
timestamp 1680363874
transform 1 0 236 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3807
timestamp 1680363874
transform 1 0 340 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4219
timestamp 1680363874
transform 1 0 348 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3808
timestamp 1680363874
transform 1 0 372 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1680363874
transform 1 0 332 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4231
timestamp 1680363874
transform 1 0 340 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3931
timestamp 1680363874
transform 1 0 324 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4298
timestamp 1680363874
transform 1 0 332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1680363874
transform 1 0 476 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1680363874
transform 1 0 452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1680363874
transform 1 0 460 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3856
timestamp 1680363874
transform 1 0 412 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4299
timestamp 1680363874
transform 1 0 436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1680363874
transform 1 0 444 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3857
timestamp 1680363874
transform 1 0 452 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1680363874
transform 1 0 524 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1680363874
transform 1 0 532 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4301
timestamp 1680363874
transform 1 0 564 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1680363874
transform 1 0 572 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3876
timestamp 1680363874
transform 1 0 436 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1680363874
transform 1 0 460 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1680363874
transform 1 0 564 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1680363874
transform 1 0 364 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1680363874
transform 1 0 356 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4392
timestamp 1680363874
transform 1 0 460 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3907
timestamp 1680363874
transform 1 0 540 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1680363874
transform 1 0 572 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1680363874
transform 1 0 548 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1680363874
transform 1 0 588 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4234
timestamp 1680363874
transform 1 0 596 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1680363874
transform 1 0 604 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3879
timestamp 1680363874
transform 1 0 604 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1680363874
transform 1 0 596 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4221
timestamp 1680363874
transform 1 0 620 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3810
timestamp 1680363874
transform 1 0 644 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1680363874
transform 1 0 668 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4303
timestamp 1680363874
transform 1 0 708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1680363874
transform 1 0 716 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3880
timestamp 1680363874
transform 1 0 708 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1680363874
transform 1 0 628 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1680363874
transform 1 0 692 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1680363874
transform 1 0 756 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4236
timestamp 1680363874
transform 1 0 740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1680363874
transform 1 0 732 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3835
timestamp 1680363874
transform 1 0 748 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1680363874
transform 1 0 740 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4305
timestamp 1680363874
transform 1 0 764 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3910
timestamp 1680363874
transform 1 0 756 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4306
timestamp 1680363874
transform 1 0 788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1680363874
transform 1 0 804 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3881
timestamp 1680363874
transform 1 0 804 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4393
timestamp 1680363874
transform 1 0 780 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3911
timestamp 1680363874
transform 1 0 796 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1680363874
transform 1 0 820 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1680363874
transform 1 0 820 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1680363874
transform 1 0 860 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4386
timestamp 1680363874
transform 1 0 812 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1680363874
transform 1 0 828 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3811
timestamp 1680363874
transform 1 0 836 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4223
timestamp 1680363874
transform 1 0 940 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1680363874
transform 1 0 932 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3859
timestamp 1680363874
transform 1 0 892 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4307
timestamp 1680363874
transform 1 0 916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1680363874
transform 1 0 924 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3912
timestamp 1680363874
transform 1 0 884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1680363874
transform 1 0 940 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4387
timestamp 1680363874
transform 1 0 940 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3775
timestamp 1680363874
transform 1 0 956 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1680363874
transform 1 0 956 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1680363874
transform 1 0 964 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4309
timestamp 1680363874
transform 1 0 980 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3861
timestamp 1680363874
transform 1 0 988 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4388
timestamp 1680363874
transform 1 0 980 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3862
timestamp 1680363874
transform 1 0 1028 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4394
timestamp 1680363874
transform 1 0 1060 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1680363874
transform 1 0 1116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1680363874
transform 1 0 1156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3792
timestamp 1680363874
transform 1 0 1204 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1680363874
transform 1 0 1180 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1680363874
transform 1 0 1220 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4239
timestamp 1680363874
transform 1 0 1180 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3837
timestamp 1680363874
transform 1 0 1228 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4312
timestamp 1680363874
transform 1 0 1228 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3913
timestamp 1680363874
transform 1 0 1260 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1680363874
transform 1 0 1188 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1680363874
transform 1 0 1276 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1680363874
transform 1 0 1308 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1680363874
transform 1 0 1324 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4240
timestamp 1680363874
transform 1 0 1316 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3935
timestamp 1680363874
transform 1 0 1316 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4241
timestamp 1680363874
transform 1 0 1340 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3838
timestamp 1680363874
transform 1 0 1348 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1680363874
transform 1 0 1380 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1680363874
transform 1 0 1380 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4224
timestamp 1680363874
transform 1 0 1388 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1680363874
transform 1 0 1356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1680363874
transform 1 0 1372 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1680363874
transform 1 0 1340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1680363874
transform 1 0 1348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1680363874
transform 1 0 1364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3864
timestamp 1680363874
transform 1 0 1372 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1680363874
transform 1 0 1340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1680363874
transform 1 0 1356 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1680363874
transform 1 0 1348 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1680363874
transform 1 0 1348 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1680363874
transform 1 0 1396 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4225
timestamp 1680363874
transform 1 0 1412 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3777
timestamp 1680363874
transform 1 0 1484 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1680363874
transform 1 0 1428 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1680363874
transform 1 0 1500 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4244
timestamp 1680363874
transform 1 0 1428 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3840
timestamp 1680363874
transform 1 0 1452 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4316
timestamp 1680363874
transform 1 0 1452 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1680363874
transform 1 0 1508 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3884
timestamp 1680363874
transform 1 0 1508 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1680363874
transform 1 0 1580 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1680363874
transform 1 0 1652 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4245
timestamp 1680363874
transform 1 0 1636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1680363874
transform 1 0 1684 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3955
timestamp 1680363874
transform 1 0 1676 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4319
timestamp 1680363874
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1680363874
transform 1 0 1772 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3778
timestamp 1680363874
transform 1 0 1812 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4247
timestamp 1680363874
transform 1 0 1804 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3841
timestamp 1680363874
transform 1 0 1828 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1680363874
transform 1 0 1852 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1680363874
transform 1 0 1884 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4248
timestamp 1680363874
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1680363874
transform 1 0 1844 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3842
timestamp 1680363874
transform 1 0 1860 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4249
timestamp 1680363874
transform 1 0 1868 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1680363874
transform 1 0 1884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1680363874
transform 1 0 1860 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1680363874
transform 1 0 1876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1680363874
transform 1 0 1884 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3886
timestamp 1680363874
transform 1 0 1860 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1680363874
transform 1 0 1860 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1680363874
transform 1 0 1876 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4251
timestamp 1680363874
transform 1 0 1924 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3887
timestamp 1680363874
transform 1 0 1924 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4324
timestamp 1680363874
transform 1 0 1948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1680363874
transform 1 0 1964 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3888
timestamp 1680363874
transform 1 0 1964 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1680363874
transform 1 0 1956 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1680363874
transform 1 0 1972 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1680363874
transform 1 0 2012 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1680363874
transform 1 0 2004 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1680363874
transform 1 0 2044 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4252
timestamp 1680363874
transform 1 0 2044 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1680363874
transform 1 0 2052 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1680363874
transform 1 0 2068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1680363874
transform 1 0 2036 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3890
timestamp 1680363874
transform 1 0 2044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1680363874
transform 1 0 2036 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1680363874
transform 1 0 2044 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1680363874
transform 1 0 2076 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1680363874
transform 1 0 2092 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4215
timestamp 1680363874
transform 1 0 2092 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1680363874
transform 1 0 2060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1680363874
transform 1 0 2076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1680363874
transform 1 0 2084 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3891
timestamp 1680363874
transform 1 0 2084 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1680363874
transform 1 0 2060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1680363874
transform 1 0 2076 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1680363874
transform 1 0 2060 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1680363874
transform 1 0 2116 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1680363874
transform 1 0 2116 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1680363874
transform 1 0 2132 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4255
timestamp 1680363874
transform 1 0 2180 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1680363874
transform 1 0 2132 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3959
timestamp 1680363874
transform 1 0 2108 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1680363874
transform 1 0 2124 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1680363874
transform 1 0 2156 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1680363874
transform 1 0 2228 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4256
timestamp 1680363874
transform 1 0 2228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1680363874
transform 1 0 2252 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3962
timestamp 1680363874
transform 1 0 2252 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1680363874
transform 1 0 2292 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4257
timestamp 1680363874
transform 1 0 2284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1680363874
transform 1 0 2268 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3845
timestamp 1680363874
transform 1 0 2292 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4258
timestamp 1680363874
transform 1 0 2308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1680363874
transform 1 0 2292 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3892
timestamp 1680363874
transform 1 0 2276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1680363874
transform 1 0 2316 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4259
timestamp 1680363874
transform 1 0 2324 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3893
timestamp 1680363874
transform 1 0 2332 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1680363874
transform 1 0 2356 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4334
timestamp 1680363874
transform 1 0 2356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1680363874
transform 1 0 2380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1680363874
transform 1 0 2412 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3894
timestamp 1680363874
transform 1 0 2412 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4261
timestamp 1680363874
transform 1 0 2420 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3782
timestamp 1680363874
transform 1 0 2436 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4262
timestamp 1680363874
transform 1 0 2452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1680363874
transform 1 0 2468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1680363874
transform 1 0 2444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1680363874
transform 1 0 2460 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3895
timestamp 1680363874
transform 1 0 2460 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1680363874
transform 1 0 2436 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1680363874
transform 1 0 2468 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4264
timestamp 1680363874
transform 1 0 2492 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3920
timestamp 1680363874
transform 1 0 2516 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4265
timestamp 1680363874
transform 1 0 2540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1680363874
transform 1 0 2556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1680363874
transform 1 0 2580 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3865
timestamp 1680363874
transform 1 0 2580 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1680363874
transform 1 0 2596 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1680363874
transform 1 0 2596 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1680363874
transform 1 0 2612 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4267
timestamp 1680363874
transform 1 0 2612 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3866
timestamp 1680363874
transform 1 0 2612 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1680363874
transform 1 0 2628 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4268
timestamp 1680363874
transform 1 0 2636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1680363874
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1680363874
transform 1 0 2620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1680363874
transform 1 0 2628 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1680363874
transform 1 0 2644 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3896
timestamp 1680363874
transform 1 0 2644 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1680363874
transform 1 0 2620 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1680363874
transform 1 0 2668 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1680363874
transform 1 0 2764 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4270
timestamp 1680363874
transform 1 0 2692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1680363874
transform 1 0 2716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1680363874
transform 1 0 2772 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3942
timestamp 1680363874
transform 1 0 2708 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1680363874
transform 1 0 2780 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4344
timestamp 1680363874
transform 1 0 2820 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3921
timestamp 1680363874
transform 1 0 2812 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1680363874
transform 1 0 2812 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1680363874
transform 1 0 2844 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4345
timestamp 1680363874
transform 1 0 2844 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3922
timestamp 1680363874
transform 1 0 2844 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4271
timestamp 1680363874
transform 1 0 2876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1680363874
transform 1 0 2884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1680363874
transform 1 0 2868 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3898
timestamp 1680363874
transform 1 0 2884 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1680363874
transform 1 0 2876 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1680363874
transform 1 0 2916 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4273
timestamp 1680363874
transform 1 0 2916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1680363874
transform 1 0 2900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1680363874
transform 1 0 2916 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1680363874
transform 1 0 2932 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3867
timestamp 1680363874
transform 1 0 2932 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4348
timestamp 1680363874
transform 1 0 2988 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3849
timestamp 1680363874
transform 1 0 3020 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4390
timestamp 1680363874
transform 1 0 3012 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1680363874
transform 1 0 3092 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3945
timestamp 1680363874
transform 1 0 3092 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4349
timestamp 1680363874
transform 1 0 3100 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3868
timestamp 1680363874
transform 1 0 3140 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1680363874
transform 1 0 3164 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4276
timestamp 1680363874
transform 1 0 3244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1680363874
transform 1 0 3156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1680363874
transform 1 0 3164 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3899
timestamp 1680363874
transform 1 0 3156 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1680363874
transform 1 0 3172 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4352
timestamp 1680363874
transform 1 0 3204 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3900
timestamp 1680363874
transform 1 0 3204 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1680363874
transform 1 0 3164 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1680363874
transform 1 0 3212 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1680363874
transform 1 0 3156 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1680363874
transform 1 0 3172 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1680363874
transform 1 0 3260 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1680363874
transform 1 0 3260 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1680363874
transform 1 0 3388 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4216
timestamp 1680363874
transform 1 0 3404 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1680363874
transform 1 0 3428 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1680363874
transform 1 0 3436 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1680363874
transform 1 0 3492 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1680363874
transform 1 0 3508 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3901
timestamp 1680363874
transform 1 0 3492 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4278
timestamp 1680363874
transform 1 0 3556 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3965
timestamp 1680363874
transform 1 0 3548 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4355
timestamp 1680363874
transform 1 0 3572 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3925
timestamp 1680363874
transform 1 0 3572 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1680363874
transform 1 0 3604 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1680363874
transform 1 0 3596 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1680363874
transform 1 0 3612 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1680363874
transform 1 0 3604 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1680363874
transform 1 0 3628 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4279
timestamp 1680363874
transform 1 0 3620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1680363874
transform 1 0 3636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1680363874
transform 1 0 3612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1680363874
transform 1 0 3628 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1680363874
transform 1 0 3644 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3948
timestamp 1680363874
transform 1 0 3612 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1680363874
transform 1 0 3644 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1680363874
transform 1 0 3668 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1680363874
transform 1 0 3684 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1680363874
transform 1 0 3732 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4281
timestamp 1680363874
transform 1 0 3772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1680363874
transform 1 0 3724 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3871
timestamp 1680363874
transform 1 0 3772 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1680363874
transform 1 0 3788 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4360
timestamp 1680363874
transform 1 0 3788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1680363874
transform 1 0 3804 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3786
timestamp 1680363874
transform 1 0 3828 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4226
timestamp 1680363874
transform 1 0 3844 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1680363874
transform 1 0 3860 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3872
timestamp 1680363874
transform 1 0 3860 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1680363874
transform 1 0 3860 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1680363874
transform 1 0 3892 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4284
timestamp 1680363874
transform 1 0 3892 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3852
timestamp 1680363874
transform 1 0 3924 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4361
timestamp 1680363874
transform 1 0 3876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1680363874
transform 1 0 3916 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3873
timestamp 1680363874
transform 1 0 3924 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1680363874
transform 1 0 3876 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1680363874
transform 1 0 3916 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1680363874
transform 1 0 3980 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4363
timestamp 1680363874
transform 1 0 3980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1680363874
transform 1 0 4028 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1680363874
transform 1 0 4060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1680363874
transform 1 0 4108 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1680363874
transform 1 0 4164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1680363874
transform 1 0 4140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1680363874
transform 1 0 4156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3874
timestamp 1680363874
transform 1 0 4164 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4227
timestamp 1680363874
transform 1 0 4180 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3966
timestamp 1680363874
transform 1 0 4172 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1680363874
transform 1 0 4204 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1680363874
transform 1 0 4244 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1680363874
transform 1 0 4196 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4287
timestamp 1680363874
transform 1 0 4196 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3875
timestamp 1680363874
transform 1 0 4196 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4368
timestamp 1680363874
transform 1 0 4244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1680363874
transform 1 0 4276 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3903
timestamp 1680363874
transform 1 0 4244 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1680363874
transform 1 0 4292 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4288
timestamp 1680363874
transform 1 0 4292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1680363874
transform 1 0 4292 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3904
timestamp 1680363874
transform 1 0 4292 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1680363874
transform 1 0 4356 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1680363874
transform 1 0 4388 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4289
timestamp 1680363874
transform 1 0 4412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1680363874
transform 1 0 4428 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1680363874
transform 1 0 4332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1680363874
transform 1 0 4380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1680363874
transform 1 0 4428 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3967
timestamp 1680363874
transform 1 0 4316 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1680363874
transform 1 0 4380 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1680363874
transform 1 0 4428 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4374
timestamp 1680363874
transform 1 0 4444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1680363874
transform 1 0 4508 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1680363874
transform 1 0 4500 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3829
timestamp 1680363874
transform 1 0 4524 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4292
timestamp 1680363874
transform 1 0 4524 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1680363874
transform 1 0 4612 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3854
timestamp 1680363874
transform 1 0 4620 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4375
timestamp 1680363874
transform 1 0 4556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1680363874
transform 1 0 4604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1680363874
transform 1 0 4612 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3949
timestamp 1680363874
transform 1 0 4588 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1680363874
transform 1 0 4612 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1680363874
transform 1 0 4644 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4294
timestamp 1680363874
transform 1 0 4636 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3855
timestamp 1680363874
transform 1 0 4644 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4378
timestamp 1680363874
transform 1 0 4660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1680363874
transform 1 0 4692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1680363874
transform 1 0 4700 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1680363874
transform 1 0 4684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1680363874
transform 1 0 4708 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3831
timestamp 1680363874
transform 1 0 4756 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4297
timestamp 1680363874
transform 1 0 4756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1680363874
transform 1 0 4756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1680363874
transform 1 0 4764 0 1 2725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_40
timestamp 1680363874
transform 1 0 24 0 1 2670
box -10 -3 10 3
use FILL  FILL_4138
timestamp 1680363874
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1680363874
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_287
timestamp 1680363874
transform 1 0 88 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4143
timestamp 1680363874
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1680363874
transform 1 0 112 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3968
timestamp 1680363874
transform 1 0 132 0 1 2675
box -3 -3 3 3
use FILL  FILL_4145
timestamp 1680363874
transform 1 0 120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1680363874
transform 1 0 128 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1680363874
transform 1 0 136 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4153
timestamp 1680363874
transform 1 0 168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1680363874
transform 1 0 176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1680363874
transform 1 0 184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1680363874
transform 1 0 192 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_41
timestamp 1680363874
transform 1 0 200 0 -1 2770
box -8 -3 32 105
use FILL  FILL_4160
timestamp 1680363874
transform 1 0 224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1680363874
transform 1 0 232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1680363874
transform 1 0 240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1680363874
transform 1 0 248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1680363874
transform 1 0 256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1680363874
transform 1 0 264 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3969
timestamp 1680363874
transform 1 0 284 0 1 2675
box -3 -3 3 3
use FILL  FILL_4169
timestamp 1680363874
transform 1 0 272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1680363874
transform 1 0 280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1680363874
transform 1 0 288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1680363874
transform 1 0 296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1680363874
transform 1 0 304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1680363874
transform 1 0 312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1680363874
transform 1 0 320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1680363874
transform 1 0 328 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_2
timestamp 1680363874
transform -1 0 456 0 -1 2770
box -5 -3 126 105
use FILL  FILL_4215
timestamp 1680363874
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_3
timestamp 1680363874
transform -1 0 584 0 -1 2770
box -5 -3 126 105
use FILL  FILL_4216
timestamp 1680363874
transform 1 0 584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1680363874
transform 1 0 592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1680363874
transform 1 0 600 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_4
timestamp 1680363874
transform -1 0 728 0 -1 2770
box -5 -3 126 105
use FILL  FILL_4219
timestamp 1680363874
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1680363874
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1680363874
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1680363874
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1680363874
transform 1 0 760 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1680363874
transform -1 0 800 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4240
timestamp 1680363874
transform 1 0 800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1680363874
transform 1 0 808 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_6
timestamp 1680363874
transform -1 0 936 0 -1 2770
box -5 -3 126 105
use FILL  FILL_4242
timestamp 1680363874
transform 1 0 936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1680363874
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1680363874
transform 1 0 952 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1680363874
transform -1 0 992 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4245
timestamp 1680363874
transform 1 0 992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1680363874
transform 1 0 1000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1680363874
transform 1 0 1008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1680363874
transform 1 0 1016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1680363874
transform 1 0 1024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1680363874
transform 1 0 1032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1680363874
transform 1 0 1040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1680363874
transform 1 0 1048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1680363874
transform 1 0 1056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1680363874
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1680363874
transform 1 0 1072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1680363874
transform 1 0 1080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1680363874
transform 1 0 1088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1680363874
transform 1 0 1096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1680363874
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1680363874
transform 1 0 1112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1680363874
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1680363874
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1680363874
transform 1 0 1136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1680363874
transform 1 0 1144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1680363874
transform 1 0 1152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1680363874
transform 1 0 1160 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_270
timestamp 1680363874
transform 1 0 1168 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4267
timestamp 1680363874
transform 1 0 1264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1680363874
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1680363874
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_293
timestamp 1680363874
transform 1 0 1288 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4290
timestamp 1680363874
transform 1 0 1304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1680363874
transform 1 0 1312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1680363874
transform 1 0 1320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1680363874
transform 1 0 1328 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_220
timestamp 1680363874
transform 1 0 1336 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4294
timestamp 1680363874
transform 1 0 1376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1680363874
transform 1 0 1384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1680363874
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1680363874
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1680363874
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_271
timestamp 1680363874
transform 1 0 1416 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4299
timestamp 1680363874
transform 1 0 1512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1680363874
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1680363874
transform 1 0 1528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1680363874
transform 1 0 1536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1680363874
transform 1 0 1544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1680363874
transform 1 0 1552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1680363874
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1680363874
transform 1 0 1568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1680363874
transform 1 0 1576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1680363874
transform 1 0 1584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1680363874
transform 1 0 1592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1680363874
transform 1 0 1600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1680363874
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1680363874
transform 1 0 1616 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3970
timestamp 1680363874
transform 1 0 1644 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_273
timestamp 1680363874
transform 1 0 1624 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4322
timestamp 1680363874
transform 1 0 1720 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3971
timestamp 1680363874
transform 1 0 1740 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_296
timestamp 1680363874
transform 1 0 1728 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4327
timestamp 1680363874
transform 1 0 1744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1680363874
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1680363874
transform 1 0 1760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1680363874
transform 1 0 1768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1680363874
transform 1 0 1776 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_297
timestamp 1680363874
transform 1 0 1784 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4332
timestamp 1680363874
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1680363874
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1680363874
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1680363874
transform 1 0 1824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1680363874
transform 1 0 1832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1680363874
transform 1 0 1840 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_223
timestamp 1680363874
transform -1 0 1888 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4338
timestamp 1680363874
transform 1 0 1888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1680363874
transform 1 0 1896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1680363874
transform 1 0 1904 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3972
timestamp 1680363874
transform 1 0 1924 0 1 2675
box -3 -3 3 3
use FILL  FILL_4341
timestamp 1680363874
transform 1 0 1912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1680363874
transform 1 0 1920 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_147
timestamp 1680363874
transform 1 0 1928 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4347
timestamp 1680363874
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1680363874
transform 1 0 1976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1680363874
transform 1 0 1984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1680363874
transform 1 0 1992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1680363874
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1680363874
transform 1 0 2008 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3973
timestamp 1680363874
transform 1 0 2028 0 1 2675
box -3 -3 3 3
use FILL  FILL_4363
timestamp 1680363874
transform 1 0 2016 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_299
timestamp 1680363874
transform -1 0 2040 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4364
timestamp 1680363874
transform 1 0 2040 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_225
timestamp 1680363874
transform -1 0 2088 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4365
timestamp 1680363874
transform 1 0 2088 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1680363874
transform -1 0 2192 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4366
timestamp 1680363874
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1680363874
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1680363874
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1680363874
transform 1 0 2216 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_300
timestamp 1680363874
transform 1 0 2224 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4376
timestamp 1680363874
transform 1 0 2240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1680363874
transform 1 0 2248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1680363874
transform 1 0 2256 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_39
timestamp 1680363874
transform 1 0 2264 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_40
timestamp 1680363874
transform 1 0 2288 0 -1 2770
box -5 -3 28 105
use FILL  FILL_4379
timestamp 1680363874
transform 1 0 2312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1680363874
transform 1 0 2320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1680363874
transform 1 0 2328 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_301
timestamp 1680363874
transform 1 0 2336 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4382
timestamp 1680363874
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1680363874
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1680363874
transform 1 0 2368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1680363874
transform 1 0 2376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1680363874
transform 1 0 2384 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_304
timestamp 1680363874
transform 1 0 2392 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4390
timestamp 1680363874
transform 1 0 2408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1680363874
transform 1 0 2416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1680363874
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_227
timestamp 1680363874
transform 1 0 2432 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4396
timestamp 1680363874
transform 1 0 2472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1680363874
transform 1 0 2480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1680363874
transform 1 0 2488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1680363874
transform 1 0 2496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1680363874
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1680363874
transform 1 0 2512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1680363874
transform 1 0 2520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1680363874
transform 1 0 2528 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_306
timestamp 1680363874
transform 1 0 2536 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4413
timestamp 1680363874
transform 1 0 2552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1680363874
transform 1 0 2560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1680363874
transform 1 0 2568 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_307
timestamp 1680363874
transform 1 0 2576 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4416
timestamp 1680363874
transform 1 0 2592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1680363874
transform 1 0 2600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1680363874
transform 1 0 2608 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_228
timestamp 1680363874
transform 1 0 2616 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4419
timestamp 1680363874
transform 1 0 2656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1680363874
transform 1 0 2664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1680363874
transform 1 0 2672 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_277
timestamp 1680363874
transform 1 0 2680 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4430
timestamp 1680363874
transform 1 0 2776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1680363874
transform 1 0 2784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1680363874
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1680363874
transform 1 0 2800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1680363874
transform 1 0 2808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1680363874
transform 1 0 2816 0 -1 2770
box -8 -3 16 105
use AND2X2  AND2X2_17
timestamp 1680363874
transform -1 0 2856 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4441
timestamp 1680363874
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1680363874
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1680363874
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1680363874
transform 1 0 2880 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_113
timestamp 1680363874
transform 1 0 2888 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4450
timestamp 1680363874
transform 1 0 2920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1680363874
transform 1 0 2928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1680363874
transform 1 0 2936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1680363874
transform 1 0 2944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1680363874
transform 1 0 2952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1680363874
transform 1 0 2960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1680363874
transform 1 0 2968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1680363874
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_115
timestamp 1680363874
transform 1 0 2984 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4465
timestamp 1680363874
transform 1 0 3016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1680363874
transform 1 0 3024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1680363874
transform 1 0 3032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1680363874
transform 1 0 3040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1680363874
transform 1 0 3048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1680363874
transform 1 0 3056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1680363874
transform 1 0 3064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1680363874
transform 1 0 3072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1680363874
transform 1 0 3080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1680363874
transform 1 0 3088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1680363874
transform 1 0 3096 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_310
timestamp 1680363874
transform 1 0 3104 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4489
timestamp 1680363874
transform 1 0 3120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1680363874
transform 1 0 3128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1680363874
transform 1 0 3136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1680363874
transform 1 0 3144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1680363874
transform 1 0 3152 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3974
timestamp 1680363874
transform 1 0 3228 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_280
timestamp 1680363874
transform -1 0 3256 0 -1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3975
timestamp 1680363874
transform 1 0 3268 0 1 2675
box -3 -3 3 3
use FILL  FILL_4494
timestamp 1680363874
transform 1 0 3256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1680363874
transform 1 0 3264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1680363874
transform 1 0 3272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1680363874
transform 1 0 3280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1680363874
transform 1 0 3288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1680363874
transform 1 0 3296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1680363874
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1680363874
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1680363874
transform 1 0 3320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1680363874
transform 1 0 3328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1680363874
transform 1 0 3336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1680363874
transform 1 0 3344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1680363874
transform 1 0 3352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1680363874
transform 1 0 3360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1680363874
transform 1 0 3368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1680363874
transform 1 0 3376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1680363874
transform 1 0 3384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1680363874
transform 1 0 3392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1680363874
transform 1 0 3400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1680363874
transform 1 0 3408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1680363874
transform 1 0 3416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1680363874
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1680363874
transform 1 0 3432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1680363874
transform 1 0 3440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1680363874
transform 1 0 3448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1680363874
transform 1 0 3456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1680363874
transform 1 0 3464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1680363874
transform 1 0 3472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1680363874
transform 1 0 3480 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_148
timestamp 1680363874
transform -1 0 3528 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4540
timestamp 1680363874
transform 1 0 3528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1680363874
transform 1 0 3536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1680363874
transform 1 0 3544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1680363874
transform 1 0 3552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1680363874
transform 1 0 3560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1680363874
transform 1 0 3568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1680363874
transform 1 0 3576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1680363874
transform 1 0 3584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1680363874
transform 1 0 3592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1680363874
transform 1 0 3600 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_149
timestamp 1680363874
transform 1 0 3608 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4562
timestamp 1680363874
transform 1 0 3648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1680363874
transform 1 0 3656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1680363874
transform 1 0 3664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1680363874
transform 1 0 3672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1680363874
transform 1 0 3680 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1680363874
transform -1 0 3784 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4578
timestamp 1680363874
transform 1 0 3784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1680363874
transform 1 0 3792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1680363874
transform 1 0 3800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1680363874
transform 1 0 3808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1680363874
transform 1 0 3816 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_44
timestamp 1680363874
transform -1 0 3848 0 -1 2770
box -8 -3 32 105
use FILL  FILL_4586
timestamp 1680363874
transform 1 0 3848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1680363874
transform 1 0 3856 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_314
timestamp 1680363874
transform 1 0 3864 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_282
timestamp 1680363874
transform 1 0 3880 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4612
timestamp 1680363874
transform 1 0 3976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1680363874
transform 1 0 3984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1680363874
transform 1 0 3992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1680363874
transform 1 0 4000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1680363874
transform 1 0 4008 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1680363874
transform 1 0 4016 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4617
timestamp 1680363874
transform 1 0 4112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1680363874
transform 1 0 4120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1680363874
transform 1 0 4128 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_153
timestamp 1680363874
transform -1 0 4176 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4623
timestamp 1680363874
transform 1 0 4176 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_284
timestamp 1680363874
transform 1 0 4184 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4632
timestamp 1680363874
transform 1 0 4280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1680363874
transform 1 0 4288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1680363874
transform 1 0 4296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1680363874
transform 1 0 4304 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_315
timestamp 1680363874
transform 1 0 4312 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_285
timestamp 1680363874
transform -1 0 4424 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_316
timestamp 1680363874
transform 1 0 4424 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4648
timestamp 1680363874
transform 1 0 4440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1680363874
transform 1 0 4448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1680363874
transform 1 0 4456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1680363874
transform 1 0 4464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1680363874
transform 1 0 4472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1680363874
transform 1 0 4480 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_46
timestamp 1680363874
transform -1 0 4512 0 -1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_286
timestamp 1680363874
transform 1 0 4512 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4668
timestamp 1680363874
transform 1 0 4608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1680363874
transform 1 0 4616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1680363874
transform 1 0 4624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1680363874
transform 1 0 4632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1680363874
transform 1 0 4640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1680363874
transform 1 0 4648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1680363874
transform 1 0 4656 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_157
timestamp 1680363874
transform 1 0 4664 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4681
timestamp 1680363874
transform 1 0 4704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1680363874
transform 1 0 4712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1680363874
transform 1 0 4720 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_318
timestamp 1680363874
transform 1 0 4728 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4684
timestamp 1680363874
transform 1 0 4744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1680363874
transform 1 0 4752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1680363874
transform 1 0 4760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1680363874
transform 1 0 4768 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_319
timestamp 1680363874
transform 1 0 4776 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4688
timestamp 1680363874
transform 1 0 4792 0 -1 2770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_41
timestamp 1680363874
transform 1 0 4851 0 1 2670
box -10 -3 10 3
use M2_M1  M2_M1_4512
timestamp 1680363874
transform 1 0 84 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4113
timestamp 1680363874
transform 1 0 92 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4414
timestamp 1680363874
transform 1 0 100 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4059
timestamp 1680363874
transform 1 0 100 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4582
timestamp 1680363874
transform 1 0 140 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1680363874
transform 1 0 204 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1680363874
transform 1 0 196 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4080
timestamp 1680363874
transform 1 0 220 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1680363874
transform 1 0 308 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1680363874
transform 1 0 236 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1680363874
transform 1 0 308 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4416
timestamp 1680363874
transform 1 0 332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1680363874
transform 1 0 340 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4060
timestamp 1680363874
transform 1 0 244 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1680363874
transform 1 0 316 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4583
timestamp 1680363874
transform 1 0 244 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4114
timestamp 1680363874
transform 1 0 300 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1680363874
transform 1 0 340 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4395
timestamp 1680363874
transform 1 0 356 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1680363874
transform 1 0 372 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4062
timestamp 1680363874
transform 1 0 380 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4513
timestamp 1680363874
transform 1 0 396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1680363874
transform 1 0 380 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4081
timestamp 1680363874
transform 1 0 388 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4396
timestamp 1680363874
transform 1 0 412 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_4063
timestamp 1680363874
transform 1 0 412 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1680363874
transform 1 0 436 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1680363874
transform 1 0 460 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4397
timestamp 1680363874
transform 1 0 452 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1680363874
transform 1 0 444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1680363874
transform 1 0 492 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1680363874
transform 1 0 476 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4064
timestamp 1680363874
transform 1 0 484 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4585
timestamp 1680363874
transform 1 0 484 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4116
timestamp 1680363874
transform 1 0 476 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1680363874
transform 1 0 492 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4420
timestamp 1680363874
transform 1 0 508 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4117
timestamp 1680363874
transform 1 0 516 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4515
timestamp 1680363874
transform 1 0 540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1680363874
transform 1 0 564 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4013
timestamp 1680363874
transform 1 0 596 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1680363874
transform 1 0 588 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1680363874
transform 1 0 612 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1680363874
transform 1 0 612 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4398
timestamp 1680363874
transform 1 0 620 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3991
timestamp 1680363874
transform 1 0 636 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4404
timestamp 1680363874
transform 1 0 612 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1680363874
transform 1 0 628 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1680363874
transform 1 0 612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1680363874
transform 1 0 636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1680363874
transform 1 0 636 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4118
timestamp 1680363874
transform 1 0 636 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1680363874
transform 1 0 700 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1680363874
transform 1 0 716 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4424
timestamp 1680363874
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1680363874
transform 1 0 716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1680363874
transform 1 0 692 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1680363874
transform 1 0 708 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4066
timestamp 1680363874
transform 1 0 716 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4426
timestamp 1680363874
transform 1 0 764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1680363874
transform 1 0 772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1680363874
transform 1 0 764 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4040
timestamp 1680363874
transform 1 0 788 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1680363874
transform 1 0 804 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4519
timestamp 1680363874
transform 1 0 788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1680363874
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4083
timestamp 1680363874
transform 1 0 796 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1680363874
transform 1 0 836 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4428
timestamp 1680363874
transform 1 0 820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1680363874
transform 1 0 828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1680363874
transform 1 0 844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1680363874
transform 1 0 860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1680363874
transform 1 0 868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1680363874
transform 1 0 884 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1680363874
transform 1 0 916 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3993
timestamp 1680363874
transform 1 0 932 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4399
timestamp 1680363874
transform 1 0 932 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_4006
timestamp 1680363874
transform 1 0 956 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4407
timestamp 1680363874
transform 1 0 948 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1680363874
transform 1 0 940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1680363874
transform 1 0 956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1680363874
transform 1 0 956 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4084
timestamp 1680363874
transform 1 0 956 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1680363874
transform 1 0 980 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1680363874
transform 1 0 1020 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1680363874
transform 1 0 1036 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4435
timestamp 1680363874
transform 1 0 988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1680363874
transform 1 0 1004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1680363874
transform 1 0 1020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1680363874
transform 1 0 1028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1680363874
transform 1 0 996 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1680363874
transform 1 0 1012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1680363874
transform 1 0 1068 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_4016
timestamp 1680363874
transform 1 0 1108 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4525
timestamp 1680363874
transform 1 0 1116 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4085
timestamp 1680363874
transform 1 0 1132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1680363874
transform 1 0 1196 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4526
timestamp 1680363874
transform 1 0 1196 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4086
timestamp 1680363874
transform 1 0 1244 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4439
timestamp 1680363874
transform 1 0 1260 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3995
timestamp 1680363874
transform 1 0 1284 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1680363874
transform 1 0 1292 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4440
timestamp 1680363874
transform 1 0 1292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1680363874
transform 1 0 1268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1680363874
transform 1 0 1284 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4067
timestamp 1680363874
transform 1 0 1292 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4529
timestamp 1680363874
transform 1 0 1308 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4018
timestamp 1680363874
transform 1 0 1340 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1680363874
transform 1 0 1332 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1680363874
transform 1 0 1348 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4441
timestamp 1680363874
transform 1 0 1388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1680363874
transform 1 0 1364 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4068
timestamp 1680363874
transform 1 0 1388 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1680363874
transform 1 0 1364 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1680363874
transform 1 0 1380 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1680363874
transform 1 0 1468 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4442
timestamp 1680363874
transform 1 0 1468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1680363874
transform 1 0 1476 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4069
timestamp 1680363874
transform 1 0 1484 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1680363874
transform 1 0 1596 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4444
timestamp 1680363874
transform 1 0 1548 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4070
timestamp 1680363874
transform 1 0 1548 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4531
timestamp 1680363874
transform 1 0 1596 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4121
timestamp 1680363874
transform 1 0 1604 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1680363874
transform 1 0 1636 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1680363874
transform 1 0 1636 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4400
timestamp 1680363874
transform 1 0 1636 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1680363874
transform 1 0 1628 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_4043
timestamp 1680363874
transform 1 0 1628 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4410
timestamp 1680363874
transform 1 0 1652 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_4020
timestamp 1680363874
transform 1 0 1716 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4411
timestamp 1680363874
transform 1 0 1724 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1680363874
transform 1 0 1716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1680363874
transform 1 0 1748 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1680363874
transform 1 0 1764 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_4008
timestamp 1680363874
transform 1 0 1772 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1680363874
transform 1 0 1788 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4446
timestamp 1680363874
transform 1 0 1772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1680363874
transform 1 0 1788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1680363874
transform 1 0 1796 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4089
timestamp 1680363874
transform 1 0 1804 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1680363874
transform 1 0 1852 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1680363874
transform 1 0 1844 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1680363874
transform 1 0 1884 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4448
timestamp 1680363874
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1680363874
transform 1 0 1852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1680363874
transform 1 0 1868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1680363874
transform 1 0 1884 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4071
timestamp 1680363874
transform 1 0 1852 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4534
timestamp 1680363874
transform 1 0 1860 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4072
timestamp 1680363874
transform 1 0 1884 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1680363874
transform 1 0 1900 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4535
timestamp 1680363874
transform 1 0 1908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1680363874
transform 1 0 1916 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4090
timestamp 1680363874
transform 1 0 1916 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4452
timestamp 1680363874
transform 1 0 1940 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3984
timestamp 1680363874
transform 1 0 1964 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4453
timestamp 1680363874
transform 1 0 2028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1680363874
transform 1 0 2044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1680363874
transform 1 0 2036 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4073
timestamp 1680363874
transform 1 0 2044 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4538
timestamp 1680363874
transform 1 0 2068 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3985
timestamp 1680363874
transform 1 0 2196 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4455
timestamp 1680363874
transform 1 0 2108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1680363874
transform 1 0 2164 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4044
timestamp 1680363874
transform 1 0 2180 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4457
timestamp 1680363874
transform 1 0 2204 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4045
timestamp 1680363874
transform 1 0 2228 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4458
timestamp 1680363874
transform 1 0 2260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1680363874
transform 1 0 2084 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4074
timestamp 1680363874
transform 1 0 2108 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1680363874
transform 1 0 2164 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4540
timestamp 1680363874
transform 1 0 2180 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4076
timestamp 1680363874
transform 1 0 2204 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1680363874
transform 1 0 2180 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1680363874
transform 1 0 2220 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1680363874
transform 1 0 2284 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1680363874
transform 1 0 2308 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1680363874
transform 1 0 2300 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1680363874
transform 1 0 2316 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1680363874
transform 1 0 2348 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4459
timestamp 1680363874
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1680363874
transform 1 0 2380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1680363874
transform 1 0 2300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1680363874
transform 1 0 2396 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3977
timestamp 1680363874
transform 1 0 2420 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1680363874
transform 1 0 2452 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4461
timestamp 1680363874
transform 1 0 2444 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4046
timestamp 1680363874
transform 1 0 2460 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4543
timestamp 1680363874
transform 1 0 2460 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4122
timestamp 1680363874
transform 1 0 2468 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4544
timestamp 1680363874
transform 1 0 2508 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4093
timestamp 1680363874
transform 1 0 2508 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1680363874
transform 1 0 2636 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4462
timestamp 1680363874
transform 1 0 2572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1680363874
transform 1 0 2612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1680363874
transform 1 0 2620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1680363874
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1680363874
transform 1 0 2524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1680363874
transform 1 0 2612 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1680363874
transform 1 0 2628 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4094
timestamp 1680363874
transform 1 0 2572 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4548
timestamp 1680363874
transform 1 0 2652 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4095
timestamp 1680363874
transform 1 0 2628 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1680363874
transform 1 0 2644 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1680363874
transform 1 0 2612 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1680363874
transform 1 0 2700 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4466
timestamp 1680363874
transform 1 0 2700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1680363874
transform 1 0 2676 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4097
timestamp 1680363874
transform 1 0 2740 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1680363874
transform 1 0 2796 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4467
timestamp 1680363874
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4047
timestamp 1680363874
transform 1 0 2788 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4550
timestamp 1680363874
transform 1 0 2788 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4048
timestamp 1680363874
transform 1 0 2916 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4468
timestamp 1680363874
transform 1 0 2972 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1680363874
transform 1 0 2988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1680363874
transform 1 0 3012 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_4049
timestamp 1680363874
transform 1 0 3012 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4470
timestamp 1680363874
transform 1 0 3028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1680363874
transform 1 0 3076 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4098
timestamp 1680363874
transform 1 0 3076 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4471
timestamp 1680363874
transform 1 0 3100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1680363874
transform 1 0 3092 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1680363874
transform 1 0 3132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1680363874
transform 1 0 3140 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4029
timestamp 1680363874
transform 1 0 3156 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1680363874
transform 1 0 3180 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4413
timestamp 1680363874
transform 1 0 3172 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1680363874
transform 1 0 3156 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4050
timestamp 1680363874
transform 1 0 3172 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1680363874
transform 1 0 3156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1680363874
transform 1 0 3244 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1680363874
transform 1 0 3196 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1680363874
transform 1 0 3284 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4474
timestamp 1680363874
transform 1 0 3244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1680363874
transform 1 0 3276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1680363874
transform 1 0 3284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1680363874
transform 1 0 3180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1680363874
transform 1 0 3196 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4100
timestamp 1680363874
transform 1 0 3196 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1680363874
transform 1 0 3236 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1680363874
transform 1 0 3268 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4556
timestamp 1680363874
transform 1 0 3316 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4102
timestamp 1680363874
transform 1 0 3308 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1680363874
transform 1 0 3332 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1680363874
transform 1 0 3412 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4477
timestamp 1680363874
transform 1 0 3436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1680363874
transform 1 0 3492 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4052
timestamp 1680363874
transform 1 0 3508 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1680363874
transform 1 0 3524 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4479
timestamp 1680363874
transform 1 0 3532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1680363874
transform 1 0 3516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1680363874
transform 1 0 3524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1680363874
transform 1 0 3540 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4126
timestamp 1680363874
transform 1 0 3516 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4560
timestamp 1680363874
transform 1 0 3556 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4127
timestamp 1680363874
transform 1 0 3588 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4480
timestamp 1680363874
transform 1 0 3628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1680363874
transform 1 0 3660 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1680363874
transform 1 0 3716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1680363874
transform 1 0 3724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1680363874
transform 1 0 3764 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4000
timestamp 1680363874
transform 1 0 3788 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4483
timestamp 1680363874
transform 1 0 3804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1680363874
transform 1 0 3820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1680363874
transform 1 0 3796 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1680363874
transform 1 0 3812 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4103
timestamp 1680363874
transform 1 0 3812 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4485
timestamp 1680363874
transform 1 0 3852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1680363874
transform 1 0 3860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1680363874
transform 1 0 3876 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4032
timestamp 1680363874
transform 1 0 3900 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4563
timestamp 1680363874
transform 1 0 3892 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4033
timestamp 1680363874
transform 1 0 3932 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4488
timestamp 1680363874
transform 1 0 3924 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4054
timestamp 1680363874
transform 1 0 3932 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4489
timestamp 1680363874
transform 1 0 3948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1680363874
transform 1 0 3916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1680363874
transform 1 0 3932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1680363874
transform 1 0 3940 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4104
timestamp 1680363874
transform 1 0 3940 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1680363874
transform 1 0 3980 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1680363874
transform 1 0 4004 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4589
timestamp 1680363874
transform 1 0 4004 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1680363874
transform 1 0 4044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1680363874
transform 1 0 4060 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4105
timestamp 1680363874
transform 1 0 4092 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1680363874
transform 1 0 4100 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1680363874
transform 1 0 4132 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4492
timestamp 1680363874
transform 1 0 4116 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4057
timestamp 1680363874
transform 1 0 4124 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4493
timestamp 1680363874
transform 1 0 4132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1680363874
transform 1 0 4100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1680363874
transform 1 0 4108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1680363874
transform 1 0 4124 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4106
timestamp 1680363874
transform 1 0 4116 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4570
timestamp 1680363874
transform 1 0 4148 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4035
timestamp 1680363874
transform 1 0 4156 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1680363874
transform 1 0 4188 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4494
timestamp 1680363874
transform 1 0 4172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1680363874
transform 1 0 4188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1680363874
transform 1 0 4180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1680363874
transform 1 0 4204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1680363874
transform 1 0 4228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1680363874
transform 1 0 4236 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4107
timestamp 1680363874
transform 1 0 4236 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1680363874
transform 1 0 4292 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1680363874
transform 1 0 4284 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4498
timestamp 1680363874
transform 1 0 4292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1680363874
transform 1 0 4268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1680363874
transform 1 0 4284 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4108
timestamp 1680363874
transform 1 0 4284 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1680363874
transform 1 0 4324 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4499
timestamp 1680363874
transform 1 0 4332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1680363874
transform 1 0 4340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1680363874
transform 1 0 4356 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4078
timestamp 1680363874
transform 1 0 4348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1680363874
transform 1 0 4348 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1680363874
transform 1 0 4388 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1680363874
transform 1 0 4420 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4502
timestamp 1680363874
transform 1 0 4388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1680363874
transform 1 0 4404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1680363874
transform 1 0 4412 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4079
timestamp 1680363874
transform 1 0 4388 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4575
timestamp 1680363874
transform 1 0 4396 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4109
timestamp 1680363874
transform 1 0 4372 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1680363874
transform 1 0 4404 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1680363874
transform 1 0 4436 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4576
timestamp 1680363874
transform 1 0 4444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1680363874
transform 1 0 4452 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4111
timestamp 1680363874
transform 1 0 4444 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1680363874
transform 1 0 4484 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4590
timestamp 1680363874
transform 1 0 4492 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4129
timestamp 1680363874
transform 1 0 4476 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1680363874
transform 1 0 4516 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4505
timestamp 1680363874
transform 1 0 4556 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4011
timestamp 1680363874
transform 1 0 4580 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1680363874
transform 1 0 4588 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4506
timestamp 1680363874
transform 1 0 4580 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1680363874
transform 1 0 4588 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4037
timestamp 1680363874
transform 1 0 4612 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4507
timestamp 1680363874
transform 1 0 4612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1680363874
transform 1 0 4604 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1680363874
transform 1 0 4636 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1680363874
transform 1 0 4652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1680363874
transform 1 0 4676 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4012
timestamp 1680363874
transform 1 0 4708 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4510
timestamp 1680363874
transform 1 0 4700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1680363874
transform 1 0 4756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1680363874
transform 1 0 4780 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4131
timestamp 1680363874
transform 1 0 4780 0 1 2585
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_42
timestamp 1680363874
transform 1 0 48 0 1 2570
box -10 -3 10 3
use FILL  FILL_4689
timestamp 1680363874
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1680363874
transform 1 0 80 0 1 2570
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1680363874
transform 1 0 88 0 1 2570
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1680363874
transform 1 0 96 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1680363874
transform 1 0 104 0 1 2570
box -7 -3 39 105
use FILL  FILL_4696
timestamp 1680363874
transform 1 0 136 0 1 2570
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1680363874
transform 1 0 144 0 1 2570
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1680363874
transform 1 0 152 0 1 2570
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1680363874
transform 1 0 160 0 1 2570
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1680363874
transform 1 0 168 0 1 2570
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1680363874
transform 1 0 176 0 1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_35
timestamp 1680363874
transform 1 0 184 0 1 2570
box -8 -3 32 105
use FILL  FILL_4707
timestamp 1680363874
transform 1 0 208 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4132
timestamp 1680363874
transform 1 0 228 0 1 2575
box -3 -3 3 3
use FILL  FILL_4708
timestamp 1680363874
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1680363874
transform 1 0 224 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4133
timestamp 1680363874
transform 1 0 292 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1680363874
transform 1 0 348 0 1 2575
box -3 -3 3 3
use FAX1  FAX1_7
timestamp 1680363874
transform -1 0 352 0 1 2570
box -5 -3 126 105
use FILL  FILL_4710
timestamp 1680363874
transform 1 0 352 0 1 2570
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1680363874
transform 1 0 360 0 1 2570
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1680363874
transform 1 0 368 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_6
timestamp 1680363874
transform -1 0 408 0 1 2570
box -7 -3 39 105
use FILL  FILL_4719
timestamp 1680363874
transform 1 0 408 0 1 2570
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1680363874
transform 1 0 416 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4135
timestamp 1680363874
transform 1 0 436 0 1 2575
box -3 -3 3 3
use FILL  FILL_4721
timestamp 1680363874
transform 1 0 424 0 1 2570
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1680363874
transform 1 0 432 0 1 2570
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1680363874
transform 1 0 440 0 1 2570
box -8 -3 16 105
use AND2X1  AND2X1_0
timestamp 1680363874
transform -1 0 480 0 1 2570
box -8 -3 40 105
use FILL  FILL_4724
timestamp 1680363874
transform 1 0 480 0 1 2570
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1680363874
transform 1 0 488 0 1 2570
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1680363874
transform 1 0 496 0 1 2570
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1680363874
transform 1 0 504 0 1 2570
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1680363874
transform 1 0 512 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1680363874
transform -1 0 552 0 1 2570
box -7 -3 39 105
use FILL  FILL_4740
timestamp 1680363874
transform 1 0 552 0 1 2570
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1680363874
transform 1 0 560 0 1 2570
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1680363874
transform 1 0 568 0 1 2570
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1680363874
transform 1 0 576 0 1 2570
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1680363874
transform 1 0 584 0 1 2570
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1680363874
transform 1 0 592 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1680363874
transform 1 0 600 0 1 2570
box -8 -3 40 105
use FILL  FILL_4754
timestamp 1680363874
transform 1 0 632 0 1 2570
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1680363874
transform 1 0 640 0 1 2570
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1680363874
transform 1 0 648 0 1 2570
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1680363874
transform 1 0 656 0 1 2570
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1680363874
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1680363874
transform 1 0 672 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_160
timestamp 1680363874
transform -1 0 720 0 1 2570
box -8 -3 46 105
use FILL  FILL_4765
timestamp 1680363874
transform 1 0 720 0 1 2570
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1680363874
transform 1 0 728 0 1 2570
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1680363874
transform 1 0 736 0 1 2570
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1680363874
transform 1 0 744 0 1 2570
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1680363874
transform 1 0 752 0 1 2570
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1680363874
transform 1 0 760 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_9
timestamp 1680363874
transform -1 0 800 0 1 2570
box -7 -3 39 105
use FILL  FILL_4778
timestamp 1680363874
transform 1 0 800 0 1 2570
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1680363874
transform 1 0 808 0 1 2570
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1680363874
transform 1 0 816 0 1 2570
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1680363874
transform 1 0 824 0 1 2570
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1680363874
transform 1 0 832 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_161
timestamp 1680363874
transform -1 0 880 0 1 2570
box -8 -3 46 105
use FILL  FILL_4790
timestamp 1680363874
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1680363874
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1680363874
transform 1 0 896 0 1 2570
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1680363874
transform 1 0 904 0 1 2570
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1680363874
transform 1 0 912 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1680363874
transform -1 0 952 0 1 2570
box -8 -3 40 105
use FILL  FILL_4802
timestamp 1680363874
transform 1 0 952 0 1 2570
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1680363874
transform 1 0 960 0 1 2570
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1680363874
transform 1 0 968 0 1 2570
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1680363874
transform 1 0 976 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_162
timestamp 1680363874
transform -1 0 1024 0 1 2570
box -8 -3 46 105
use FILL  FILL_4809
timestamp 1680363874
transform 1 0 1024 0 1 2570
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1680363874
transform 1 0 1032 0 1 2570
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1680363874
transform 1 0 1040 0 1 2570
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1680363874
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1680363874
transform 1 0 1056 0 1 2570
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1680363874
transform 1 0 1064 0 1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_36
timestamp 1680363874
transform -1 0 1096 0 1 2570
box -8 -3 32 105
use FILL  FILL_4821
timestamp 1680363874
transform 1 0 1096 0 1 2570
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1680363874
transform 1 0 1104 0 1 2570
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1680363874
transform 1 0 1112 0 1 2570
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1680363874
transform 1 0 1120 0 1 2570
box -8 -3 16 105
use XOR2X1  XOR2X1_1
timestamp 1680363874
transform -1 0 1184 0 1 2570
box -8 -3 64 105
use FILL  FILL_4828
timestamp 1680363874
transform 1 0 1184 0 1 2570
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1680363874
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1680363874
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1680363874
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1680363874
transform 1 0 1216 0 1 2570
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1680363874
transform 1 0 1224 0 1 2570
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1680363874
transform 1 0 1232 0 1 2570
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1680363874
transform 1 0 1240 0 1 2570
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1680363874
transform 1 0 1248 0 1 2570
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1680363874
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4136
timestamp 1680363874
transform 1 0 1308 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_232
timestamp 1680363874
transform 1 0 1264 0 1 2570
box -8 -3 46 105
use FILL  FILL_4850
timestamp 1680363874
transform 1 0 1304 0 1 2570
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1680363874
transform 1 0 1312 0 1 2570
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1680363874
transform 1 0 1320 0 1 2570
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1680363874
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1680363874
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1680363874
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4137
timestamp 1680363874
transform 1 0 1420 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_288
timestamp 1680363874
transform 1 0 1352 0 1 2570
box -8 -3 104 105
use FILL  FILL_4862
timestamp 1680363874
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_322
timestamp 1680363874
transform 1 0 1456 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1680363874
transform -1 0 1488 0 1 2570
box -9 -3 26 105
use FILL  FILL_4871
timestamp 1680363874
transform 1 0 1488 0 1 2570
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1680363874
transform 1 0 1496 0 1 2570
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1680363874
transform 1 0 1504 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4138
timestamp 1680363874
transform 1 0 1572 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_289
timestamp 1680363874
transform -1 0 1608 0 1 2570
box -8 -3 104 105
use FILL  FILL_4874
timestamp 1680363874
transform 1 0 1608 0 1 2570
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1680363874
transform 1 0 1616 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1680363874
transform -1 0 1656 0 1 2570
box -8 -3 40 105
use FILL  FILL_4886
timestamp 1680363874
transform 1 0 1656 0 1 2570
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1680363874
transform 1 0 1664 0 1 2570
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1680363874
transform 1 0 1672 0 1 2570
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1680363874
transform 1 0 1680 0 1 2570
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1680363874
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1680363874
transform -1 0 1728 0 1 2570
box -8 -3 40 105
use FILL  FILL_4895
timestamp 1680363874
transform 1 0 1728 0 1 2570
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1680363874
transform 1 0 1736 0 1 2570
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1680363874
transform 1 0 1744 0 1 2570
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1680363874
transform 1 0 1752 0 1 2570
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1680363874
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_165
timestamp 1680363874
transform -1 0 1808 0 1 2570
box -8 -3 46 105
use FILL  FILL_4900
timestamp 1680363874
transform 1 0 1808 0 1 2570
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1680363874
transform 1 0 1816 0 1 2570
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1680363874
transform 1 0 1824 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4139
timestamp 1680363874
transform 1 0 1844 0 1 2575
box -3 -3 3 3
use FILL  FILL_4907
timestamp 1680363874
transform 1 0 1832 0 1 2570
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1680363874
transform 1 0 1840 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4140
timestamp 1680363874
transform 1 0 1860 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_166
timestamp 1680363874
transform -1 0 1888 0 1 2570
box -8 -3 46 105
use FILL  FILL_4910
timestamp 1680363874
transform 1 0 1888 0 1 2570
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1680363874
transform 1 0 1896 0 1 2570
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1680363874
transform 1 0 1904 0 1 2570
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1680363874
transform 1 0 1912 0 1 2570
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1680363874
transform 1 0 1920 0 1 2570
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1680363874
transform 1 0 1928 0 1 2570
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1680363874
transform 1 0 1936 0 1 2570
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1680363874
transform 1 0 1944 0 1 2570
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1680363874
transform 1 0 1952 0 1 2570
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1680363874
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1680363874
transform 1 0 1968 0 1 2570
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1680363874
transform 1 0 1976 0 1 2570
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1680363874
transform 1 0 1984 0 1 2570
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1680363874
transform 1 0 1992 0 1 2570
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1680363874
transform 1 0 2000 0 1 2570
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1680363874
transform 1 0 2008 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_237
timestamp 1680363874
transform -1 0 2056 0 1 2570
box -8 -3 46 105
use FILL  FILL_4941
timestamp 1680363874
transform 1 0 2056 0 1 2570
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1680363874
transform 1 0 2064 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_291
timestamp 1680363874
transform 1 0 2072 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1680363874
transform 1 0 2168 0 1 2570
box -8 -3 104 105
use FILL  FILL_4951
timestamp 1680363874
transform 1 0 2264 0 1 2570
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1680363874
transform 1 0 2272 0 1 2570
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1680363874
transform 1 0 2280 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_293
timestamp 1680363874
transform 1 0 2288 0 1 2570
box -8 -3 104 105
use FILL  FILL_4972
timestamp 1680363874
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_328
timestamp 1680363874
transform 1 0 2392 0 1 2570
box -9 -3 26 105
use FILL  FILL_4973
timestamp 1680363874
transform 1 0 2408 0 1 2570
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1680363874
transform 1 0 2416 0 1 2570
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1680363874
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1680363874
transform 1 0 2432 0 1 2570
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1680363874
transform 1 0 2440 0 1 2570
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1680363874
transform 1 0 2448 0 1 2570
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1680363874
transform 1 0 2456 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_329
timestamp 1680363874
transform -1 0 2480 0 1 2570
box -9 -3 26 105
use FILL  FILL_4987
timestamp 1680363874
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1680363874
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1680363874
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1680363874
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_295
timestamp 1680363874
transform 1 0 2512 0 1 2570
box -8 -3 104 105
use OAI22X1  OAI22X1_240
timestamp 1680363874
transform 1 0 2608 0 1 2570
box -8 -3 46 105
use FILL  FILL_4994
timestamp 1680363874
transform 1 0 2648 0 1 2570
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1680363874
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_297
timestamp 1680363874
transform 1 0 2664 0 1 2570
box -8 -3 104 105
use FILL  FILL_5000
timestamp 1680363874
transform 1 0 2760 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_332
timestamp 1680363874
transform 1 0 2768 0 1 2570
box -9 -3 26 105
use FILL  FILL_5002
timestamp 1680363874
transform 1 0 2784 0 1 2570
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1680363874
transform 1 0 2792 0 1 2570
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1680363874
transform 1 0 2800 0 1 2570
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1680363874
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1680363874
transform 1 0 2816 0 1 2570
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1680363874
transform 1 0 2824 0 1 2570
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1680363874
transform 1 0 2832 0 1 2570
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1680363874
transform 1 0 2840 0 1 2570
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1680363874
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1680363874
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1680363874
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1680363874
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1680363874
transform 1 0 2880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1680363874
transform 1 0 2888 0 1 2570
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1680363874
transform 1 0 2896 0 1 2570
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1680363874
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1680363874
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1680363874
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1680363874
transform 1 0 2928 0 1 2570
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1680363874
transform 1 0 2936 0 1 2570
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1680363874
transform 1 0 2944 0 1 2570
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1680363874
transform 1 0 2952 0 1 2570
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1680363874
transform 1 0 2960 0 1 2570
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1680363874
transform 1 0 2968 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_123
timestamp 1680363874
transform 1 0 2976 0 1 2570
box -8 -3 34 105
use FILL  FILL_5042
timestamp 1680363874
transform 1 0 3008 0 1 2570
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1680363874
transform 1 0 3016 0 1 2570
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1680363874
transform 1 0 3024 0 1 2570
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1680363874
transform 1 0 3032 0 1 2570
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1680363874
transform 1 0 3040 0 1 2570
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1680363874
transform 1 0 3048 0 1 2570
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1680363874
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1680363874
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1680363874
transform 1 0 3072 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_167
timestamp 1680363874
transform 1 0 3080 0 1 2570
box -8 -3 46 105
use FILL  FILL_5062
timestamp 1680363874
transform 1 0 3120 0 1 2570
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1680363874
transform 1 0 3128 0 1 2570
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1680363874
transform 1 0 3136 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_124
timestamp 1680363874
transform 1 0 3144 0 1 2570
box -8 -3 34 105
use FILL  FILL_5065
timestamp 1680363874
transform 1 0 3176 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1680363874
transform 1 0 3184 0 1 2570
box -8 -3 104 105
use FILL  FILL_5074
timestamp 1680363874
transform 1 0 3280 0 1 2570
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1680363874
transform 1 0 3288 0 1 2570
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1680363874
transform 1 0 3296 0 1 2570
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1680363874
transform 1 0 3304 0 1 2570
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1680363874
transform 1 0 3312 0 1 2570
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1680363874
transform 1 0 3320 0 1 2570
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1680363874
transform 1 0 3328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1680363874
transform 1 0 3336 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_335
timestamp 1680363874
transform 1 0 3344 0 1 2570
box -9 -3 26 105
use FILL  FILL_5093
timestamp 1680363874
transform 1 0 3360 0 1 2570
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1680363874
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1680363874
transform 1 0 3376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1680363874
transform 1 0 3384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1680363874
transform 1 0 3392 0 1 2570
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1680363874
transform 1 0 3400 0 1 2570
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1680363874
transform 1 0 3408 0 1 2570
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1680363874
transform 1 0 3416 0 1 2570
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1680363874
transform 1 0 3424 0 1 2570
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1680363874
transform 1 0 3432 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_336
timestamp 1680363874
transform -1 0 3456 0 1 2570
box -9 -3 26 105
use FILL  FILL_5109
timestamp 1680363874
transform 1 0 3456 0 1 2570
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1680363874
transform 1 0 3464 0 1 2570
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1680363874
transform 1 0 3472 0 1 2570
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1680363874
transform 1 0 3480 0 1 2570
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1680363874
transform 1 0 3488 0 1 2570
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1680363874
transform 1 0 3496 0 1 2570
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1680363874
transform 1 0 3504 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_170
timestamp 1680363874
transform -1 0 3552 0 1 2570
box -8 -3 46 105
use FILL  FILL_5118
timestamp 1680363874
transform 1 0 3552 0 1 2570
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1680363874
transform 1 0 3560 0 1 2570
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1680363874
transform 1 0 3568 0 1 2570
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1680363874
transform 1 0 3576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1680363874
transform 1 0 3584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1680363874
transform 1 0 3592 0 1 2570
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1680363874
transform 1 0 3600 0 1 2570
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1680363874
transform 1 0 3608 0 1 2570
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1680363874
transform 1 0 3616 0 1 2570
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1680363874
transform 1 0 3624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1680363874
transform 1 0 3632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1680363874
transform 1 0 3640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1680363874
transform 1 0 3648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1680363874
transform 1 0 3656 0 1 2570
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1680363874
transform 1 0 3664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1680363874
transform 1 0 3672 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_337
timestamp 1680363874
transform 1 0 3680 0 1 2570
box -9 -3 26 105
use FILL  FILL_5140
timestamp 1680363874
transform 1 0 3696 0 1 2570
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1680363874
transform 1 0 3704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1680363874
transform 1 0 3712 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_47
timestamp 1680363874
transform -1 0 3744 0 1 2570
box -8 -3 32 105
use FILL  FILL_5143
timestamp 1680363874
transform 1 0 3744 0 1 2570
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1680363874
transform 1 0 3752 0 1 2570
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1680363874
transform 1 0 3760 0 1 2570
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1680363874
transform 1 0 3768 0 1 2570
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1680363874
transform 1 0 3776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1680363874
transform 1 0 3784 0 1 2570
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1680363874
transform 1 0 3792 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4141
timestamp 1680363874
transform 1 0 3820 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_171
timestamp 1680363874
transform 1 0 3800 0 1 2570
box -8 -3 46 105
use FILL  FILL_5158
timestamp 1680363874
transform 1 0 3840 0 1 2570
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1680363874
transform 1 0 3848 0 1 2570
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1680363874
transform 1 0 3856 0 1 2570
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1680363874
transform 1 0 3864 0 1 2570
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1680363874
transform 1 0 3872 0 1 2570
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1680363874
transform 1 0 3880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1680363874
transform 1 0 3888 0 1 2570
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1680363874
transform 1 0 3896 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_173
timestamp 1680363874
transform 1 0 3904 0 1 2570
box -8 -3 46 105
use FILL  FILL_5175
timestamp 1680363874
transform 1 0 3944 0 1 2570
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1680363874
transform 1 0 3952 0 1 2570
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1680363874
transform 1 0 3960 0 1 2570
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1680363874
transform 1 0 3968 0 1 2570
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1680363874
transform 1 0 3976 0 1 2570
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1680363874
transform 1 0 3984 0 1 2570
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1680363874
transform 1 0 3992 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_48
timestamp 1680363874
transform 1 0 4000 0 1 2570
box -8 -3 32 105
use FILL  FILL_5189
timestamp 1680363874
transform 1 0 4024 0 1 2570
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1680363874
transform 1 0 4032 0 1 2570
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1680363874
transform 1 0 4040 0 1 2570
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1680363874
transform 1 0 4048 0 1 2570
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1680363874
transform 1 0 4056 0 1 2570
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1680363874
transform 1 0 4064 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_340
timestamp 1680363874
transform -1 0 4088 0 1 2570
box -9 -3 26 105
use FILL  FILL_5201
timestamp 1680363874
transform 1 0 4088 0 1 2570
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1680363874
transform 1 0 4096 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_241
timestamp 1680363874
transform 1 0 4104 0 1 2570
box -8 -3 46 105
use FILL  FILL_5207
timestamp 1680363874
transform 1 0 4144 0 1 2570
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1680363874
transform 1 0 4152 0 1 2570
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1680363874
transform 1 0 4160 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_176
timestamp 1680363874
transform -1 0 4208 0 1 2570
box -8 -3 46 105
use FILL  FILL_5213
timestamp 1680363874
transform 1 0 4208 0 1 2570
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1680363874
transform 1 0 4216 0 1 2570
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1680363874
transform 1 0 4224 0 1 2570
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1680363874
transform 1 0 4232 0 1 2570
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1680363874
transform 1 0 4240 0 1 2570
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1680363874
transform 1 0 4248 0 1 2570
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1680363874
transform 1 0 4256 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_242
timestamp 1680363874
transform 1 0 4264 0 1 2570
box -8 -3 46 105
use FILL  FILL_5230
timestamp 1680363874
transform 1 0 4304 0 1 2570
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1680363874
transform 1 0 4312 0 1 2570
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1680363874
transform 1 0 4320 0 1 2570
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1680363874
transform 1 0 4328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1680363874
transform 1 0 4336 0 1 2570
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1680363874
transform 1 0 4344 0 1 2570
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1680363874
transform 1 0 4352 0 1 2570
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1680363874
transform 1 0 4360 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_178
timestamp 1680363874
transform -1 0 4408 0 1 2570
box -8 -3 46 105
use FILL  FILL_5243
timestamp 1680363874
transform 1 0 4408 0 1 2570
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1680363874
transform 1 0 4416 0 1 2570
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1680363874
transform 1 0 4424 0 1 2570
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1680363874
transform 1 0 4432 0 1 2570
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1680363874
transform 1 0 4440 0 1 2570
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1680363874
transform 1 0 4448 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_50
timestamp 1680363874
transform -1 0 4480 0 1 2570
box -8 -3 32 105
use FILL  FILL_5249
timestamp 1680363874
transform 1 0 4480 0 1 2570
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1680363874
transform 1 0 4488 0 1 2570
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1680363874
transform 1 0 4496 0 1 2570
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1680363874
transform 1 0 4504 0 1 2570
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1680363874
transform 1 0 4512 0 1 2570
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1680363874
transform 1 0 4520 0 1 2570
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1680363874
transform 1 0 4528 0 1 2570
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1680363874
transform 1 0 4536 0 1 2570
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1680363874
transform 1 0 4544 0 1 2570
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1680363874
transform 1 0 4552 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_343
timestamp 1680363874
transform -1 0 4576 0 1 2570
box -9 -3 26 105
use FILL  FILL_5263
timestamp 1680363874
transform 1 0 4576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1680363874
transform 1 0 4584 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_179
timestamp 1680363874
transform -1 0 4632 0 1 2570
box -8 -3 46 105
use FILL  FILL_5265
timestamp 1680363874
transform 1 0 4632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1680363874
transform 1 0 4640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1680363874
transform 1 0 4648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1680363874
transform 1 0 4656 0 1 2570
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1680363874
transform 1 0 4664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1680363874
transform 1 0 4672 0 1 2570
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1680363874
transform 1 0 4680 0 1 2570
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1680363874
transform 1 0 4688 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_304
timestamp 1680363874
transform -1 0 4792 0 1 2570
box -8 -3 104 105
use FILL  FILL_5276
timestamp 1680363874
transform 1 0 4792 0 1 2570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_43
timestamp 1680363874
transform 1 0 4827 0 1 2570
box -10 -3 10 3
use M3_M2  M3_M2_4142
timestamp 1680363874
transform 1 0 76 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1680363874
transform 1 0 76 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4597
timestamp 1680363874
transform 1 0 84 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4231
timestamp 1680363874
transform 1 0 84 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1680363874
transform 1 0 84 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1680363874
transform 1 0 116 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1680363874
transform 1 0 100 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4680
timestamp 1680363874
transform 1 0 100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1680363874
transform 1 0 140 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1680363874
transform 1 0 156 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1680363874
transform 1 0 164 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4165
timestamp 1680363874
transform 1 0 196 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1680363874
transform 1 0 180 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4593
timestamp 1680363874
transform 1 0 188 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1680363874
transform 1 0 180 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4212
timestamp 1680363874
transform 1 0 188 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1680363874
transform 1 0 284 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4599
timestamp 1680363874
transform 1 0 292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1680363874
transform 1 0 276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1680363874
transform 1 0 284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1680363874
transform 1 0 300 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4181
timestamp 1680363874
transform 1 0 332 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1680363874
transform 1 0 340 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1680363874
transform 1 0 324 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4684
timestamp 1680363874
transform 1 0 340 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1680363874
transform 1 0 332 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1680363874
transform 1 0 364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1680363874
transform 1 0 356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4259
timestamp 1680363874
transform 1 0 356 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1680363874
transform 1 0 396 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4784
timestamp 1680363874
transform 1 0 396 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4182
timestamp 1680363874
transform 1 0 412 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1680363874
transform 1 0 436 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4601
timestamp 1680363874
transform 1 0 412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1680363874
transform 1 0 428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1680363874
transform 1 0 436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1680363874
transform 1 0 420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1680363874
transform 1 0 436 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4260
timestamp 1680363874
transform 1 0 428 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1680363874
transform 1 0 436 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4688
timestamp 1680363874
transform 1 0 460 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4145
timestamp 1680363874
transform 1 0 540 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4604
timestamp 1680363874
transform 1 0 516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1680363874
transform 1 0 532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1680363874
transform 1 0 524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1680363874
transform 1 0 540 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4299
timestamp 1680363874
transform 1 0 540 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1680363874
transform 1 0 604 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1680363874
transform 1 0 612 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4606
timestamp 1680363874
transform 1 0 620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1680363874
transform 1 0 612 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4261
timestamp 1680363874
transform 1 0 612 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4692
timestamp 1680363874
transform 1 0 636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1680363874
transform 1 0 652 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_4184
timestamp 1680363874
transform 1 0 732 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4607
timestamp 1680363874
transform 1 0 732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1680363874
transform 1 0 740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1680363874
transform 1 0 756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1680363874
transform 1 0 764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1680363874
transform 1 0 764 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4216
timestamp 1680363874
transform 1 0 780 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4695
timestamp 1680363874
transform 1 0 788 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4217
timestamp 1680363874
transform 1 0 820 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4696
timestamp 1680363874
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4262
timestamp 1680363874
transform 1 0 812 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4609
timestamp 1680363874
transform 1 0 828 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4147
timestamp 1680363874
transform 1 0 868 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1680363874
transform 1 0 860 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4610
timestamp 1680363874
transform 1 0 860 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4263
timestamp 1680363874
transform 1 0 860 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4786
timestamp 1680363874
transform 1 0 884 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1680363874
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1680363874
transform 1 0 940 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4264
timestamp 1680363874
transform 1 0 940 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4611
timestamp 1680363874
transform 1 0 956 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4233
timestamp 1680363874
transform 1 0 964 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1680363874
transform 1 0 956 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4699
timestamp 1680363874
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4148
timestamp 1680363874
transform 1 0 1012 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1680363874
transform 1 0 1004 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4612
timestamp 1680363874
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1680363874
transform 1 0 1020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1680363874
transform 1 0 996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1680363874
transform 1 0 1012 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4266
timestamp 1680363874
transform 1 0 1012 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1680363874
transform 1 0 1004 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1680363874
transform 1 0 1036 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1680363874
transform 1 0 1044 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4702
timestamp 1680363874
transform 1 0 1060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1680363874
transform 1 0 1076 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1680363874
transform 1 0 1084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1680363874
transform 1 0 1100 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4234
timestamp 1680363874
transform 1 0 1084 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1680363874
transform 1 0 1108 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4703
timestamp 1680363874
transform 1 0 1108 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4302
timestamp 1680363874
transform 1 0 1148 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4704
timestamp 1680363874
transform 1 0 1180 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4267
timestamp 1680363874
transform 1 0 1180 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4787
timestamp 1680363874
transform 1 0 1196 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1680363874
transform 1 0 1180 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1680363874
transform 1 0 1188 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_4303
timestamp 1680363874
transform 1 0 1196 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1680363874
transform 1 0 1268 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1680363874
transform 1 0 1252 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4616
timestamp 1680363874
transform 1 0 1252 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4219
timestamp 1680363874
transform 1 0 1260 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4617
timestamp 1680363874
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1680363874
transform 1 0 1260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1680363874
transform 1 0 1276 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4268
timestamp 1680363874
transform 1 0 1284 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4618
timestamp 1680363874
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4304
timestamp 1680363874
transform 1 0 1308 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4707
timestamp 1680363874
transform 1 0 1324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1680363874
transform 1 0 1332 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4269
timestamp 1680363874
transform 1 0 1332 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4709
timestamp 1680363874
transform 1 0 1356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4235
timestamp 1680363874
transform 1 0 1396 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4710
timestamp 1680363874
transform 1 0 1404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1680363874
transform 1 0 1428 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4188
timestamp 1680363874
transform 1 0 1468 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1680363874
transform 1 0 1508 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1680363874
transform 1 0 1500 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4619
timestamp 1680363874
transform 1 0 1460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1680363874
transform 1 0 1468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1680363874
transform 1 0 1484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1680363874
transform 1 0 1500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1680363874
transform 1 0 1508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1680363874
transform 1 0 1476 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4236
timestamp 1680363874
transform 1 0 1484 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4713
timestamp 1680363874
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4237
timestamp 1680363874
transform 1 0 1508 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1680363874
transform 1 0 1516 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1680363874
transform 1 0 1580 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4624
timestamp 1680363874
transform 1 0 1564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1680363874
transform 1 0 1580 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4238
timestamp 1680363874
transform 1 0 1548 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4714
timestamp 1680363874
transform 1 0 1556 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1680363874
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4220
timestamp 1680363874
transform 1 0 1588 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4716
timestamp 1680363874
transform 1 0 1588 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4168
timestamp 1680363874
transform 1 0 1604 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4626
timestamp 1680363874
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4190
timestamp 1680363874
transform 1 0 1612 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4717
timestamp 1680363874
transform 1 0 1636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1680363874
transform 1 0 1660 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4151
timestamp 1680363874
transform 1 0 1692 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1680363874
transform 1 0 1700 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4628
timestamp 1680363874
transform 1 0 1684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1680363874
transform 1 0 1700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1680363874
transform 1 0 1676 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1680363874
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4270
timestamp 1680363874
transform 1 0 1684 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1680363874
transform 1 0 1724 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1680363874
transform 1 0 1796 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1680363874
transform 1 0 1804 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4679
timestamp 1680363874
transform 1 0 1740 0 1 2533
box -2 -2 2 2
use M3_M2  M3_M2_4239
timestamp 1680363874
transform 1 0 1740 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4720
timestamp 1680363874
transform 1 0 1764 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4271
timestamp 1680363874
transform 1 0 1764 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1680363874
transform 1 0 1756 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1680363874
transform 1 0 1740 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1680363874
transform 1 0 1844 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1680363874
transform 1 0 1860 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4721
timestamp 1680363874
transform 1 0 1860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1680363874
transform 1 0 1956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1680363874
transform 1 0 1956 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1680363874
transform 1 0 1972 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1680363874
transform 1 0 1964 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1680363874
transform 1 0 1988 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4240
timestamp 1680363874
transform 1 0 2012 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4630
timestamp 1680363874
transform 1 0 2028 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4337
timestamp 1680363874
transform 1 0 2020 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1680363874
transform 1 0 2068 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4631
timestamp 1680363874
transform 1 0 2140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1680363874
transform 1 0 2148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1680363874
transform 1 0 2164 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4241
timestamp 1680363874
transform 1 0 2148 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4724
timestamp 1680363874
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1680363874
transform 1 0 2172 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4272
timestamp 1680363874
transform 1 0 2156 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1680363874
transform 1 0 2188 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4634
timestamp 1680363874
transform 1 0 2188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1680363874
transform 1 0 2188 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4273
timestamp 1680363874
transform 1 0 2188 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4635
timestamp 1680363874
transform 1 0 2260 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4242
timestamp 1680363874
transform 1 0 2260 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1680363874
transform 1 0 2356 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4636
timestamp 1680363874
transform 1 0 2308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1680363874
transform 1 0 2356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1680363874
transform 1 0 2396 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4192
timestamp 1680363874
transform 1 0 2460 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4637
timestamp 1680363874
transform 1 0 2444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1680363874
transform 1 0 2460 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4338
timestamp 1680363874
transform 1 0 2436 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4729
timestamp 1680363874
transform 1 0 2452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1680363874
transform 1 0 2468 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4156
timestamp 1680363874
transform 1 0 2500 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1680363874
transform 1 0 2492 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4639
timestamp 1680363874
transform 1 0 2492 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4274
timestamp 1680363874
transform 1 0 2500 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1680363874
transform 1 0 2548 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4640
timestamp 1680363874
transform 1 0 2516 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4243
timestamp 1680363874
transform 1 0 2516 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4731
timestamp 1680363874
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4244
timestamp 1680363874
transform 1 0 2588 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1680363874
transform 1 0 2540 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1680363874
transform 1 0 2620 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4641
timestamp 1680363874
transform 1 0 2620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1680363874
transform 1 0 2612 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4195
timestamp 1680363874
transform 1 0 2636 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4733
timestamp 1680363874
transform 1 0 2628 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4171
timestamp 1680363874
transform 1 0 2652 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1680363874
transform 1 0 2652 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4642
timestamp 1680363874
transform 1 0 2676 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4245
timestamp 1680363874
transform 1 0 2676 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4734
timestamp 1680363874
transform 1 0 2700 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4246
timestamp 1680363874
transform 1 0 2756 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1680363874
transform 1 0 2676 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1680363874
transform 1 0 2668 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1680363874
transform 1 0 2700 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1680363874
transform 1 0 2788 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4643
timestamp 1680363874
transform 1 0 2788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1680363874
transform 1 0 2780 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4277
timestamp 1680363874
transform 1 0 2780 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4736
timestamp 1680363874
transform 1 0 2820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1680363874
transform 1 0 2836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1680363874
transform 1 0 2876 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1680363874
transform 1 0 2884 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4247
timestamp 1680363874
transform 1 0 2868 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4790
timestamp 1680363874
transform 1 0 2868 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4278
timestamp 1680363874
transform 1 0 2884 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1680363874
transform 1 0 2876 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4738
timestamp 1680363874
transform 1 0 2900 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4248
timestamp 1680363874
transform 1 0 2916 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4791
timestamp 1680363874
transform 1 0 2916 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4197
timestamp 1680363874
transform 1 0 3060 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4646
timestamp 1680363874
transform 1 0 3052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1680363874
transform 1 0 3060 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4249
timestamp 1680363874
transform 1 0 3052 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4739
timestamp 1680363874
transform 1 0 3076 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4172
timestamp 1680363874
transform 1 0 3092 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4648
timestamp 1680363874
transform 1 0 3092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1680363874
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4221
timestamp 1680363874
transform 1 0 3108 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1680363874
transform 1 0 3100 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1680363874
transform 1 0 3092 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1680363874
transform 1 0 3132 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1680363874
transform 1 0 3132 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4649
timestamp 1680363874
transform 1 0 3140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1680363874
transform 1 0 3132 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4323
timestamp 1680363874
transform 1 0 3124 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4792
timestamp 1680363874
transform 1 0 3156 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4159
timestamp 1680363874
transform 1 0 3172 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4742
timestamp 1680363874
transform 1 0 3172 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4280
timestamp 1680363874
transform 1 0 3172 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1680363874
transform 1 0 3204 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4650
timestamp 1680363874
transform 1 0 3204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1680363874
transform 1 0 3220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1680363874
transform 1 0 3228 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4281
timestamp 1680363874
transform 1 0 3228 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1680363874
transform 1 0 3220 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1680363874
transform 1 0 3244 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4651
timestamp 1680363874
transform 1 0 3260 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4160
timestamp 1680363874
transform 1 0 3284 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1680363874
transform 1 0 3276 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4745
timestamp 1680363874
transform 1 0 3284 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4173
timestamp 1680363874
transform 1 0 3324 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1680363874
transform 1 0 3300 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4652
timestamp 1680363874
transform 1 0 3324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1680363874
transform 1 0 3332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1680363874
transform 1 0 3316 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4282
timestamp 1680363874
transform 1 0 3332 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1680363874
transform 1 0 3380 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4654
timestamp 1680363874
transform 1 0 3404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1680363874
transform 1 0 3436 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4326
timestamp 1680363874
transform 1 0 3420 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1680363874
transform 1 0 3420 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1680363874
transform 1 0 3492 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4748
timestamp 1680363874
transform 1 0 3508 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4174
timestamp 1680363874
transform 1 0 3540 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1680363874
transform 1 0 3540 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4749
timestamp 1680363874
transform 1 0 3540 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4250
timestamp 1680363874
transform 1 0 3556 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4793
timestamp 1680363874
transform 1 0 3556 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4226
timestamp 1680363874
transform 1 0 3580 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4655
timestamp 1680363874
transform 1 0 3588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1680363874
transform 1 0 3572 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4311
timestamp 1680363874
transform 1 0 3572 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1680363874
transform 1 0 3596 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4656
timestamp 1680363874
transform 1 0 3596 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4251
timestamp 1680363874
transform 1 0 3588 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1680363874
transform 1 0 3612 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4657
timestamp 1680363874
transform 1 0 3620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1680363874
transform 1 0 3708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1680363874
transform 1 0 3612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1680363874
transform 1 0 3628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1680363874
transform 1 0 3684 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4283
timestamp 1680363874
transform 1 0 3612 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1680363874
transform 1 0 3628 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1680363874
transform 1 0 3692 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1680363874
transform 1 0 3708 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1680363874
transform 1 0 3724 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4753
timestamp 1680363874
transform 1 0 3732 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4284
timestamp 1680363874
transform 1 0 3732 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1680363874
transform 1 0 3748 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1680363874
transform 1 0 3788 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4659
timestamp 1680363874
transform 1 0 3788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1680363874
transform 1 0 3804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1680363874
transform 1 0 3812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1680363874
transform 1 0 3796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1680363874
transform 1 0 3812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4286
timestamp 1680363874
transform 1 0 3780 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1680363874
transform 1 0 3812 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1680363874
transform 1 0 3884 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4662
timestamp 1680363874
transform 1 0 3884 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4203
timestamp 1680363874
transform 1 0 3916 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4663
timestamp 1680363874
transform 1 0 3916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1680363874
transform 1 0 3908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1680363874
transform 1 0 3916 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4312
timestamp 1680363874
transform 1 0 3900 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1680363874
transform 1 0 3916 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4664
timestamp 1680363874
transform 1 0 3956 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1680363874
transform 1 0 3964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1680363874
transform 1 0 3948 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1680363874
transform 1 0 3964 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4288
timestamp 1680363874
transform 1 0 3940 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1680363874
transform 1 0 3964 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1680363874
transform 1 0 3940 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4760
timestamp 1680363874
transform 1 0 4020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1680363874
transform 1 0 4036 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4290
timestamp 1680363874
transform 1 0 4036 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1680363874
transform 1 0 4028 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4666
timestamp 1680363874
transform 1 0 4060 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4329
timestamp 1680363874
transform 1 0 4084 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1680363874
transform 1 0 4140 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4667
timestamp 1680363874
transform 1 0 4140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1680363874
transform 1 0 4108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1680363874
transform 1 0 4124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1680363874
transform 1 0 4140 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4314
timestamp 1680363874
transform 1 0 4108 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1680363874
transform 1 0 4132 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1680363874
transform 1 0 4108 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1680363874
transform 1 0 4140 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1680363874
transform 1 0 4196 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4668
timestamp 1680363874
transform 1 0 4204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1680363874
transform 1 0 4196 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4252
timestamp 1680363874
transform 1 0 4204 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1680363874
transform 1 0 4228 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4669
timestamp 1680363874
transform 1 0 4228 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4291
timestamp 1680363874
transform 1 0 4220 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1680363874
transform 1 0 4236 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1680363874
transform 1 0 4252 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4596
timestamp 1680363874
transform 1 0 4252 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1680363874
transform 1 0 4244 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4292
timestamp 1680363874
transform 1 0 4244 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1680363874
transform 1 0 4276 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1680363874
transform 1 0 4268 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4670
timestamp 1680363874
transform 1 0 4268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1680363874
transform 1 0 4268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1680363874
transform 1 0 4276 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4316
timestamp 1680363874
transform 1 0 4276 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1680363874
transform 1 0 4292 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1680363874
transform 1 0 4316 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1680363874
transform 1 0 4308 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4671
timestamp 1680363874
transform 1 0 4316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1680363874
transform 1 0 4332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1680363874
transform 1 0 4340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1680363874
transform 1 0 4308 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4253
timestamp 1680363874
transform 1 0 4316 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4770
timestamp 1680363874
transform 1 0 4324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1680363874
transform 1 0 4340 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4293
timestamp 1680363874
transform 1 0 4340 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1680363874
transform 1 0 4332 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1680363874
transform 1 0 4340 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1680363874
transform 1 0 4412 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1680363874
transform 1 0 4484 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1680363874
transform 1 0 4396 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4674
timestamp 1680363874
transform 1 0 4484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1680363874
transform 1 0 4396 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1680363874
transform 1 0 4404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1680363874
transform 1 0 4436 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4294
timestamp 1680363874
transform 1 0 4396 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1680363874
transform 1 0 4436 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1680363874
transform 1 0 4404 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1680363874
transform 1 0 4428 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1680363874
transform 1 0 4500 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1680363874
transform 1 0 4516 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1680363874
transform 1 0 4580 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4675
timestamp 1680363874
transform 1 0 4516 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4255
timestamp 1680363874
transform 1 0 4516 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4775
timestamp 1680363874
transform 1 0 4564 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4296
timestamp 1680363874
transform 1 0 4564 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1680363874
transform 1 0 4580 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1680363874
transform 1 0 4636 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1680363874
transform 1 0 4612 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4676
timestamp 1680363874
transform 1 0 4636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1680363874
transform 1 0 4604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1680363874
transform 1 0 4612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1680363874
transform 1 0 4628 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4256
timestamp 1680363874
transform 1 0 4636 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4779
timestamp 1680363874
transform 1 0 4644 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4319
timestamp 1680363874
transform 1 0 4644 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1680363874
transform 1 0 4620 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1680363874
transform 1 0 4660 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4677
timestamp 1680363874
transform 1 0 4684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1680363874
transform 1 0 4676 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4257
timestamp 1680363874
transform 1 0 4684 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4781
timestamp 1680363874
transform 1 0 4692 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4297
timestamp 1680363874
transform 1 0 4676 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4678
timestamp 1680363874
transform 1 0 4788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1680363874
transform 1 0 4764 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4320
timestamp 1680363874
transform 1 0 4708 0 1 2505
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_44
timestamp 1680363874
transform 1 0 24 0 1 2470
box -10 -3 10 3
use FILL  FILL_4690
timestamp 1680363874
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1680363874
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1680363874
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1680363874
transform 1 0 96 0 -1 2570
box -7 -3 39 105
use FILL  FILL_4697
timestamp 1680363874
transform 1 0 128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1680363874
transform 1 0 136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1680363874
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1680363874
transform 1 0 152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1680363874
transform 1 0 160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1680363874
transform 1 0 168 0 -1 2570
box -8 -3 16 105
use FAX1  FAX1_8
timestamp 1680363874
transform -1 0 296 0 -1 2570
box -5 -3 126 105
use FILL  FILL_4712
timestamp 1680363874
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1680363874
transform 1 0 304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1680363874
transform 1 0 312 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_10
timestamp 1680363874
transform -1 0 352 0 -1 2570
box -8 -3 40 105
use FILL  FILL_4715
timestamp 1680363874
transform 1 0 352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1680363874
transform 1 0 360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1680363874
transform 1 0 368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1680363874
transform 1 0 376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1680363874
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1680363874
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_158
timestamp 1680363874
transform -1 0 440 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4729
timestamp 1680363874
transform 1 0 440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1680363874
transform 1 0 448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1680363874
transform 1 0 456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1680363874
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1680363874
transform 1 0 472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1680363874
transform 1 0 480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1680363874
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1680363874
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_159
timestamp 1680363874
transform -1 0 544 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4742
timestamp 1680363874
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1680363874
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1680363874
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1680363874
transform 1 0 568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1680363874
transform 1 0 576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1680363874
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1680363874
transform 1 0 592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1680363874
transform 1 0 600 0 -1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_8
timestamp 1680363874
transform 1 0 608 0 -1 2570
box -7 -3 39 105
use FILL  FILL_4757
timestamp 1680363874
transform 1 0 640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1680363874
transform 1 0 648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1680363874
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1680363874
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1680363874
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1680363874
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1680363874
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1680363874
transform 1 0 696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1680363874
transform 1 0 704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1680363874
transform 1 0 712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1680363874
transform 1 0 720 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_119
timestamp 1680363874
transform 1 0 728 0 -1 2570
box -8 -3 34 105
use FILL  FILL_4781
timestamp 1680363874
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1680363874
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1680363874
transform 1 0 776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1680363874
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1680363874
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_320
timestamp 1680363874
transform -1 0 816 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4786
timestamp 1680363874
transform 1 0 816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1680363874
transform 1 0 824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1680363874
transform 1 0 832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1680363874
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_10
timestamp 1680363874
transform 1 0 848 0 -1 2570
box -7 -3 39 105
use FILL  FILL_4793
timestamp 1680363874
transform 1 0 880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1680363874
transform 1 0 888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1680363874
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1680363874
transform 1 0 904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1680363874
transform 1 0 912 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_120
timestamp 1680363874
transform -1 0 952 0 -1 2570
box -8 -3 34 105
use FILL  FILL_4803
timestamp 1680363874
transform 1 0 952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1680363874
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1680363874
transform 1 0 968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1680363874
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1680363874
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_163
timestamp 1680363874
transform -1 0 1032 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4813
timestamp 1680363874
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1680363874
transform 1 0 1040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1680363874
transform 1 0 1048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1680363874
transform 1 0 1056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1680363874
transform 1 0 1064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1680363874
transform 1 0 1072 0 -1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_11
timestamp 1680363874
transform -1 0 1112 0 -1 2570
box -7 -3 39 105
use FILL  FILL_4826
timestamp 1680363874
transform 1 0 1112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1680363874
transform 1 0 1120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1680363874
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1680363874
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1680363874
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1680363874
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1680363874
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1680363874
transform 1 0 1168 0 -1 2570
box -8 -3 40 105
use FILL  FILL_4837
timestamp 1680363874
transform 1 0 1200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1680363874
transform 1 0 1208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1680363874
transform 1 0 1216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1680363874
transform 1 0 1224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1680363874
transform 1 0 1232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1680363874
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_233
timestamp 1680363874
transform 1 0 1248 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4851
timestamp 1680363874
transform 1 0 1288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1680363874
transform 1 0 1296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1680363874
transform 1 0 1304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1680363874
transform 1 0 1312 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_321
timestamp 1680363874
transform 1 0 1320 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4859
timestamp 1680363874
transform 1 0 1336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1680363874
transform 1 0 1344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1680363874
transform 1 0 1352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1680363874
transform 1 0 1360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1680363874
transform 1 0 1368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1680363874
transform 1 0 1376 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_164
timestamp 1680363874
transform 1 0 1384 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4867
timestamp 1680363874
transform 1 0 1424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1680363874
transform 1 0 1432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1680363874
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1680363874
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1680363874
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_234
timestamp 1680363874
transform -1 0 1504 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4876
timestamp 1680363874
transform 1 0 1504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1680363874
transform 1 0 1512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1680363874
transform 1 0 1520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1680363874
transform 1 0 1528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1680363874
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_235
timestamp 1680363874
transform 1 0 1544 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4881
timestamp 1680363874
transform 1 0 1584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1680363874
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1680363874
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1680363874
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_324
timestamp 1680363874
transform 1 0 1616 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4887
timestamp 1680363874
transform 1 0 1632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1680363874
transform 1 0 1640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1680363874
transform 1 0 1648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1680363874
transform 1 0 1656 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_236
timestamp 1680363874
transform 1 0 1664 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4903
timestamp 1680363874
transform 1 0 1704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1680363874
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1680363874
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_290
timestamp 1680363874
transform 1 0 1728 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4906
timestamp 1680363874
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1680363874
transform 1 0 1832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1680363874
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_325
timestamp 1680363874
transform 1 0 1848 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4912
timestamp 1680363874
transform 1 0 1864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1680363874
transform 1 0 1872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1680363874
transform 1 0 1880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1680363874
transform 1 0 1888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1680363874
transform 1 0 1896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1680363874
transform 1 0 1904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1680363874
transform 1 0 1912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1680363874
transform 1 0 1920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1680363874
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1680363874
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1680363874
transform 1 0 1944 0 -1 2570
box -8 -3 40 105
use FILL  FILL_4933
timestamp 1680363874
transform 1 0 1976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1680363874
transform 1 0 1984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1680363874
transform 1 0 1992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1680363874
transform 1 0 2000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1680363874
transform 1 0 2008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1680363874
transform 1 0 2016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1680363874
transform 1 0 2024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1680363874
transform 1 0 2032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1680363874
transform 1 0 2040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1680363874
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1680363874
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1680363874
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1680363874
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1680363874
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1680363874
transform 1 0 2088 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_326
timestamp 1680363874
transform -1 0 2112 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4955
timestamp 1680363874
transform 1 0 2112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1680363874
transform 1 0 2120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1680363874
transform 1 0 2128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1680363874
transform 1 0 2136 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_238
timestamp 1680363874
transform -1 0 2184 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4959
timestamp 1680363874
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1680363874
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1680363874
transform 1 0 2200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1680363874
transform 1 0 2208 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4346
timestamp 1680363874
transform 1 0 2228 0 1 2475
box -3 -3 3 3
use FILL  FILL_4963
timestamp 1680363874
transform 1 0 2216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1680363874
transform 1 0 2224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1680363874
transform 1 0 2232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1680363874
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_327
timestamp 1680363874
transform -1 0 2264 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4967
timestamp 1680363874
transform 1 0 2264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1680363874
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1680363874
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1680363874
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4347
timestamp 1680363874
transform 1 0 2316 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_294
timestamp 1680363874
transform 1 0 2296 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4975
timestamp 1680363874
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1680363874
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1680363874
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1680363874
transform 1 0 2416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1680363874
transform 1 0 2424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1680363874
transform 1 0 2432 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_239
timestamp 1680363874
transform 1 0 2440 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4988
timestamp 1680363874
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1680363874
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1680363874
transform 1 0 2496 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_296
timestamp 1680363874
transform 1 0 2504 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_330
timestamp 1680363874
transform 1 0 2600 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1680363874
transform 1 0 2616 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4995
timestamp 1680363874
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1680363874
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1680363874
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1680363874
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_298
timestamp 1680363874
transform 1 0 2664 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5001
timestamp 1680363874
transform 1 0 2760 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_333
timestamp 1680363874
transform 1 0 2768 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5003
timestamp 1680363874
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1680363874
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1680363874
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_121
timestamp 1680363874
transform 1 0 2808 0 -1 2570
box -8 -3 34 105
use M3_M2  M3_M2_4348
timestamp 1680363874
transform 1 0 2852 0 1 2475
box -3 -3 3 3
use FILL  FILL_5013
timestamp 1680363874
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1680363874
transform 1 0 2848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1680363874
transform 1 0 2856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1680363874
transform 1 0 2864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1680363874
transform 1 0 2872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1680363874
transform 1 0 2880 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_122
timestamp 1680363874
transform 1 0 2888 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5029
timestamp 1680363874
transform 1 0 2920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1680363874
transform 1 0 2928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1680363874
transform 1 0 2936 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4349
timestamp 1680363874
transform 1 0 2956 0 1 2475
box -3 -3 3 3
use FILL  FILL_5035
timestamp 1680363874
transform 1 0 2944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1680363874
transform 1 0 2952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1680363874
transform 1 0 2960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1680363874
transform 1 0 2968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1680363874
transform 1 0 2976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1680363874
transform 1 0 2984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1680363874
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1680363874
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1680363874
transform 1 0 3008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1680363874
transform 1 0 3016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1680363874
transform 1 0 3024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1680363874
transform 1 0 3032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1680363874
transform 1 0 3040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1680363874
transform 1 0 3048 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_334
timestamp 1680363874
transform 1 0 3056 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5061
timestamp 1680363874
transform 1 0 3072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1680363874
transform 1 0 3080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1680363874
transform 1 0 3088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1680363874
transform 1 0 3096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1680363874
transform 1 0 3104 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_168
timestamp 1680363874
transform 1 0 3112 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5070
timestamp 1680363874
transform 1 0 3152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1680363874
transform 1 0 3160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1680363874
transform 1 0 3168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1680363874
transform 1 0 3176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1680363874
transform 1 0 3184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1680363874
transform 1 0 3192 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_125
timestamp 1680363874
transform -1 0 3232 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5077
timestamp 1680363874
transform 1 0 3232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1680363874
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1680363874
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1680363874
transform 1 0 3256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1680363874
transform 1 0 3264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1680363874
transform 1 0 3272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1680363874
transform 1 0 3280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1680363874
transform 1 0 3288 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_169
timestamp 1680363874
transform -1 0 3336 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5092
timestamp 1680363874
transform 1 0 3336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1680363874
transform 1 0 3344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1680363874
transform 1 0 3352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1680363874
transform 1 0 3360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1680363874
transform 1 0 3368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1680363874
transform 1 0 3376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1680363874
transform 1 0 3384 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4350
timestamp 1680363874
transform 1 0 3444 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_300
timestamp 1680363874
transform 1 0 3392 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5114
timestamp 1680363874
transform 1 0 3488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1680363874
transform 1 0 3496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1680363874
transform 1 0 3504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1680363874
transform 1 0 3512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1680363874
transform 1 0 3520 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_126
timestamp 1680363874
transform 1 0 3528 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5123
timestamp 1680363874
transform 1 0 3560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1680363874
transform 1 0 3568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1680363874
transform 1 0 3576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1680363874
transform 1 0 3584 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4351
timestamp 1680363874
transform 1 0 3612 0 1 2475
box -3 -3 3 3
use OAI21X1  OAI21X1_127
timestamp 1680363874
transform -1 0 3624 0 -1 2570
box -8 -3 34 105
use M3_M2  M3_M2_4352
timestamp 1680363874
transform 1 0 3636 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_301
timestamp 1680363874
transform -1 0 3720 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5145
timestamp 1680363874
transform 1 0 3720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1680363874
transform 1 0 3728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1680363874
transform 1 0 3736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1680363874
transform 1 0 3744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1680363874
transform 1 0 3752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1680363874
transform 1 0 3760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1680363874
transform 1 0 3768 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4353
timestamp 1680363874
transform 1 0 3812 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_172
timestamp 1680363874
transform 1 0 3776 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5159
timestamp 1680363874
transform 1 0 3816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1680363874
transform 1 0 3824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1680363874
transform 1 0 3832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1680363874
transform 1 0 3840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1680363874
transform 1 0 3848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1680363874
transform 1 0 3856 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_338
timestamp 1680363874
transform 1 0 3864 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5170
timestamp 1680363874
transform 1 0 3880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1680363874
transform 1 0 3888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1680363874
transform 1 0 3896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1680363874
transform 1 0 3904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1680363874
transform 1 0 3912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1680363874
transform 1 0 3920 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_174
timestamp 1680363874
transform 1 0 3928 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5182
timestamp 1680363874
transform 1 0 3968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1680363874
transform 1 0 3976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1680363874
transform 1 0 3984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1680363874
transform 1 0 3992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1680363874
transform 1 0 4000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1680363874
transform 1 0 4008 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_339
timestamp 1680363874
transform 1 0 4016 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5193
timestamp 1680363874
transform 1 0 4032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1680363874
transform 1 0 4040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1680363874
transform 1 0 4048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1680363874
transform 1 0 4056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1680363874
transform 1 0 4064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1680363874
transform 1 0 4072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1680363874
transform 1 0 4080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1680363874
transform 1 0 4088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1680363874
transform 1 0 4096 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_175
timestamp 1680363874
transform -1 0 4144 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5209
timestamp 1680363874
transform 1 0 4144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1680363874
transform 1 0 4152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1680363874
transform 1 0 4160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1680363874
transform 1 0 4168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1680363874
transform 1 0 4176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1680363874
transform 1 0 4184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1680363874
transform 1 0 4192 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_49
timestamp 1680363874
transform -1 0 4224 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5221
timestamp 1680363874
transform 1 0 4224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1680363874
transform 1 0 4232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1680363874
transform 1 0 4240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1680363874
transform 1 0 4248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1680363874
transform 1 0 4256 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_341
timestamp 1680363874
transform 1 0 4264 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5236
timestamp 1680363874
transform 1 0 4280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1680363874
transform 1 0 4288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1680363874
transform 1 0 4296 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_177
timestamp 1680363874
transform 1 0 4304 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5239
timestamp 1680363874
transform 1 0 4344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1680363874
transform 1 0 4352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1680363874
transform 1 0 4360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1680363874
transform 1 0 4368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1680363874
transform 1 0 4376 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_342
timestamp 1680363874
transform 1 0 4384 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_302
timestamp 1680363874
transform -1 0 4496 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5255
timestamp 1680363874
transform 1 0 4496 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_303
timestamp 1680363874
transform 1 0 4504 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5268
timestamp 1680363874
transform 1 0 4600 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_180
timestamp 1680363874
transform -1 0 4648 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5269
timestamp 1680363874
transform 1 0 4648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1680363874
transform 1 0 4656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1680363874
transform 1 0 4664 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_344
timestamp 1680363874
transform -1 0 4688 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5278
timestamp 1680363874
transform 1 0 4688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1680363874
transform 1 0 4696 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_305
timestamp 1680363874
transform -1 0 4800 0 -1 2570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_45
timestamp 1680363874
transform 1 0 4851 0 1 2470
box -10 -3 10 3
use M2_M1  M2_M1_4925
timestamp 1680363874
transform 1 0 92 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1680363874
transform 1 0 116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1680363874
transform 1 0 124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1680363874
transform 1 0 164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1680363874
transform 1 0 172 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4356
timestamp 1680363874
transform 1 0 204 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4830
timestamp 1680363874
transform 1 0 204 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4495
timestamp 1680363874
transform 1 0 204 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4929
timestamp 1680363874
transform 1 0 268 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4496
timestamp 1680363874
transform 1 0 268 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1680363874
transform 1 0 300 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4831
timestamp 1680363874
transform 1 0 300 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4395
timestamp 1680363874
transform 1 0 324 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4807
timestamp 1680363874
transform 1 0 324 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4463
timestamp 1680363874
transform 1 0 316 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4930
timestamp 1680363874
transform 1 0 324 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1680363874
transform 1 0 340 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4464
timestamp 1680363874
transform 1 0 340 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1680363874
transform 1 0 364 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1680363874
transform 1 0 364 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4808
timestamp 1680363874
transform 1 0 364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1680363874
transform 1 0 356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1680363874
transform 1 0 348 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4497
timestamp 1680363874
transform 1 0 348 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1680363874
transform 1 0 364 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1680363874
transform 1 0 380 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4809
timestamp 1680363874
transform 1 0 388 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1680363874
transform 1 0 388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1680363874
transform 1 0 420 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4373
timestamp 1680363874
transform 1 0 436 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4799
timestamp 1680363874
transform 1 0 436 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4405
timestamp 1680363874
transform 1 0 436 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4835
timestamp 1680363874
transform 1 0 444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1680363874
transform 1 0 492 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4533
timestamp 1680363874
transform 1 0 492 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1680363874
transform 1 0 500 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4810
timestamp 1680363874
transform 1 0 500 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1680363874
transform 1 0 508 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4398
timestamp 1680363874
transform 1 0 524 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1680363874
transform 1 0 524 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1680363874
transform 1 0 564 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1680363874
transform 1 0 580 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4934
timestamp 1680363874
transform 1 0 572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1680363874
transform 1 0 636 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1680363874
transform 1 0 620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1680363874
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4466
timestamp 1680363874
transform 1 0 636 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1680363874
transform 1 0 628 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1680363874
transform 1 0 620 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4936
timestamp 1680363874
transform 1 0 652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1680363874
transform 1 0 668 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4500
timestamp 1680363874
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4838
timestamp 1680363874
transform 1 0 708 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4501
timestamp 1680363874
transform 1 0 740 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1680363874
transform 1 0 756 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4938
timestamp 1680363874
transform 1 0 772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1680363874
transform 1 0 804 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4375
timestamp 1680363874
transform 1 0 836 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4812
timestamp 1680363874
transform 1 0 836 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4467
timestamp 1680363874
transform 1 0 828 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4840
timestamp 1680363874
transform 1 0 860 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4468
timestamp 1680363874
transform 1 0 860 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4939
timestamp 1680363874
transform 1 0 876 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4502
timestamp 1680363874
transform 1 0 876 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4940
timestamp 1680363874
transform 1 0 900 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4376
timestamp 1680363874
transform 1 0 940 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4813
timestamp 1680363874
transform 1 0 940 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1680363874
transform 1 0 948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1680363874
transform 1 0 948 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4408
timestamp 1680363874
transform 1 0 1012 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1680363874
transform 1 0 1004 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1680363874
transform 1 0 1044 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1680363874
transform 1 0 1068 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1680363874
transform 1 0 1060 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4814
timestamp 1680363874
transform 1 0 1068 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1680363874
transform 1 0 1044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1680363874
transform 1 0 1052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1680363874
transform 1 0 1068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1680363874
transform 1 0 1036 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1680363874
transform 1 0 1076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1680363874
transform 1 0 1100 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1680363874
transform 1 0 1108 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4378
timestamp 1680363874
transform 1 0 1164 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4800
timestamp 1680363874
transform 1 0 1148 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1680363874
transform 1 0 1164 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1680363874
transform 1 0 1140 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4400
timestamp 1680363874
transform 1 0 1172 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4816
timestamp 1680363874
transform 1 0 1172 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1680363874
transform 1 0 1180 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4410
timestamp 1680363874
transform 1 0 1220 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4946
timestamp 1680363874
transform 1 0 1212 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4535
timestamp 1680363874
transform 1 0 1212 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4846
timestamp 1680363874
transform 1 0 1268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1680363874
transform 1 0 1236 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4504
timestamp 1680363874
transform 1 0 1236 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1680363874
transform 1 0 1252 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1680363874
transform 1 0 1276 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4847
timestamp 1680363874
transform 1 0 1324 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4411
timestamp 1680363874
transform 1 0 1372 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4848
timestamp 1680363874
transform 1 0 1356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1680363874
transform 1 0 1372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1680363874
transform 1 0 1388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1680363874
transform 1 0 1340 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4469
timestamp 1680363874
transform 1 0 1348 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1680363874
transform 1 0 1356 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1680363874
transform 1 0 1388 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1680363874
transform 1 0 1428 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1680363874
transform 1 0 1420 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1680363874
transform 1 0 1436 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4851
timestamp 1680363874
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1680363874
transform 1 0 1436 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4439
timestamp 1680363874
transform 1 0 1444 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4853
timestamp 1680363874
transform 1 0 1452 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4440
timestamp 1680363874
transform 1 0 1476 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4949
timestamp 1680363874
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1680363874
transform 1 0 1428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1680363874
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1680363874
transform 1 0 1460 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4471
timestamp 1680363874
transform 1 0 1468 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1680363874
transform 1 0 1500 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1680363874
transform 1 0 1500 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1680363874
transform 1 0 1580 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4854
timestamp 1680363874
transform 1 0 1564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1680363874
transform 1 0 1516 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4472
timestamp 1680363874
transform 1 0 1564 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1680363874
transform 1 0 1580 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1680363874
transform 1 0 1612 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4855
timestamp 1680363874
transform 1 0 1612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1680363874
transform 1 0 1652 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4536
timestamp 1680363874
transform 1 0 1668 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_5009
timestamp 1680363874
transform 1 0 1676 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1680363874
transform 1 0 1796 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1680363874
transform 1 0 1732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1680363874
transform 1 0 1788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1680363874
transform 1 0 1708 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4473
timestamp 1680363874
transform 1 0 1780 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1680363874
transform 1 0 1788 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1680363874
transform 1 0 1844 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1680363874
transform 1 0 1828 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4802
timestamp 1680363874
transform 1 0 1852 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1680363874
transform 1 0 1852 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1680363874
transform 1 0 1860 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1680363874
transform 1 0 1844 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4442
timestamp 1680363874
transform 1 0 1852 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1680363874
transform 1 0 1860 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_5010
timestamp 1680363874
transform 1 0 1860 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4359
timestamp 1680363874
transform 1 0 1884 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4803
timestamp 1680363874
transform 1 0 1876 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1680363874
transform 1 0 1900 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4380
timestamp 1680363874
transform 1 0 1932 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4804
timestamp 1680363874
transform 1 0 1924 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1680363874
transform 1 0 1932 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1680363874
transform 1 0 1940 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4354
timestamp 1680363874
transform 1 0 1964 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4860
timestamp 1680363874
transform 1 0 1980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1680363874
transform 1 0 1996 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4443
timestamp 1680363874
transform 1 0 2004 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4821
timestamp 1680363874
transform 1 0 2020 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1680363874
transform 1 0 2012 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4475
timestamp 1680363874
transform 1 0 1980 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4955
timestamp 1680363874
transform 1 0 1988 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4476
timestamp 1680363874
transform 1 0 2004 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1680363874
transform 1 0 1980 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1680363874
transform 1 0 2052 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1680363874
transform 1 0 2044 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4805
timestamp 1680363874
transform 1 0 2060 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4415
timestamp 1680363874
transform 1 0 2060 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1680363874
transform 1 0 2084 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1680363874
transform 1 0 2068 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4863
timestamp 1680363874
transform 1 0 2076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1680363874
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4538
timestamp 1680363874
transform 1 0 2052 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4822
timestamp 1680363874
transform 1 0 2100 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4478
timestamp 1680363874
transform 1 0 2100 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1680363874
transform 1 0 2156 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4864
timestamp 1680363874
transform 1 0 2172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1680363874
transform 1 0 2164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1680363874
transform 1 0 2212 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4479
timestamp 1680363874
transform 1 0 2220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1680363874
transform 1 0 2252 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4865
timestamp 1680363874
transform 1 0 2236 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4445
timestamp 1680363874
transform 1 0 2244 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4866
timestamp 1680363874
transform 1 0 2252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1680363874
transform 1 0 2244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4480
timestamp 1680363874
transform 1 0 2252 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4960
timestamp 1680363874
transform 1 0 2260 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4539
timestamp 1680363874
transform 1 0 2268 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4823
timestamp 1680363874
transform 1 0 2284 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1680363874
transform 1 0 2300 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4384
timestamp 1680363874
transform 1 0 2364 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1680363874
transform 1 0 2340 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4867
timestamp 1680363874
transform 1 0 2340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1680363874
transform 1 0 2316 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4385
timestamp 1680363874
transform 1 0 2412 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4868
timestamp 1680363874
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1680363874
transform 1 0 2420 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4540
timestamp 1680363874
transform 1 0 2404 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1680363874
transform 1 0 2420 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4962
timestamp 1680363874
transform 1 0 2436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1680363874
transform 1 0 2452 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4386
timestamp 1680363874
transform 1 0 2492 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1680363874
transform 1 0 2516 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1680363874
transform 1 0 2508 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4871
timestamp 1680363874
transform 1 0 2492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1680363874
transform 1 0 2508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1680363874
transform 1 0 2500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1680363874
transform 1 0 2516 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1680363874
transform 1 0 2596 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4388
timestamp 1680363874
transform 1 0 2612 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1680363874
transform 1 0 2612 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1680363874
transform 1 0 2628 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1680363874
transform 1 0 2620 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4874
timestamp 1680363874
transform 1 0 2628 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4421
timestamp 1680363874
transform 1 0 2692 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4875
timestamp 1680363874
transform 1 0 2676 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4447
timestamp 1680363874
transform 1 0 2684 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4876
timestamp 1680363874
transform 1 0 2692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1680363874
transform 1 0 2652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1680363874
transform 1 0 2668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1680363874
transform 1 0 2684 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4542
timestamp 1680363874
transform 1 0 2652 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1680363874
transform 1 0 2724 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1680363874
transform 1 0 2780 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4877
timestamp 1680363874
transform 1 0 2732 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4448
timestamp 1680363874
transform 1 0 2740 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4878
timestamp 1680363874
transform 1 0 2780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1680363874
transform 1 0 2708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1680363874
transform 1 0 2724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1680363874
transform 1 0 2740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1680363874
transform 1 0 2756 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4511
timestamp 1680363874
transform 1 0 2788 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1680363874
transform 1 0 2804 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1680363874
transform 1 0 2756 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1680363874
transform 1 0 2860 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1680363874
transform 1 0 2876 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4879
timestamp 1680363874
transform 1 0 2868 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4361
timestamp 1680363874
transform 1 0 2900 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4880
timestamp 1680363874
transform 1 0 2916 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4362
timestamp 1680363874
transform 1 0 2932 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4825
timestamp 1680363874
transform 1 0 2932 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4450
timestamp 1680363874
transform 1 0 2932 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1680363874
transform 1 0 2948 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4972
timestamp 1680363874
transform 1 0 2948 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1680363874
transform 1 0 2972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1680363874
transform 1 0 3012 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4451
timestamp 1680363874
transform 1 0 3036 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4973
timestamp 1680363874
transform 1 0 3036 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1680363874
transform 1 0 3076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1680363874
transform 1 0 3052 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4513
timestamp 1680363874
transform 1 0 3052 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1680363874
transform 1 0 3092 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4883
timestamp 1680363874
transform 1 0 3140 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4544
timestamp 1680363874
transform 1 0 3156 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1680363874
transform 1 0 3172 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4827
timestamp 1680363874
transform 1 0 3188 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1680363874
transform 1 0 3172 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4452
timestamp 1680363874
transform 1 0 3188 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1680363874
transform 1 0 3172 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1680363874
transform 1 0 3212 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4885
timestamp 1680363874
transform 1 0 3204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1680363874
transform 1 0 3212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1680363874
transform 1 0 3284 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4453
timestamp 1680363874
transform 1 0 3308 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4976
timestamp 1680363874
transform 1 0 3308 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4515
timestamp 1680363874
transform 1 0 3308 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1680363874
transform 1 0 3324 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4887
timestamp 1680363874
transform 1 0 3324 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4516
timestamp 1680363874
transform 1 0 3340 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1680363874
transform 1 0 3332 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4977
timestamp 1680363874
transform 1 0 3380 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4481
timestamp 1680363874
transform 1 0 3404 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_5005
timestamp 1680363874
transform 1 0 3396 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4364
timestamp 1680363874
transform 1 0 3428 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1680363874
transform 1 0 3452 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1680363874
transform 1 0 3500 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1680363874
transform 1 0 3468 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4888
timestamp 1680363874
transform 1 0 3468 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4454
timestamp 1680363874
transform 1 0 3492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1680363874
transform 1 0 3508 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4889
timestamp 1680363874
transform 1 0 3500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1680363874
transform 1 0 3508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1680363874
transform 1 0 3420 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4517
timestamp 1680363874
transform 1 0 3436 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1680363874
transform 1 0 3460 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1680363874
transform 1 0 3532 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4891
timestamp 1680363874
transform 1 0 3556 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4519
timestamp 1680363874
transform 1 0 3556 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1680363874
transform 1 0 3556 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4892
timestamp 1680363874
transform 1 0 3596 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4455
timestamp 1680363874
transform 1 0 3612 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4979
timestamp 1680363874
transform 1 0 3572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1680363874
transform 1 0 3580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4520
timestamp 1680363874
transform 1 0 3572 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1680363874
transform 1 0 3596 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4981
timestamp 1680363874
transform 1 0 3612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4521
timestamp 1680363874
transform 1 0 3604 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4893
timestamp 1680363874
transform 1 0 3636 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4549
timestamp 1680363874
transform 1 0 3668 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4894
timestamp 1680363874
transform 1 0 3684 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4367
timestamp 1680363874
transform 1 0 3708 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4982
timestamp 1680363874
transform 1 0 3700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1680363874
transform 1 0 3764 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4368
timestamp 1680363874
transform 1 0 3788 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1680363874
transform 1 0 3812 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1680363874
transform 1 0 3804 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1680363874
transform 1 0 3836 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4896
timestamp 1680363874
transform 1 0 3812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1680363874
transform 1 0 3828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1680363874
transform 1 0 3836 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1680363874
transform 1 0 3804 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1680363874
transform 1 0 3844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1680363874
transform 1 0 3852 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4522
timestamp 1680363874
transform 1 0 3844 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4899
timestamp 1680363874
transform 1 0 3908 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4456
timestamp 1680363874
transform 1 0 3940 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4986
timestamp 1680363874
transform 1 0 3940 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4523
timestamp 1680363874
transform 1 0 3900 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1680363874
transform 1 0 3876 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1680363874
transform 1 0 3924 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4900
timestamp 1680363874
transform 1 0 3956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1680363874
transform 1 0 4020 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4457
timestamp 1680363874
transform 1 0 4044 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1680363874
transform 1 0 4124 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1680363874
transform 1 0 4116 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4902
timestamp 1680363874
transform 1 0 4060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1680363874
transform 1 0 4116 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4483
timestamp 1680363874
transform 1 0 4020 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4987
timestamp 1680363874
transform 1 0 4044 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4524
timestamp 1680363874
transform 1 0 4044 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4988
timestamp 1680363874
transform 1 0 4140 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4525
timestamp 1680363874
transform 1 0 4140 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1680363874
transform 1 0 4156 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4904
timestamp 1680363874
transform 1 0 4156 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4391
timestamp 1680363874
transform 1 0 4172 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4989
timestamp 1680363874
transform 1 0 4172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1680363874
transform 1 0 4204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1680363874
transform 1 0 4244 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4484
timestamp 1680363874
transform 1 0 4292 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1680363874
transform 1 0 4308 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4906
timestamp 1680363874
transform 1 0 4308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1680363874
transform 1 0 4324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1680363874
transform 1 0 4340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1680363874
transform 1 0 4300 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4485
timestamp 1680363874
transform 1 0 4308 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4991
timestamp 1680363874
transform 1 0 4316 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4369
timestamp 1680363874
transform 1 0 4356 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4909
timestamp 1680363874
transform 1 0 4356 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4526
timestamp 1680363874
transform 1 0 4356 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1680363874
transform 1 0 4348 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1680363874
transform 1 0 4380 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1680363874
transform 1 0 4396 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1680363874
transform 1 0 4412 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1680363874
transform 1 0 4420 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1680363874
transform 1 0 4436 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4828
timestamp 1680363874
transform 1 0 4444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1680363874
transform 1 0 4404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1680363874
transform 1 0 4412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1680363874
transform 1 0 4428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1680363874
transform 1 0 4396 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4487
timestamp 1680363874
transform 1 0 4404 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4993
timestamp 1680363874
transform 1 0 4420 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4488
timestamp 1680363874
transform 1 0 4428 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1680363874
transform 1 0 4420 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1680363874
transform 1 0 4412 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1680363874
transform 1 0 4444 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4994
timestamp 1680363874
transform 1 0 4444 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4403
timestamp 1680363874
transform 1 0 4500 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4913
timestamp 1680363874
transform 1 0 4500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1680363874
transform 1 0 4516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1680363874
transform 1 0 4492 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4393
timestamp 1680363874
transform 1 0 4556 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1680363874
transform 1 0 4548 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4996
timestamp 1680363874
transform 1 0 4548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4554
timestamp 1680363874
transform 1 0 4548 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1680363874
transform 1 0 4588 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1680363874
transform 1 0 4564 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4915
timestamp 1680363874
transform 1 0 4572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1680363874
transform 1 0 4588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1680363874
transform 1 0 4564 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4489
timestamp 1680363874
transform 1 0 4572 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4998
timestamp 1680363874
transform 1 0 4580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4490
timestamp 1680363874
transform 1 0 4588 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4917
timestamp 1680363874
transform 1 0 4604 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4491
timestamp 1680363874
transform 1 0 4604 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_5007
timestamp 1680363874
transform 1 0 4604 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4461
timestamp 1680363874
transform 1 0 4628 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4999
timestamp 1680363874
transform 1 0 4628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4528
timestamp 1680363874
transform 1 0 4628 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_5000
timestamp 1680363874
transform 1 0 4644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1680363874
transform 1 0 4660 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4492
timestamp 1680363874
transform 1 0 4660 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1680363874
transform 1 0 4652 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1680363874
transform 1 0 4676 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4919
timestamp 1680363874
transform 1 0 4676 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4436
timestamp 1680363874
transform 1 0 4692 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4920
timestamp 1680363874
transform 1 0 4692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1680363874
transform 1 0 4676 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4493
timestamp 1680363874
transform 1 0 4684 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1680363874
transform 1 0 4676 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1680363874
transform 1 0 4732 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4921
timestamp 1680363874
transform 1 0 4708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1680363874
transform 1 0 4716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1680363874
transform 1 0 4732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1680363874
transform 1 0 4708 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4531
timestamp 1680363874
transform 1 0 4708 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1680363874
transform 1 0 4700 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1680363874
transform 1 0 4740 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1680363874
transform 1 0 4732 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_5003
timestamp 1680363874
transform 1 0 4740 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4532
timestamp 1680363874
transform 1 0 4740 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1680363874
transform 1 0 4724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1680363874
transform 1 0 4756 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4806
timestamp 1680363874
transform 1 0 4756 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4438
timestamp 1680363874
transform 1 0 4756 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_5004
timestamp 1680363874
transform 1 0 4756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1680363874
transform 1 0 4764 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4557
timestamp 1680363874
transform 1 0 4764 0 1 2385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_46
timestamp 1680363874
transform 1 0 48 0 1 2370
box -10 -3 10 3
use FILL  FILL_5280
timestamp 1680363874
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1680363874
transform 1 0 80 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_345
timestamp 1680363874
transform 1 0 88 0 1 2370
box -9 -3 26 105
use FILL  FILL_5284
timestamp 1680363874
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1680363874
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1680363874
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1680363874
transform 1 0 128 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_346
timestamp 1680363874
transform 1 0 136 0 1 2370
box -9 -3 26 105
use FILL  FILL_5290
timestamp 1680363874
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1680363874
transform 1 0 160 0 1 2370
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1680363874
transform 1 0 168 0 1 2370
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1680363874
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1680363874
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1680363874
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1680363874
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1680363874
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1680363874
transform 1 0 216 0 1 2370
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1680363874
transform 1 0 224 0 1 2370
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1680363874
transform 1 0 232 0 1 2370
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1680363874
transform 1 0 240 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_347
timestamp 1680363874
transform 1 0 248 0 1 2370
box -9 -3 26 105
use FILL  FILL_5302
timestamp 1680363874
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1680363874
transform 1 0 272 0 1 2370
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1680363874
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1680363874
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1680363874
transform 1 0 296 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_37
timestamp 1680363874
transform 1 0 304 0 1 2370
box -8 -3 32 105
use FILL  FILL_5307
timestamp 1680363874
transform 1 0 328 0 1 2370
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1680363874
transform 1 0 336 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_348
timestamp 1680363874
transform 1 0 344 0 1 2370
box -9 -3 26 105
use NAND2X1  NAND2X1_38
timestamp 1680363874
transform -1 0 384 0 1 2370
box -8 -3 32 105
use FILL  FILL_5309
timestamp 1680363874
transform 1 0 384 0 1 2370
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1680363874
transform 1 0 392 0 1 2370
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1680363874
transform 1 0 400 0 1 2370
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1680363874
transform 1 0 408 0 1 2370
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1680363874
transform 1 0 416 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_18
timestamp 1680363874
transform -1 0 456 0 1 2370
box -8 -3 40 105
use FILL  FILL_5314
timestamp 1680363874
transform 1 0 456 0 1 2370
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1680363874
transform 1 0 464 0 1 2370
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1680363874
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1680363874
transform 1 0 480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1680363874
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1680363874
transform 1 0 496 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_349
timestamp 1680363874
transform 1 0 504 0 1 2370
box -9 -3 26 105
use FILL  FILL_5328
timestamp 1680363874
transform 1 0 520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1680363874
transform 1 0 528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1680363874
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1680363874
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1680363874
transform 1 0 552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1680363874
transform 1 0 560 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_351
timestamp 1680363874
transform 1 0 568 0 1 2370
box -9 -3 26 105
use FILL  FILL_5340
timestamp 1680363874
transform 1 0 584 0 1 2370
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1680363874
transform 1 0 592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5342
timestamp 1680363874
transform 1 0 600 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_129
timestamp 1680363874
transform 1 0 608 0 1 2370
box -8 -3 34 105
use FILL  FILL_5343
timestamp 1680363874
transform 1 0 640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1680363874
transform 1 0 648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1680363874
transform 1 0 656 0 1 2370
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1680363874
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1680363874
transform 1 0 672 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_352
timestamp 1680363874
transform 1 0 680 0 1 2370
box -9 -3 26 105
use FILL  FILL_5348
timestamp 1680363874
transform 1 0 696 0 1 2370
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1680363874
transform 1 0 704 0 1 2370
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1680363874
transform 1 0 712 0 1 2370
box -8 -3 16 105
use FILL  FILL_5351
timestamp 1680363874
transform 1 0 720 0 1 2370
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1680363874
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_5353
timestamp 1680363874
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_5354
timestamp 1680363874
transform 1 0 744 0 1 2370
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1680363874
transform 1 0 752 0 1 2370
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1680363874
transform 1 0 760 0 1 2370
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1680363874
transform 1 0 768 0 1 2370
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1680363874
transform 1 0 776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1680363874
transform 1 0 784 0 1 2370
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1680363874
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1680363874
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_5370
timestamp 1680363874
transform 1 0 808 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_39
timestamp 1680363874
transform 1 0 816 0 1 2370
box -8 -3 32 105
use FILL  FILL_5372
timestamp 1680363874
transform 1 0 840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5377
timestamp 1680363874
transform 1 0 848 0 1 2370
box -8 -3 16 105
use FILL  FILL_5379
timestamp 1680363874
transform 1 0 856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5381
timestamp 1680363874
transform 1 0 864 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_354
timestamp 1680363874
transform 1 0 872 0 1 2370
box -9 -3 26 105
use FILL  FILL_5383
timestamp 1680363874
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5384
timestamp 1680363874
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5385
timestamp 1680363874
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5386
timestamp 1680363874
transform 1 0 912 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_40
timestamp 1680363874
transform 1 0 920 0 1 2370
box -8 -3 32 105
use FILL  FILL_5387
timestamp 1680363874
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5388
timestamp 1680363874
transform 1 0 952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5389
timestamp 1680363874
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5390
timestamp 1680363874
transform 1 0 968 0 1 2370
box -8 -3 16 105
use FILL  FILL_5391
timestamp 1680363874
transform 1 0 976 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_41
timestamp 1680363874
transform -1 0 1008 0 1 2370
box -5 -3 28 105
use FILL  FILL_5392
timestamp 1680363874
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5396
timestamp 1680363874
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5398
timestamp 1680363874
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5400
timestamp 1680363874
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_130
timestamp 1680363874
transform 1 0 1040 0 1 2370
box -8 -3 34 105
use FILL  FILL_5401
timestamp 1680363874
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_5404
timestamp 1680363874
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use FILL  FILL_5406
timestamp 1680363874
transform 1 0 1088 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_355
timestamp 1680363874
transform -1 0 1112 0 1 2370
box -9 -3 26 105
use FILL  FILL_5407
timestamp 1680363874
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5412
timestamp 1680363874
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5413
timestamp 1680363874
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_5414
timestamp 1680363874
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_20
timestamp 1680363874
transform 1 0 1144 0 1 2370
box -8 -3 40 105
use FILL  FILL_5415
timestamp 1680363874
transform 1 0 1176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5420
timestamp 1680363874
transform 1 0 1184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5422
timestamp 1680363874
transform 1 0 1192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5424
timestamp 1680363874
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5426
timestamp 1680363874
transform 1 0 1208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5428
timestamp 1680363874
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4558
timestamp 1680363874
transform 1 0 1236 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_306
timestamp 1680363874
transform 1 0 1224 0 1 2370
box -8 -3 104 105
use FILL  FILL_5429
timestamp 1680363874
transform 1 0 1320 0 1 2370
box -8 -3 16 105
use FILL  FILL_5430
timestamp 1680363874
transform 1 0 1328 0 1 2370
box -8 -3 16 105
use FILL  FILL_5431
timestamp 1680363874
transform 1 0 1336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5432
timestamp 1680363874
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_182
timestamp 1680363874
transform 1 0 1352 0 1 2370
box -8 -3 46 105
use FILL  FILL_5433
timestamp 1680363874
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_5434
timestamp 1680363874
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_5435
timestamp 1680363874
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_5450
timestamp 1680363874
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_243
timestamp 1680363874
transform 1 0 1424 0 1 2370
box -8 -3 46 105
use FILL  FILL_5452
timestamp 1680363874
transform 1 0 1464 0 1 2370
box -8 -3 16 105
use FILL  FILL_5453
timestamp 1680363874
transform 1 0 1472 0 1 2370
box -8 -3 16 105
use FILL  FILL_5454
timestamp 1680363874
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5455
timestamp 1680363874
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5456
timestamp 1680363874
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1680363874
transform 1 0 1504 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_357
timestamp 1680363874
transform 1 0 1600 0 1 2370
box -9 -3 26 105
use FILL  FILL_5457
timestamp 1680363874
transform 1 0 1616 0 1 2370
box -8 -3 16 105
use FILL  FILL_5458
timestamp 1680363874
transform 1 0 1624 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4559
timestamp 1680363874
transform 1 0 1644 0 1 2375
box -3 -3 3 3
use FILL  FILL_5459
timestamp 1680363874
transform 1 0 1632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5460
timestamp 1680363874
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5461
timestamp 1680363874
transform 1 0 1648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5462
timestamp 1680363874
transform 1 0 1656 0 1 2370
box -8 -3 16 105
use FILL  FILL_5463
timestamp 1680363874
transform 1 0 1664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5464
timestamp 1680363874
transform 1 0 1672 0 1 2370
box -8 -3 16 105
use FILL  FILL_5465
timestamp 1680363874
transform 1 0 1680 0 1 2370
box -8 -3 16 105
use FILL  FILL_5475
timestamp 1680363874
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_310
timestamp 1680363874
transform 1 0 1696 0 1 2370
box -8 -3 104 105
use FILL  FILL_5477
timestamp 1680363874
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5491
timestamp 1680363874
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use FILL  FILL_5493
timestamp 1680363874
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_5495
timestamp 1680363874
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_23
timestamp 1680363874
transform -1 0 1856 0 1 2370
box -8 -3 40 105
use FILL  FILL_5496
timestamp 1680363874
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5503
timestamp 1680363874
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_5505
timestamp 1680363874
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use FILL  FILL_5507
timestamp 1680363874
transform 1 0 1880 0 1 2370
box -8 -3 16 105
use FILL  FILL_5508
timestamp 1680363874
transform 1 0 1888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5509
timestamp 1680363874
transform 1 0 1896 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_24
timestamp 1680363874
transform 1 0 1904 0 1 2370
box -8 -3 40 105
use FILL  FILL_5510
timestamp 1680363874
transform 1 0 1936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5515
timestamp 1680363874
transform 1 0 1944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5517
timestamp 1680363874
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5519
timestamp 1680363874
transform 1 0 1960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5521
timestamp 1680363874
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_184
timestamp 1680363874
transform 1 0 1976 0 1 2370
box -8 -3 46 105
use FILL  FILL_5522
timestamp 1680363874
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5523
timestamp 1680363874
transform 1 0 2024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5524
timestamp 1680363874
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use FILL  FILL_5525
timestamp 1680363874
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_5526
timestamp 1680363874
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_5527
timestamp 1680363874
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4560
timestamp 1680363874
transform 1 0 2076 0 1 2375
box -3 -3 3 3
use NAND3X1  NAND3X1_26
timestamp 1680363874
transform 1 0 2064 0 1 2370
box -8 -3 40 105
use FILL  FILL_5528
timestamp 1680363874
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5529
timestamp 1680363874
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5530
timestamp 1680363874
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5531
timestamp 1680363874
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5532
timestamp 1680363874
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use FILL  FILL_5533
timestamp 1680363874
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_5534
timestamp 1680363874
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5535
timestamp 1680363874
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5536
timestamp 1680363874
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_5537
timestamp 1680363874
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_5538
timestamp 1680363874
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5539
timestamp 1680363874
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5540
timestamp 1680363874
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5544
timestamp 1680363874
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5546
timestamp 1680363874
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5548
timestamp 1680363874
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_244
timestamp 1680363874
transform 1 0 2224 0 1 2370
box -8 -3 46 105
use FILL  FILL_5550
timestamp 1680363874
transform 1 0 2264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5551
timestamp 1680363874
transform 1 0 2272 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4561
timestamp 1680363874
transform 1 0 2292 0 1 2375
box -3 -3 3 3
use FILL  FILL_5554
timestamp 1680363874
transform 1 0 2280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5556
timestamp 1680363874
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use FILL  FILL_5558
timestamp 1680363874
transform 1 0 2296 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_313
timestamp 1680363874
transform 1 0 2304 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_359
timestamp 1680363874
transform 1 0 2400 0 1 2370
box -9 -3 26 105
use FILL  FILL_5560
timestamp 1680363874
transform 1 0 2416 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_360
timestamp 1680363874
transform -1 0 2440 0 1 2370
box -9 -3 26 105
use FILL  FILL_5561
timestamp 1680363874
transform 1 0 2440 0 1 2370
box -8 -3 16 105
use FILL  FILL_5568
timestamp 1680363874
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_5570
timestamp 1680363874
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_5572
timestamp 1680363874
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_5574
timestamp 1680363874
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_246
timestamp 1680363874
transform 1 0 2480 0 1 2370
box -8 -3 46 105
use FILL  FILL_5576
timestamp 1680363874
transform 1 0 2520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5578
timestamp 1680363874
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5580
timestamp 1680363874
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5582
timestamp 1680363874
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5584
timestamp 1680363874
transform 1 0 2552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5586
timestamp 1680363874
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5588
timestamp 1680363874
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5590
timestamp 1680363874
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_5592
timestamp 1680363874
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_5593
timestamp 1680363874
transform 1 0 2592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5594
timestamp 1680363874
transform 1 0 2600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5595
timestamp 1680363874
transform 1 0 2608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5596
timestamp 1680363874
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_5597
timestamp 1680363874
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_5599
timestamp 1680363874
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5601
timestamp 1680363874
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4562
timestamp 1680363874
transform 1 0 2684 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_249
timestamp 1680363874
transform 1 0 2648 0 1 2370
box -8 -3 46 105
use FILL  FILL_5603
timestamp 1680363874
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use FILL  FILL_5604
timestamp 1680363874
transform 1 0 2696 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4563
timestamp 1680363874
transform 1 0 2740 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_250
timestamp 1680363874
transform 1 0 2704 0 1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4564
timestamp 1680363874
transform 1 0 2812 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_315
timestamp 1680363874
transform 1 0 2744 0 1 2370
box -8 -3 104 105
use FILL  FILL_5605
timestamp 1680363874
transform 1 0 2840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5629
timestamp 1680363874
transform 1 0 2848 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_362
timestamp 1680363874
transform 1 0 2856 0 1 2370
box -9 -3 26 105
use FILL  FILL_5630
timestamp 1680363874
transform 1 0 2872 0 1 2370
box -8 -3 16 105
use FILL  FILL_5631
timestamp 1680363874
transform 1 0 2880 0 1 2370
box -8 -3 16 105
use FILL  FILL_5634
timestamp 1680363874
transform 1 0 2888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5636
timestamp 1680363874
transform 1 0 2896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5638
timestamp 1680363874
transform 1 0 2904 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_363
timestamp 1680363874
transform -1 0 2928 0 1 2370
box -9 -3 26 105
use FILL  FILL_5639
timestamp 1680363874
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use FILL  FILL_5642
timestamp 1680363874
transform 1 0 2936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5644
timestamp 1680363874
transform 1 0 2944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5646
timestamp 1680363874
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5648
timestamp 1680363874
transform 1 0 2960 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_131
timestamp 1680363874
transform 1 0 2968 0 1 2370
box -8 -3 34 105
use FILL  FILL_5650
timestamp 1680363874
transform 1 0 3000 0 1 2370
box -8 -3 16 105
use FILL  FILL_5651
timestamp 1680363874
transform 1 0 3008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5654
timestamp 1680363874
transform 1 0 3016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5656
timestamp 1680363874
transform 1 0 3024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5658
timestamp 1680363874
transform 1 0 3032 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_316
timestamp 1680363874
transform 1 0 3040 0 1 2370
box -8 -3 104 105
use FILL  FILL_5660
timestamp 1680363874
transform 1 0 3136 0 1 2370
box -8 -3 16 105
use FILL  FILL_5670
timestamp 1680363874
transform 1 0 3144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5672
timestamp 1680363874
transform 1 0 3152 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_134
timestamp 1680363874
transform 1 0 3160 0 1 2370
box -8 -3 34 105
use FILL  FILL_5674
timestamp 1680363874
transform 1 0 3192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5675
timestamp 1680363874
transform 1 0 3200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5676
timestamp 1680363874
transform 1 0 3208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5677
timestamp 1680363874
transform 1 0 3216 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_317
timestamp 1680363874
transform -1 0 3320 0 1 2370
box -8 -3 104 105
use FILL  FILL_5678
timestamp 1680363874
transform 1 0 3320 0 1 2370
box -8 -3 16 105
use FILL  FILL_5695
timestamp 1680363874
transform 1 0 3328 0 1 2370
box -8 -3 16 105
use FILL  FILL_5697
timestamp 1680363874
transform 1 0 3336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5698
timestamp 1680363874
transform 1 0 3344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5699
timestamp 1680363874
transform 1 0 3352 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_52
timestamp 1680363874
transform -1 0 3384 0 1 2370
box -8 -3 32 105
use FILL  FILL_5700
timestamp 1680363874
transform 1 0 3384 0 1 2370
box -8 -3 16 105
use FILL  FILL_5705
timestamp 1680363874
transform 1 0 3392 0 1 2370
box -8 -3 16 105
use FILL  FILL_5706
timestamp 1680363874
transform 1 0 3400 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_318
timestamp 1680363874
transform 1 0 3408 0 1 2370
box -8 -3 104 105
use FILL  FILL_5707
timestamp 1680363874
transform 1 0 3504 0 1 2370
box -8 -3 16 105
use FILL  FILL_5708
timestamp 1680363874
transform 1 0 3512 0 1 2370
box -8 -3 16 105
use FILL  FILL_5709
timestamp 1680363874
transform 1 0 3520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5713
timestamp 1680363874
transform 1 0 3528 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_367
timestamp 1680363874
transform -1 0 3552 0 1 2370
box -9 -3 26 105
use FILL  FILL_5714
timestamp 1680363874
transform 1 0 3552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5719
timestamp 1680363874
transform 1 0 3560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5721
timestamp 1680363874
transform 1 0 3568 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_185
timestamp 1680363874
transform 1 0 3576 0 1 2370
box -8 -3 46 105
use FILL  FILL_5722
timestamp 1680363874
transform 1 0 3616 0 1 2370
box -8 -3 16 105
use FILL  FILL_5725
timestamp 1680363874
transform 1 0 3624 0 1 2370
box -8 -3 16 105
use FILL  FILL_5727
timestamp 1680363874
transform 1 0 3632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5729
timestamp 1680363874
transform 1 0 3640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5731
timestamp 1680363874
transform 1 0 3648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5733
timestamp 1680363874
transform 1 0 3656 0 1 2370
box -8 -3 16 105
use FILL  FILL_5735
timestamp 1680363874
transform 1 0 3664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5736
timestamp 1680363874
transform 1 0 3672 0 1 2370
box -8 -3 16 105
use FILL  FILL_5737
timestamp 1680363874
transform 1 0 3680 0 1 2370
box -8 -3 16 105
use FILL  FILL_5738
timestamp 1680363874
transform 1 0 3688 0 1 2370
box -8 -3 16 105
use FILL  FILL_5739
timestamp 1680363874
transform 1 0 3696 0 1 2370
box -8 -3 16 105
use FILL  FILL_5740
timestamp 1680363874
transform 1 0 3704 0 1 2370
box -8 -3 16 105
use FILL  FILL_5741
timestamp 1680363874
transform 1 0 3712 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_368
timestamp 1680363874
transform 1 0 3720 0 1 2370
box -9 -3 26 105
use FILL  FILL_5742
timestamp 1680363874
transform 1 0 3736 0 1 2370
box -8 -3 16 105
use FILL  FILL_5746
timestamp 1680363874
transform 1 0 3744 0 1 2370
box -8 -3 16 105
use FILL  FILL_5748
timestamp 1680363874
transform 1 0 3752 0 1 2370
box -8 -3 16 105
use FILL  FILL_5750
timestamp 1680363874
transform 1 0 3760 0 1 2370
box -8 -3 16 105
use FILL  FILL_5752
timestamp 1680363874
transform 1 0 3768 0 1 2370
box -8 -3 16 105
use FILL  FILL_5754
timestamp 1680363874
transform 1 0 3776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5756
timestamp 1680363874
transform 1 0 3784 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_188
timestamp 1680363874
transform 1 0 3792 0 1 2370
box -8 -3 46 105
use FILL  FILL_5757
timestamp 1680363874
transform 1 0 3832 0 1 2370
box -8 -3 16 105
use FILL  FILL_5760
timestamp 1680363874
transform 1 0 3840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5762
timestamp 1680363874
transform 1 0 3848 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_320
timestamp 1680363874
transform -1 0 3952 0 1 2370
box -8 -3 104 105
use FILL  FILL_5763
timestamp 1680363874
transform 1 0 3952 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_321
timestamp 1680363874
transform -1 0 4056 0 1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4565
timestamp 1680363874
transform 1 0 4084 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_322
timestamp 1680363874
transform -1 0 4152 0 1 2370
box -8 -3 104 105
use FILL  FILL_5764
timestamp 1680363874
transform 1 0 4152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5791
timestamp 1680363874
transform 1 0 4160 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4566
timestamp 1680363874
transform 1 0 4196 0 1 2375
box -3 -3 3 3
use INVX2  INVX2_370
timestamp 1680363874
transform 1 0 4168 0 1 2370
box -9 -3 26 105
use FILL  FILL_5792
timestamp 1680363874
transform 1 0 4184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5795
timestamp 1680363874
transform 1 0 4192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5797
timestamp 1680363874
transform 1 0 4200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5799
timestamp 1680363874
transform 1 0 4208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5801
timestamp 1680363874
transform 1 0 4216 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1680363874
transform -1 0 4248 0 1 2370
box -8 -3 32 105
use FILL  FILL_5802
timestamp 1680363874
transform 1 0 4248 0 1 2370
box -8 -3 16 105
use FILL  FILL_5803
timestamp 1680363874
transform 1 0 4256 0 1 2370
box -8 -3 16 105
use FILL  FILL_5804
timestamp 1680363874
transform 1 0 4264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5807
timestamp 1680363874
transform 1 0 4272 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4567
timestamp 1680363874
transform 1 0 4292 0 1 2375
box -3 -3 3 3
use FILL  FILL_5809
timestamp 1680363874
transform 1 0 4280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5811
timestamp 1680363874
transform 1 0 4288 0 1 2370
box -8 -3 16 105
use FILL  FILL_5813
timestamp 1680363874
transform 1 0 4296 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4568
timestamp 1680363874
transform 1 0 4316 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_192
timestamp 1680363874
transform 1 0 4304 0 1 2370
box -8 -3 46 105
use FILL  FILL_5815
timestamp 1680363874
transform 1 0 4344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5820
timestamp 1680363874
transform 1 0 4352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5821
timestamp 1680363874
transform 1 0 4360 0 1 2370
box -8 -3 16 105
use FILL  FILL_5822
timestamp 1680363874
transform 1 0 4368 0 1 2370
box -8 -3 16 105
use FILL  FILL_5823
timestamp 1680363874
transform 1 0 4376 0 1 2370
box -8 -3 16 105
use FILL  FILL_5825
timestamp 1680363874
transform 1 0 4384 0 1 2370
box -8 -3 16 105
use FILL  FILL_5827
timestamp 1680363874
transform 1 0 4392 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_252
timestamp 1680363874
transform 1 0 4400 0 1 2370
box -8 -3 46 105
use FILL  FILL_5829
timestamp 1680363874
transform 1 0 4440 0 1 2370
box -8 -3 16 105
use FILL  FILL_5830
timestamp 1680363874
transform 1 0 4448 0 1 2370
box -8 -3 16 105
use FILL  FILL_5831
timestamp 1680363874
transform 1 0 4456 0 1 2370
box -8 -3 16 105
use FILL  FILL_5832
timestamp 1680363874
transform 1 0 4464 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4569
timestamp 1680363874
transform 1 0 4492 0 1 2375
box -3 -3 3 3
use FILL  FILL_5833
timestamp 1680363874
transform 1 0 4472 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_193
timestamp 1680363874
transform -1 0 4520 0 1 2370
box -8 -3 46 105
use FILL  FILL_5834
timestamp 1680363874
transform 1 0 4520 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4570
timestamp 1680363874
transform 1 0 4540 0 1 2375
box -3 -3 3 3
use FILL  FILL_5839
timestamp 1680363874
transform 1 0 4528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5841
timestamp 1680363874
transform 1 0 4536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5843
timestamp 1680363874
transform 1 0 4544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5844
timestamp 1680363874
transform 1 0 4552 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_253
timestamp 1680363874
transform -1 0 4600 0 1 2370
box -8 -3 46 105
use FILL  FILL_5845
timestamp 1680363874
transform 1 0 4600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5849
timestamp 1680363874
transform 1 0 4608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5851
timestamp 1680363874
transform 1 0 4616 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_57
timestamp 1680363874
transform 1 0 4624 0 1 2370
box -8 -3 32 105
use FILL  FILL_5853
timestamp 1680363874
transform 1 0 4648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5854
timestamp 1680363874
transform 1 0 4656 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4571
timestamp 1680363874
transform 1 0 4676 0 1 2375
box -3 -3 3 3
use FILL  FILL_5855
timestamp 1680363874
transform 1 0 4664 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_373
timestamp 1680363874
transform 1 0 4672 0 1 2370
box -9 -3 26 105
use FILL  FILL_5857
timestamp 1680363874
transform 1 0 4688 0 1 2370
box -8 -3 16 105
use FILL  FILL_5858
timestamp 1680363874
transform 1 0 4696 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4572
timestamp 1680363874
transform 1 0 4716 0 1 2375
box -3 -3 3 3
use FILL  FILL_5859
timestamp 1680363874
transform 1 0 4704 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_195
timestamp 1680363874
transform 1 0 4712 0 1 2370
box -8 -3 46 105
use FILL  FILL_5860
timestamp 1680363874
transform 1 0 4752 0 1 2370
box -8 -3 16 105
use FILL  FILL_5861
timestamp 1680363874
transform 1 0 4760 0 1 2370
box -8 -3 16 105
use FILL  FILL_5862
timestamp 1680363874
transform 1 0 4768 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_374
timestamp 1680363874
transform 1 0 4776 0 1 2370
box -9 -3 26 105
use FILL  FILL_5863
timestamp 1680363874
transform 1 0 4792 0 1 2370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_47
timestamp 1680363874
transform 1 0 4827 0 1 2370
box -10 -3 10 3
use M2_M1  M2_M1_5183
timestamp 1680363874
transform 1 0 92 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1680363874
transform 1 0 116 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4636
timestamp 1680363874
transform 1 0 124 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5198
timestamp 1680363874
transform 1 0 124 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_4721
timestamp 1680363874
transform 1 0 116 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5184
timestamp 1680363874
transform 1 0 140 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4690
timestamp 1680363874
transform 1 0 140 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1680363874
transform 1 0 156 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5185
timestamp 1680363874
transform 1 0 156 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4604
timestamp 1680363874
transform 1 0 196 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5014
timestamp 1680363874
transform 1 0 204 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4605
timestamp 1680363874
transform 1 0 276 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5023
timestamp 1680363874
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1680363874
transform 1 0 180 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4615
timestamp 1680363874
transform 1 0 300 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1680363874
transform 1 0 324 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5024
timestamp 1680363874
transform 1 0 316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1680363874
transform 1 0 292 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1680363874
transform 1 0 300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1680363874
transform 1 0 188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1680363874
transform 1 0 172 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_4722
timestamp 1680363874
transform 1 0 180 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1680363874
transform 1 0 204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1680363874
transform 1 0 300 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1680363874
transform 1 0 260 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1680363874
transform 1 0 300 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5093
timestamp 1680363874
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1680363874
transform 1 0 324 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4724
timestamp 1680363874
transform 1 0 324 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5025
timestamp 1680363874
transform 1 0 348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1680363874
transform 1 0 356 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4607
timestamp 1680363874
transform 1 0 372 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5094
timestamp 1680363874
transform 1 0 364 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4693
timestamp 1680363874
transform 1 0 356 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1680363874
transform 1 0 364 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5015
timestamp 1680363874
transform 1 0 388 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4616
timestamp 1680363874
transform 1 0 484 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5095
timestamp 1680363874
transform 1 0 476 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1680363874
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1680363874
transform 1 0 492 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4694
timestamp 1680363874
transform 1 0 380 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1680363874
transform 1 0 436 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1680363874
transform 1 0 476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1680363874
transform 1 0 420 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5027
timestamp 1680363874
transform 1 0 516 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4638
timestamp 1680363874
transform 1 0 516 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1680363874
transform 1 0 508 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5098
timestamp 1680363874
transform 1 0 532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1680363874
transform 1 0 548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1680363874
transform 1 0 556 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4639
timestamp 1680363874
transform 1 0 548 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1680363874
transform 1 0 556 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1680363874
transform 1 0 580 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1680363874
transform 1 0 572 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1680363874
transform 1 0 748 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1680363874
transform 1 0 636 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5016
timestamp 1680363874
transform 1 0 644 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1680363874
transform 1 0 604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1680363874
transform 1 0 620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1680363874
transform 1 0 636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1680363874
transform 1 0 748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1680363874
transform 1 0 588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1680363874
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1680363874
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1680363874
transform 1 0 628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1680363874
transform 1 0 732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1680363874
transform 1 0 740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1680363874
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4697
timestamp 1680363874
transform 1 0 636 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1680363874
transform 1 0 740 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1680363874
transform 1 0 700 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5106
timestamp 1680363874
transform 1 0 772 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4699
timestamp 1680363874
transform 1 0 764 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1680363874
transform 1 0 756 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5107
timestamp 1680363874
transform 1 0 844 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4640
timestamp 1680363874
transform 1 0 852 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1680363874
transform 1 0 876 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5017
timestamp 1680363874
transform 1 0 900 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4610
timestamp 1680363874
transform 1 0 948 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1680363874
transform 1 0 988 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1680363874
transform 1 0 996 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5034
timestamp 1680363874
transform 1 0 1004 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1680363874
transform 1 0 988 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1680363874
transform 1 0 996 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1680363874
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4700
timestamp 1680363874
transform 1 0 1020 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5035
timestamp 1680363874
transform 1 0 1036 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4612
timestamp 1680363874
transform 1 0 1068 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5036
timestamp 1680363874
transform 1 0 1068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1680363874
transform 1 0 1060 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4641
timestamp 1680363874
transform 1 0 1068 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5112
timestamp 1680363874
transform 1 0 1076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1680363874
transform 1 0 1068 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4701
timestamp 1680363874
transform 1 0 1060 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1680363874
transform 1 0 1092 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1680363874
transform 1 0 1108 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5113
timestamp 1680363874
transform 1 0 1148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1680363874
transform 1 0 1156 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4703
timestamp 1680363874
transform 1 0 1148 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5190
timestamp 1680363874
transform 1 0 1188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1680363874
transform 1 0 1228 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4573
timestamp 1680363874
transform 1 0 1252 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5191
timestamp 1680363874
transform 1 0 1244 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1680363874
transform 1 0 1228 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1680363874
transform 1 0 1236 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_4704
timestamp 1680363874
transform 1 0 1244 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1680363874
transform 1 0 1228 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5037
timestamp 1680363874
transform 1 0 1324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1680363874
transform 1 0 1316 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4642
timestamp 1680363874
transform 1 0 1324 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5116
timestamp 1680363874
transform 1 0 1332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1680363874
transform 1 0 1348 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4619
timestamp 1680363874
transform 1 0 1396 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5118
timestamp 1680363874
transform 1 0 1396 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4574
timestamp 1680363874
transform 1 0 1428 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1680363874
transform 1 0 1532 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1680363874
transform 1 0 1452 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5038
timestamp 1680363874
transform 1 0 1524 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4643
timestamp 1680363874
transform 1 0 1460 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5119
timestamp 1680363874
transform 1 0 1476 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4585
timestamp 1680363874
transform 1 0 1596 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5039
timestamp 1680363874
transform 1 0 1596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1680363874
transform 1 0 1620 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4705
timestamp 1680363874
transform 1 0 1588 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1680363874
transform 1 0 1620 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5121
timestamp 1680363874
transform 1 0 1684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4575
timestamp 1680363874
transform 1 0 1708 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5012
timestamp 1680363874
transform 1 0 1700 0 1 2355
box -2 -2 2 2
use M3_M2  M3_M2_4586
timestamp 1680363874
transform 1 0 1708 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5192
timestamp 1680363874
transform 1 0 1716 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4707
timestamp 1680363874
transform 1 0 1716 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5013
timestamp 1680363874
transform 1 0 1732 0 1 2355
box -2 -2 2 2
use M3_M2  M3_M2_4587
timestamp 1680363874
transform 1 0 1812 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1680363874
transform 1 0 1868 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1680363874
transform 1 0 1860 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1680363874
transform 1 0 1908 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5122
timestamp 1680363874
transform 1 0 1908 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1680363874
transform 1 0 1908 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4644
timestamp 1680363874
transform 1 0 1948 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1680363874
transform 1 0 1972 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5202
timestamp 1680363874
transform 1 0 1964 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1680363874
transform 1 0 1980 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4645
timestamp 1680363874
transform 1 0 1980 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5123
timestamp 1680363874
transform 1 0 2028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1680363874
transform 1 0 2060 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4666
timestamp 1680363874
transform 1 0 2012 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1680363874
transform 1 0 2028 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1680363874
transform 1 0 2092 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5088
timestamp 1680363874
transform 1 0 2092 0 1 2333
box -2 -2 2 2
use M3_M2  M3_M2_4622
timestamp 1680363874
transform 1 0 2116 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1680363874
transform 1 0 2140 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5125
timestamp 1680363874
transform 1 0 2140 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4646
timestamp 1680363874
transform 1 0 2164 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1680363874
transform 1 0 2108 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5041
timestamp 1680363874
transform 1 0 2220 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4576
timestamp 1680363874
transform 1 0 2236 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1680363874
transform 1 0 2260 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5126
timestamp 1680363874
transform 1 0 2228 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4624
timestamp 1680363874
transform 1 0 2244 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5042
timestamp 1680363874
transform 1 0 2252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1680363874
transform 1 0 2268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1680363874
transform 1 0 2244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1680363874
transform 1 0 2260 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4667
timestamp 1680363874
transform 1 0 2244 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5129
timestamp 1680363874
transform 1 0 2284 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4591
timestamp 1680363874
transform 1 0 2316 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5044
timestamp 1680363874
transform 1 0 2324 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4592
timestamp 1680363874
transform 1 0 2420 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5045
timestamp 1680363874
transform 1 0 2412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1680363874
transform 1 0 2348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1680363874
transform 1 0 2404 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4647
timestamp 1680363874
transform 1 0 2412 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5046
timestamp 1680363874
transform 1 0 2500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1680363874
transform 1 0 2516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1680363874
transform 1 0 2524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1680363874
transform 1 0 2492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1680363874
transform 1 0 2508 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4668
timestamp 1680363874
transform 1 0 2492 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1680363874
transform 1 0 2508 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5134
timestamp 1680363874
transform 1 0 2532 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4669
timestamp 1680363874
transform 1 0 2532 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5049
timestamp 1680363874
transform 1 0 2548 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4648
timestamp 1680363874
transform 1 0 2564 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1680363874
transform 1 0 2556 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1680363874
transform 1 0 2604 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5050
timestamp 1680363874
transform 1 0 2604 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4625
timestamp 1680363874
transform 1 0 2612 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5051
timestamp 1680363874
transform 1 0 2620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1680363874
transform 1 0 2596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1680363874
transform 1 0 2612 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4670
timestamp 1680363874
transform 1 0 2612 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1680363874
transform 1 0 2628 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5137
timestamp 1680363874
transform 1 0 2636 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4671
timestamp 1680363874
transform 1 0 2636 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5052
timestamp 1680363874
transform 1 0 2676 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4594
timestamp 1680363874
transform 1 0 2692 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5194
timestamp 1680363874
transform 1 0 2732 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4595
timestamp 1680363874
transform 1 0 2764 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5138
timestamp 1680363874
transform 1 0 2852 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4672
timestamp 1680363874
transform 1 0 2852 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5195
timestamp 1680363874
transform 1 0 2860 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1680363874
transform 1 0 2884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1680363874
transform 1 0 2900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1680363874
transform 1 0 2916 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4673
timestamp 1680363874
transform 1 0 2908 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5054
timestamp 1680363874
transform 1 0 2932 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4732
timestamp 1680363874
transform 1 0 2956 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5140
timestamp 1680363874
transform 1 0 2972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1680363874
transform 1 0 3004 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1680363874
transform 1 0 3108 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4627
timestamp 1680363874
transform 1 0 3116 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5141
timestamp 1680363874
transform 1 0 3124 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4674
timestamp 1680363874
transform 1 0 3116 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1680363874
transform 1 0 3140 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5142
timestamp 1680363874
transform 1 0 3140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1680363874
transform 1 0 3204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1680363874
transform 1 0 3236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1680363874
transform 1 0 3268 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4649
timestamp 1680363874
transform 1 0 3260 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5058
timestamp 1680363874
transform 1 0 3300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1680363874
transform 1 0 3292 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4650
timestamp 1680363874
transform 1 0 3300 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5144
timestamp 1680363874
transform 1 0 3316 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4675
timestamp 1680363874
transform 1 0 3316 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1680363874
transform 1 0 3316 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5059
timestamp 1680363874
transform 1 0 3340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1680363874
transform 1 0 3364 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4711
timestamp 1680363874
transform 1 0 3356 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1680363874
transform 1 0 3388 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5060
timestamp 1680363874
transform 1 0 3404 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4629
timestamp 1680363874
transform 1 0 3484 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5145
timestamp 1680363874
transform 1 0 3444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1680363874
transform 1 0 3484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1680363874
transform 1 0 3492 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4676
timestamp 1680363874
transform 1 0 3444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1680363874
transform 1 0 3492 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1680363874
transform 1 0 3484 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1680363874
transform 1 0 3532 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5061
timestamp 1680363874
transform 1 0 3532 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4651
timestamp 1680363874
transform 1 0 3532 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1680363874
transform 1 0 3548 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5148
timestamp 1680363874
transform 1 0 3556 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4597
timestamp 1680363874
transform 1 0 3588 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5062
timestamp 1680363874
transform 1 0 3580 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4652
timestamp 1680363874
transform 1 0 3580 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5149
timestamp 1680363874
transform 1 0 3588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1680363874
transform 1 0 3628 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1680363874
transform 1 0 3620 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4631
timestamp 1680363874
transform 1 0 3628 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5150
timestamp 1680363874
transform 1 0 3636 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4678
timestamp 1680363874
transform 1 0 3652 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5151
timestamp 1680363874
transform 1 0 3668 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4734
timestamp 1680363874
transform 1 0 3668 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5064
timestamp 1680363874
transform 1 0 3684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1680363874
transform 1 0 3692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1680363874
transform 1 0 3708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1680363874
transform 1 0 3676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1680363874
transform 1 0 3700 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4653
timestamp 1680363874
transform 1 0 3708 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5154
timestamp 1680363874
transform 1 0 3716 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4713
timestamp 1680363874
transform 1 0 3692 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1680363874
transform 1 0 3708 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1680363874
transform 1 0 3716 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5155
timestamp 1680363874
transform 1 0 3732 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4715
timestamp 1680363874
transform 1 0 3732 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5067
timestamp 1680363874
transform 1 0 3756 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4716
timestamp 1680363874
transform 1 0 3756 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1680363874
transform 1 0 3804 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5068
timestamp 1680363874
transform 1 0 3828 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4599
timestamp 1680363874
transform 1 0 3836 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5069
timestamp 1680363874
transform 1 0 3836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1680363874
transform 1 0 3804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1680363874
transform 1 0 3820 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4654
timestamp 1680363874
transform 1 0 3828 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5158
timestamp 1680363874
transform 1 0 3836 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4679
timestamp 1680363874
transform 1 0 3820 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1680363874
transform 1 0 3892 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1680363874
transform 1 0 3892 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1680363874
transform 1 0 3908 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1680363874
transform 1 0 3908 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1680363874
transform 1 0 3964 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5021
timestamp 1680363874
transform 1 0 3964 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1680363874
transform 1 0 3956 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4657
timestamp 1680363874
transform 1 0 3964 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1680363874
transform 1 0 3956 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1680363874
transform 1 0 3956 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1680363874
transform 1 0 3988 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5071
timestamp 1680363874
transform 1 0 3988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1680363874
transform 1 0 4004 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1680363874
transform 1 0 3980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1680363874
transform 1 0 3996 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4658
timestamp 1680363874
transform 1 0 4004 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1680363874
transform 1 0 3980 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1680363874
transform 1 0 4020 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5073
timestamp 1680363874
transform 1 0 4036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1680363874
transform 1 0 4028 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4737
timestamp 1680363874
transform 1 0 4028 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1680363874
transform 1 0 4044 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1680363874
transform 1 0 4068 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5162
timestamp 1680363874
transform 1 0 4068 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1680363874
transform 1 0 4108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1680363874
transform 1 0 4116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1680363874
transform 1 0 4100 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4682
timestamp 1680363874
transform 1 0 4092 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1680363874
transform 1 0 4108 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1680363874
transform 1 0 4132 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5164
timestamp 1680363874
transform 1 0 4124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1680363874
transform 1 0 4140 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4683
timestamp 1680363874
transform 1 0 4196 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1680363874
transform 1 0 4236 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5076
timestamp 1680363874
transform 1 0 4236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1680363874
transform 1 0 4252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1680363874
transform 1 0 4220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1680363874
transform 1 0 4228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1680363874
transform 1 0 4244 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4684
timestamp 1680363874
transform 1 0 4220 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1680363874
transform 1 0 4252 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1680363874
transform 1 0 4252 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1680363874
transform 1 0 4244 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5169
timestamp 1680363874
transform 1 0 4284 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4719
timestamp 1680363874
transform 1 0 4292 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5078
timestamp 1680363874
transform 1 0 4316 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4579
timestamp 1680363874
transform 1 0 4340 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1680363874
transform 1 0 4332 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5079
timestamp 1680363874
transform 1 0 4332 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4661
timestamp 1680363874
transform 1 0 4332 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1680363874
transform 1 0 4348 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5022
timestamp 1680363874
transform 1 0 4356 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1680363874
transform 1 0 4356 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4686
timestamp 1680363874
transform 1 0 4356 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1680363874
transform 1 0 4364 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1680363874
transform 1 0 4452 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1680363874
transform 1 0 4484 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1680363874
transform 1 0 4428 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1680363874
transform 1 0 4444 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5080
timestamp 1680363874
transform 1 0 4508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1680363874
transform 1 0 4420 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1680363874
transform 1 0 4428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1680363874
transform 1 0 4468 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4687
timestamp 1680363874
transform 1 0 4468 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5081
timestamp 1680363874
transform 1 0 4548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1680363874
transform 1 0 4564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1680363874
transform 1 0 4556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1680363874
transform 1 0 4572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1680363874
transform 1 0 4588 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4662
timestamp 1680363874
transform 1 0 4588 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5176
timestamp 1680363874
transform 1 0 4620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1680363874
transform 1 0 4636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1680363874
transform 1 0 4652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1680363874
transform 1 0 4660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1680363874
transform 1 0 4644 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4663
timestamp 1680363874
transform 1 0 4652 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5178
timestamp 1680363874
transform 1 0 4660 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4720
timestamp 1680363874
transform 1 0 4636 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5087
timestamp 1680363874
transform 1 0 4788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1680363874
transform 1 0 4692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1680363874
transform 1 0 4700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1680363874
transform 1 0 4708 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4664
timestamp 1680363874
transform 1 0 4716 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5182
timestamp 1680363874
transform 1 0 4756 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4688
timestamp 1680363874
transform 1 0 4700 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1680363874
transform 1 0 4756 0 1 2315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_48
timestamp 1680363874
transform 1 0 24 0 1 2270
box -10 -3 10 3
use M3_M2  M3_M2_4744
timestamp 1680363874
transform 1 0 84 0 1 2275
box -3 -3 3 3
use FILL  FILL_5281
timestamp 1680363874
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1680363874
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1680363874
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_17
timestamp 1680363874
transform -1 0 128 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5289
timestamp 1680363874
transform 1 0 128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1680363874
transform 1 0 136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1680363874
transform 1 0 144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1680363874
transform 1 0 152 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_19
timestamp 1680363874
transform -1 0 192 0 -1 2370
box -8 -3 40 105
use FAX1  FAX1_9
timestamp 1680363874
transform -1 0 312 0 -1 2370
box -5 -3 126 105
use FILL  FILL_5323
timestamp 1680363874
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_128
timestamp 1680363874
transform -1 0 352 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5324
timestamp 1680363874
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1680363874
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1680363874
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FAX1  FAX1_10
timestamp 1680363874
transform -1 0 496 0 -1 2370
box -5 -3 126 105
use FILL  FILL_5327
timestamp 1680363874
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1680363874
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1680363874
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1680363874
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1680363874
transform 1 0 528 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_350
timestamp 1680363874
transform -1 0 552 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5337
timestamp 1680363874
transform 1 0 552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1680363874
transform 1 0 560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1680363874
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_353
timestamp 1680363874
transform 1 0 576 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_181
timestamp 1680363874
transform 1 0 592 0 -1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4745
timestamp 1680363874
transform 1 0 692 0 1 2275
box -3 -3 3 3
use FAX1  FAX1_11
timestamp 1680363874
transform -1 0 752 0 -1 2370
box -5 -3 126 105
use FILL  FILL_5357
timestamp 1680363874
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1680363874
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1680363874
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1680363874
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1680363874
transform 1 0 784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5367
timestamp 1680363874
transform 1 0 792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1680363874
transform 1 0 800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1680363874
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1680363874
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1680363874
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1680363874
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5376
timestamp 1680363874
transform 1 0 840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5378
timestamp 1680363874
transform 1 0 848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5380
timestamp 1680363874
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5382
timestamp 1680363874
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5393
timestamp 1680363874
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5394
timestamp 1680363874
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FAX1  FAX1_12
timestamp 1680363874
transform -1 0 1008 0 -1 2370
box -5 -3 126 105
use FILL  FILL_5395
timestamp 1680363874
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5397
timestamp 1680363874
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5399
timestamp 1680363874
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5402
timestamp 1680363874
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use AND2X2  AND2X2_18
timestamp 1680363874
transform -1 0 1072 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5403
timestamp 1680363874
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5405
timestamp 1680363874
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5408
timestamp 1680363874
transform 1 0 1088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5409
timestamp 1680363874
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5410
timestamp 1680363874
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5411
timestamp 1680363874
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5416
timestamp 1680363874
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1680363874
transform -1 0 1160 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5417
timestamp 1680363874
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5418
timestamp 1680363874
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5419
timestamp 1680363874
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5421
timestamp 1680363874
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5423
timestamp 1680363874
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5425
timestamp 1680363874
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4746
timestamp 1680363874
transform 1 0 1220 0 1 2275
box -3 -3 3 3
use FILL  FILL_5427
timestamp 1680363874
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_22
timestamp 1680363874
transform 1 0 1216 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5436
timestamp 1680363874
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5437
timestamp 1680363874
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5438
timestamp 1680363874
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5439
timestamp 1680363874
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5440
timestamp 1680363874
transform 1 0 1280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5441
timestamp 1680363874
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5442
timestamp 1680363874
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5443
timestamp 1680363874
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4747
timestamp 1680363874
transform 1 0 1332 0 1 2275
box -3 -3 3 3
use AOI22X1  AOI22X1_183
timestamp 1680363874
transform 1 0 1312 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5444
timestamp 1680363874
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5445
timestamp 1680363874
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5446
timestamp 1680363874
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5447
timestamp 1680363874
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5448
timestamp 1680363874
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_356
timestamp 1680363874
transform -1 0 1408 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5449
timestamp 1680363874
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5451
timestamp 1680363874
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5466
timestamp 1680363874
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5467
timestamp 1680363874
transform 1 0 1432 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_308
timestamp 1680363874
transform -1 0 1536 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5468
timestamp 1680363874
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5469
timestamp 1680363874
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5470
timestamp 1680363874
transform 1 0 1552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5471
timestamp 1680363874
transform 1 0 1560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5472
timestamp 1680363874
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5473
timestamp 1680363874
transform 1 0 1576 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_309
timestamp 1680363874
transform 1 0 1584 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5474
timestamp 1680363874
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5476
timestamp 1680363874
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5478
timestamp 1680363874
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5479
timestamp 1680363874
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5480
timestamp 1680363874
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5481
timestamp 1680363874
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5482
timestamp 1680363874
transform 1 0 1728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5483
timestamp 1680363874
transform 1 0 1736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5484
timestamp 1680363874
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5485
timestamp 1680363874
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5486
timestamp 1680363874
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5487
timestamp 1680363874
transform 1 0 1768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5488
timestamp 1680363874
transform 1 0 1776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5489
timestamp 1680363874
transform 1 0 1784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5490
timestamp 1680363874
transform 1 0 1792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5492
timestamp 1680363874
transform 1 0 1800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5494
timestamp 1680363874
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5497
timestamp 1680363874
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5498
timestamp 1680363874
transform 1 0 1824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5499
timestamp 1680363874
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5500
timestamp 1680363874
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5501
timestamp 1680363874
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5502
timestamp 1680363874
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5504
timestamp 1680363874
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5506
timestamp 1680363874
transform 1 0 1872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5511
timestamp 1680363874
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_25
timestamp 1680363874
transform -1 0 1920 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5512
timestamp 1680363874
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5513
timestamp 1680363874
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5514
timestamp 1680363874
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5516
timestamp 1680363874
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5518
timestamp 1680363874
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5520
timestamp 1680363874
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_311
timestamp 1680363874
transform 1 0 1968 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5541
timestamp 1680363874
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5542
timestamp 1680363874
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_312
timestamp 1680363874
transform 1 0 2080 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_358
timestamp 1680363874
transform 1 0 2176 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5543
timestamp 1680363874
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5545
timestamp 1680363874
transform 1 0 2200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5547
timestamp 1680363874
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5549
timestamp 1680363874
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5552
timestamp 1680363874
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_245
timestamp 1680363874
transform -1 0 2272 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5553
timestamp 1680363874
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5555
timestamp 1680363874
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5557
timestamp 1680363874
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5559
timestamp 1680363874
transform 1 0 2296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5562
timestamp 1680363874
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_314
timestamp 1680363874
transform 1 0 2312 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5563
timestamp 1680363874
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5564
timestamp 1680363874
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5565
timestamp 1680363874
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5566
timestamp 1680363874
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5567
timestamp 1680363874
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5569
timestamp 1680363874
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5571
timestamp 1680363874
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5573
timestamp 1680363874
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5575
timestamp 1680363874
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_247
timestamp 1680363874
transform 1 0 2480 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5577
timestamp 1680363874
transform 1 0 2520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5579
timestamp 1680363874
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5581
timestamp 1680363874
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5583
timestamp 1680363874
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5585
timestamp 1680363874
transform 1 0 2552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5587
timestamp 1680363874
transform 1 0 2560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5589
timestamp 1680363874
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5591
timestamp 1680363874
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_248
timestamp 1680363874
transform 1 0 2584 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5598
timestamp 1680363874
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5600
timestamp 1680363874
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5602
timestamp 1680363874
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5606
timestamp 1680363874
transform 1 0 2648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5607
timestamp 1680363874
transform 1 0 2656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5608
timestamp 1680363874
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5609
timestamp 1680363874
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5610
timestamp 1680363874
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_361
timestamp 1680363874
transform 1 0 2688 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5611
timestamp 1680363874
transform 1 0 2704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5612
timestamp 1680363874
transform 1 0 2712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5613
timestamp 1680363874
transform 1 0 2720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5614
timestamp 1680363874
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4748
timestamp 1680363874
transform 1 0 2748 0 1 2275
box -3 -3 3 3
use FILL  FILL_5615
timestamp 1680363874
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5616
timestamp 1680363874
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5617
timestamp 1680363874
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5618
timestamp 1680363874
transform 1 0 2760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5619
timestamp 1680363874
transform 1 0 2768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5620
timestamp 1680363874
transform 1 0 2776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5621
timestamp 1680363874
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5622
timestamp 1680363874
transform 1 0 2792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5623
timestamp 1680363874
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5624
timestamp 1680363874
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5625
timestamp 1680363874
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5626
timestamp 1680363874
transform 1 0 2824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5627
timestamp 1680363874
transform 1 0 2832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5628
timestamp 1680363874
transform 1 0 2840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5632
timestamp 1680363874
transform 1 0 2848 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_41
timestamp 1680363874
transform -1 0 2880 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5633
timestamp 1680363874
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5635
timestamp 1680363874
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5637
timestamp 1680363874
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5640
timestamp 1680363874
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_364
timestamp 1680363874
transform 1 0 2912 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5641
timestamp 1680363874
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5643
timestamp 1680363874
transform 1 0 2936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5645
timestamp 1680363874
transform 1 0 2944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5647
timestamp 1680363874
transform 1 0 2952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5649
timestamp 1680363874
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5652
timestamp 1680363874
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_132
timestamp 1680363874
transform 1 0 2976 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5653
timestamp 1680363874
transform 1 0 3008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5655
timestamp 1680363874
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5657
timestamp 1680363874
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5659
timestamp 1680363874
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5661
timestamp 1680363874
transform 1 0 3040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5662
timestamp 1680363874
transform 1 0 3048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5663
timestamp 1680363874
transform 1 0 3056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5664
timestamp 1680363874
transform 1 0 3064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5665
timestamp 1680363874
transform 1 0 3072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5666
timestamp 1680363874
transform 1 0 3080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5667
timestamp 1680363874
transform 1 0 3088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5668
timestamp 1680363874
transform 1 0 3096 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_133
timestamp 1680363874
transform -1 0 3136 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5669
timestamp 1680363874
transform 1 0 3136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5671
timestamp 1680363874
transform 1 0 3144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5673
timestamp 1680363874
transform 1 0 3152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5679
timestamp 1680363874
transform 1 0 3160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5680
timestamp 1680363874
transform 1 0 3168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5681
timestamp 1680363874
transform 1 0 3176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5682
timestamp 1680363874
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5683
timestamp 1680363874
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_51
timestamp 1680363874
transform -1 0 3224 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5684
timestamp 1680363874
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5685
timestamp 1680363874
transform 1 0 3232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5686
timestamp 1680363874
transform 1 0 3240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5687
timestamp 1680363874
transform 1 0 3248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5688
timestamp 1680363874
transform 1 0 3256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5689
timestamp 1680363874
transform 1 0 3264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5690
timestamp 1680363874
transform 1 0 3272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5691
timestamp 1680363874
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_365
timestamp 1680363874
transform -1 0 3304 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5692
timestamp 1680363874
transform 1 0 3304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5693
timestamp 1680363874
transform 1 0 3312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5694
timestamp 1680363874
transform 1 0 3320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5696
timestamp 1680363874
transform 1 0 3328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5701
timestamp 1680363874
transform 1 0 3336 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_53
timestamp 1680363874
transform -1 0 3368 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5702
timestamp 1680363874
transform 1 0 3368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5703
timestamp 1680363874
transform 1 0 3376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5704
timestamp 1680363874
transform 1 0 3384 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_319
timestamp 1680363874
transform 1 0 3392 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5710
timestamp 1680363874
transform 1 0 3488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5711
timestamp 1680363874
transform 1 0 3496 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_366
timestamp 1680363874
transform -1 0 3520 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5712
timestamp 1680363874
transform 1 0 3520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5715
timestamp 1680363874
transform 1 0 3528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5716
timestamp 1680363874
transform 1 0 3536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5717
timestamp 1680363874
transform 1 0 3544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5718
timestamp 1680363874
transform 1 0 3552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5720
timestamp 1680363874
transform 1 0 3560 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_186
timestamp 1680363874
transform 1 0 3568 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5723
timestamp 1680363874
transform 1 0 3608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5724
timestamp 1680363874
transform 1 0 3616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5726
timestamp 1680363874
transform 1 0 3624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5728
timestamp 1680363874
transform 1 0 3632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5730
timestamp 1680363874
transform 1 0 3640 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4749
timestamp 1680363874
transform 1 0 3660 0 1 2275
box -3 -3 3 3
use FILL  FILL_5732
timestamp 1680363874
transform 1 0 3648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5734
timestamp 1680363874
transform 1 0 3656 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_369
timestamp 1680363874
transform 1 0 3664 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_187
timestamp 1680363874
transform -1 0 3720 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5743
timestamp 1680363874
transform 1 0 3720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5744
timestamp 1680363874
transform 1 0 3728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5745
timestamp 1680363874
transform 1 0 3736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5747
timestamp 1680363874
transform 1 0 3744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5749
timestamp 1680363874
transform 1 0 3752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5751
timestamp 1680363874
transform 1 0 3760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5753
timestamp 1680363874
transform 1 0 3768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5755
timestamp 1680363874
transform 1 0 3776 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_189
timestamp 1680363874
transform 1 0 3784 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5758
timestamp 1680363874
transform 1 0 3824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5759
timestamp 1680363874
transform 1 0 3832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5761
timestamp 1680363874
transform 1 0 3840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5765
timestamp 1680363874
transform 1 0 3848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5766
timestamp 1680363874
transform 1 0 3856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5767
timestamp 1680363874
transform 1 0 3864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5768
timestamp 1680363874
transform 1 0 3872 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_54
timestamp 1680363874
transform -1 0 3904 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5769
timestamp 1680363874
transform 1 0 3904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5770
timestamp 1680363874
transform 1 0 3912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5771
timestamp 1680363874
transform 1 0 3920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5772
timestamp 1680363874
transform 1 0 3928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5773
timestamp 1680363874
transform 1 0 3936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5774
timestamp 1680363874
transform 1 0 3944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5775
timestamp 1680363874
transform 1 0 3952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5776
timestamp 1680363874
transform 1 0 3960 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_251
timestamp 1680363874
transform 1 0 3968 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5777
timestamp 1680363874
transform 1 0 4008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5778
timestamp 1680363874
transform 1 0 4016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5779
timestamp 1680363874
transform 1 0 4024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5780
timestamp 1680363874
transform 1 0 4032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5781
timestamp 1680363874
transform 1 0 4040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5782
timestamp 1680363874
transform 1 0 4048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5783
timestamp 1680363874
transform 1 0 4056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5784
timestamp 1680363874
transform 1 0 4064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5785
timestamp 1680363874
transform 1 0 4072 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_190
timestamp 1680363874
transform -1 0 4120 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5786
timestamp 1680363874
transform 1 0 4120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5787
timestamp 1680363874
transform 1 0 4128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5788
timestamp 1680363874
transform 1 0 4136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5789
timestamp 1680363874
transform 1 0 4144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5790
timestamp 1680363874
transform 1 0 4152 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4750
timestamp 1680363874
transform 1 0 4180 0 1 2275
box -3 -3 3 3
use INVX2  INVX2_371
timestamp 1680363874
transform 1 0 4160 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5793
timestamp 1680363874
transform 1 0 4176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5794
timestamp 1680363874
transform 1 0 4184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5796
timestamp 1680363874
transform 1 0 4192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5798
timestamp 1680363874
transform 1 0 4200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5800
timestamp 1680363874
transform 1 0 4208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5805
timestamp 1680363874
transform 1 0 4216 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_191
timestamp 1680363874
transform 1 0 4224 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5806
timestamp 1680363874
transform 1 0 4264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5808
timestamp 1680363874
transform 1 0 4272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5810
timestamp 1680363874
transform 1 0 4280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5812
timestamp 1680363874
transform 1 0 4288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5814
timestamp 1680363874
transform 1 0 4296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5816
timestamp 1680363874
transform 1 0 4304 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_372
timestamp 1680363874
transform 1 0 4312 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5817
timestamp 1680363874
transform 1 0 4328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5818
timestamp 1680363874
transform 1 0 4336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5819
timestamp 1680363874
transform 1 0 4344 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_56
timestamp 1680363874
transform 1 0 4352 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5824
timestamp 1680363874
transform 1 0 4376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5826
timestamp 1680363874
transform 1 0 4384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5828
timestamp 1680363874
transform 1 0 4392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5835
timestamp 1680363874
transform 1 0 4400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5836
timestamp 1680363874
transform 1 0 4408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5837
timestamp 1680363874
transform 1 0 4416 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_323
timestamp 1680363874
transform -1 0 4520 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5838
timestamp 1680363874
transform 1 0 4520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5840
timestamp 1680363874
transform 1 0 4528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5842
timestamp 1680363874
transform 1 0 4536 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_254
timestamp 1680363874
transform 1 0 4544 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5846
timestamp 1680363874
transform 1 0 4584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5847
timestamp 1680363874
transform 1 0 4592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5848
timestamp 1680363874
transform 1 0 4600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5850
timestamp 1680363874
transform 1 0 4608 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4751
timestamp 1680363874
transform 1 0 4628 0 1 2275
box -3 -3 3 3
use FILL  FILL_5852
timestamp 1680363874
transform 1 0 4616 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_194
timestamp 1680363874
transform 1 0 4624 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5856
timestamp 1680363874
transform 1 0 4664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5864
timestamp 1680363874
transform 1 0 4672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5865
timestamp 1680363874
transform 1 0 4680 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_375
timestamp 1680363874
transform 1 0 4688 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_324
timestamp 1680363874
transform -1 0 4800 0 -1 2370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_49
timestamp 1680363874
transform 1 0 4851 0 1 2270
box -10 -3 10 3
use M2_M1  M2_M1_5324
timestamp 1680363874
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1680363874
transform 1 0 100 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4832
timestamp 1680363874
transform 1 0 108 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5203
timestamp 1680363874
transform 1 0 124 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1680363874
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1680363874
transform 1 0 108 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4843
timestamp 1680363874
transform 1 0 116 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5209
timestamp 1680363874
transform 1 0 140 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4844
timestamp 1680363874
transform 1 0 140 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1680363874
transform 1 0 148 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5204
timestamp 1680363874
transform 1 0 172 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1680363874
transform 1 0 180 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1680363874
transform 1 0 164 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4797
timestamp 1680363874
transform 1 0 196 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5211
timestamp 1680363874
transform 1 0 204 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1680363874
transform 1 0 244 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4754
timestamp 1680363874
transform 1 0 268 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5228
timestamp 1680363874
transform 1 0 260 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4845
timestamp 1680363874
transform 1 0 260 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5212
timestamp 1680363874
transform 1 0 300 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4833
timestamp 1680363874
transform 1 0 292 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5229
timestamp 1680363874
transform 1 0 332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1680363874
transform 1 0 324 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4886
timestamp 1680363874
transform 1 0 324 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1680363874
transform 1 0 364 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5230
timestamp 1680363874
transform 1 0 356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1680363874
transform 1 0 364 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4798
timestamp 1680363874
transform 1 0 372 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5326
timestamp 1680363874
transform 1 0 372 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4774
timestamp 1680363874
transform 1 0 428 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5213
timestamp 1680363874
transform 1 0 428 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4834
timestamp 1680363874
transform 1 0 428 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5327
timestamp 1680363874
transform 1 0 428 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1680363874
transform 1 0 420 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1680363874
transform 1 0 444 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4835
timestamp 1680363874
transform 1 0 484 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5232
timestamp 1680363874
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1680363874
transform 1 0 500 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4846
timestamp 1680363874
transform 1 0 556 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1680363874
transform 1 0 628 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1680363874
transform 1 0 716 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5233
timestamp 1680363874
transform 1 0 732 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4776
timestamp 1680363874
transform 1 0 780 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5234
timestamp 1680363874
transform 1 0 844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1680363874
transform 1 0 852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1680363874
transform 1 0 860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1680363874
transform 1 0 868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1680363874
transform 1 0 756 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4863
timestamp 1680363874
transform 1 0 820 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1680363874
transform 1 0 852 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1680363874
transform 1 0 836 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1680363874
transform 1 0 908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1680363874
transform 1 0 884 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5236
timestamp 1680363874
transform 1 0 908 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4888
timestamp 1680363874
transform 1 0 876 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1680363874
transform 1 0 948 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1680363874
transform 1 0 964 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1680363874
transform 1 0 956 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5331
timestamp 1680363874
transform 1 0 948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1680363874
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1680363874
transform 1 0 988 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1680363874
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4762
timestamp 1680363874
transform 1 0 1036 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5215
timestamp 1680363874
transform 1 0 1036 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4847
timestamp 1680363874
transform 1 0 1036 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5206
timestamp 1680363874
transform 1 0 1060 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4778
timestamp 1680363874
transform 1 0 1076 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5216
timestamp 1680363874
transform 1 0 1076 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4838
timestamp 1680363874
transform 1 0 1060 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1680363874
transform 1 0 1092 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1680363874
transform 1 0 1148 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5238
timestamp 1680363874
transform 1 0 1148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1680363874
transform 1 0 1196 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1680363874
transform 1 0 1276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1680363874
transform 1 0 1292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1680363874
transform 1 0 1308 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1680363874
transform 1 0 1300 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4802
timestamp 1680363874
transform 1 0 1332 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5241
timestamp 1680363874
transform 1 0 1332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1680363874
transform 1 0 1348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1680363874
transform 1 0 1388 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4865
timestamp 1680363874
transform 1 0 1412 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1680363874
transform 1 0 1428 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5244
timestamp 1680363874
transform 1 0 1460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1680363874
transform 1 0 1476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1680363874
transform 1 0 1428 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1680363874
transform 1 0 1436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1680363874
transform 1 0 1452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1680363874
transform 1 0 1468 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4866
timestamp 1680363874
transform 1 0 1436 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5338
timestamp 1680363874
transform 1 0 1524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1680363874
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4763
timestamp 1680363874
transform 1 0 1572 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1680363874
transform 1 0 1580 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1680363874
transform 1 0 1596 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5246
timestamp 1680363874
transform 1 0 1572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1680363874
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1680363874
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4867
timestamp 1680363874
transform 1 0 1564 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5340
timestamp 1680363874
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4805
timestamp 1680363874
transform 1 0 1612 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5249
timestamp 1680363874
transform 1 0 1612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1680363874
transform 1 0 1620 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4868
timestamp 1680363874
transform 1 0 1620 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5342
timestamp 1680363874
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4780
timestamp 1680363874
transform 1 0 1692 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1680363874
transform 1 0 1708 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5250
timestamp 1680363874
transform 1 0 1684 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1680363874
transform 1 0 1692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1680363874
transform 1 0 1708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1680363874
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1680363874
transform 1 0 1700 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1680363874
transform 1 0 1716 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4869
timestamp 1680363874
transform 1 0 1716 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1680363874
transform 1 0 1748 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5345
timestamp 1680363874
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1680363874
transform 1 0 1772 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4755
timestamp 1680363874
transform 1 0 1796 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1680363874
transform 1 0 1796 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1680363874
transform 1 0 1812 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5254
timestamp 1680363874
transform 1 0 1796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1680363874
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1680363874
transform 1 0 1788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1680363874
transform 1 0 1812 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4849
timestamp 1680363874
transform 1 0 1820 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5256
timestamp 1680363874
transform 1 0 1836 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4850
timestamp 1680363874
transform 1 0 1836 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5348
timestamp 1680363874
transform 1 0 1844 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4870
timestamp 1680363874
transform 1 0 1844 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1680363874
transform 1 0 1940 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1680363874
transform 1 0 1988 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5257
timestamp 1680363874
transform 1 0 1940 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1680363874
transform 1 0 1988 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1680363874
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4811
timestamp 1680363874
transform 1 0 2092 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5259
timestamp 1680363874
transform 1 0 2084 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4756
timestamp 1680363874
transform 1 0 2132 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1680363874
transform 1 0 2124 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5260
timestamp 1680363874
transform 1 0 2100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1680363874
transform 1 0 2116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1680363874
transform 1 0 2092 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4851
timestamp 1680363874
transform 1 0 2100 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5218
timestamp 1680363874
transform 1 0 2132 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1680363874
transform 1 0 2108 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1680363874
transform 1 0 2124 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4765
timestamp 1680363874
transform 1 0 2156 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5208
timestamp 1680363874
transform 1 0 2180 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4812
timestamp 1680363874
transform 1 0 2188 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5262
timestamp 1680363874
transform 1 0 2188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1680363874
transform 1 0 2228 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4871
timestamp 1680363874
transform 1 0 2220 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1680363874
transform 1 0 2268 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1680363874
transform 1 0 2260 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5263
timestamp 1680363874
transform 1 0 2244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1680363874
transform 1 0 2260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1680363874
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4852
timestamp 1680363874
transform 1 0 2260 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5354
timestamp 1680363874
transform 1 0 2268 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4782
timestamp 1680363874
transform 1 0 2284 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5265
timestamp 1680363874
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1680363874
transform 1 0 2340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1680363874
transform 1 0 2356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1680363874
transform 1 0 2308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1680363874
transform 1 0 2316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1680363874
transform 1 0 2332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1680363874
transform 1 0 2348 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4872
timestamp 1680363874
transform 1 0 2348 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5268
timestamp 1680363874
transform 1 0 2412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1680363874
transform 1 0 2404 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4873
timestamp 1680363874
transform 1 0 2412 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5269
timestamp 1680363874
transform 1 0 2436 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4766
timestamp 1680363874
transform 1 0 2460 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5270
timestamp 1680363874
transform 1 0 2500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1680363874
transform 1 0 2444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1680363874
transform 1 0 2460 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4814
timestamp 1680363874
transform 1 0 2556 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5271
timestamp 1680363874
transform 1 0 2556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1680363874
transform 1 0 2564 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4767
timestamp 1680363874
transform 1 0 2596 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5273
timestamp 1680363874
transform 1 0 2628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1680363874
transform 1 0 2676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1680363874
transform 1 0 2580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1680363874
transform 1 0 2596 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4758
timestamp 1680363874
transform 1 0 2708 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5275
timestamp 1680363874
transform 1 0 2708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1680363874
transform 1 0 2740 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4874
timestamp 1680363874
transform 1 0 2740 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5276
timestamp 1680363874
transform 1 0 2756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1680363874
transform 1 0 2764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1680363874
transform 1 0 2756 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4768
timestamp 1680363874
transform 1 0 2772 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5278
timestamp 1680363874
transform 1 0 2804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1680363874
transform 1 0 2780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1680363874
transform 1 0 2796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1680363874
transform 1 0 2812 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4889
timestamp 1680363874
transform 1 0 2820 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1680363874
transform 1 0 2868 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5369
timestamp 1680363874
transform 1 0 2868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1680363874
transform 1 0 2900 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1680363874
transform 1 0 2884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1680363874
transform 1 0 2908 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4752
timestamp 1680363874
transform 1 0 2948 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1680363874
transform 1 0 2956 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5221
timestamp 1680363874
transform 1 0 2948 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1680363874
transform 1 0 2956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1680363874
transform 1 0 2972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1680363874
transform 1 0 2988 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4753
timestamp 1680363874
transform 1 0 3004 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_5222
timestamp 1680363874
transform 1 0 3004 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4816
timestamp 1680363874
transform 1 0 3036 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1680363874
transform 1 0 3052 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1680363874
transform 1 0 3060 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1680363874
transform 1 0 3076 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5223
timestamp 1680363874
transform 1 0 3068 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1680363874
transform 1 0 3052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1680363874
transform 1 0 3036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1680363874
transform 1 0 3044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1680363874
transform 1 0 3076 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4818
timestamp 1680363874
transform 1 0 3108 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1680363874
transform 1 0 3124 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5373
timestamp 1680363874
transform 1 0 3116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1680363874
transform 1 0 3132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1680363874
transform 1 0 3156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1680363874
transform 1 0 3172 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4819
timestamp 1680363874
transform 1 0 3212 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5285
timestamp 1680363874
transform 1 0 3204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1680363874
transform 1 0 3212 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4820
timestamp 1680363874
transform 1 0 3244 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1680363874
transform 1 0 3284 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1680363874
transform 1 0 3276 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5287
timestamp 1680363874
transform 1 0 3268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1680363874
transform 1 0 3284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1680363874
transform 1 0 3276 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4875
timestamp 1680363874
transform 1 0 3284 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5377
timestamp 1680363874
transform 1 0 3324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1680363874
transform 1 0 3340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1680363874
transform 1 0 3364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1680363874
transform 1 0 3380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1680363874
transform 1 0 3356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1680363874
transform 1 0 3372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1680363874
transform 1 0 3380 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4890
timestamp 1680363874
transform 1 0 3380 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5292
timestamp 1680363874
transform 1 0 3420 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4876
timestamp 1680363874
transform 1 0 3460 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1680363874
transform 1 0 3476 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5293
timestamp 1680363874
transform 1 0 3476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1680363874
transform 1 0 3492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1680363874
transform 1 0 3508 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1680363874
transform 1 0 3484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1680363874
transform 1 0 3500 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4853
timestamp 1680363874
transform 1 0 3508 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1680363874
transform 1 0 3524 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5296
timestamp 1680363874
transform 1 0 3524 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1680363874
transform 1 0 3516 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4877
timestamp 1680363874
transform 1 0 3500 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1680363874
transform 1 0 3532 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1680363874
transform 1 0 3532 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1680363874
transform 1 0 3596 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1680363874
transform 1 0 3588 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5297
timestamp 1680363874
transform 1 0 3580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1680363874
transform 1 0 3596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1680363874
transform 1 0 3612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1680363874
transform 1 0 3588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1680363874
transform 1 0 3604 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4855
timestamp 1680363874
transform 1 0 3612 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1680363874
transform 1 0 3660 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1680363874
transform 1 0 3716 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1680363874
transform 1 0 3740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1680363874
transform 1 0 3652 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5300
timestamp 1680363874
transform 1 0 3692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1680363874
transform 1 0 3740 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4878
timestamp 1680363874
transform 1 0 3740 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1680363874
transform 1 0 3764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1680363874
transform 1 0 3756 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5387
timestamp 1680363874
transform 1 0 3764 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4826
timestamp 1680363874
transform 1 0 3788 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5301
timestamp 1680363874
transform 1 0 3788 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4792
timestamp 1680363874
transform 1 0 3804 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1680363874
transform 1 0 3828 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5302
timestamp 1680363874
transform 1 0 3828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1680363874
transform 1 0 3804 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4879
timestamp 1680363874
transform 1 0 3804 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5303
timestamp 1680363874
transform 1 0 3892 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1680363874
transform 1 0 3908 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4793
timestamp 1680363874
transform 1 0 3948 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5304
timestamp 1680363874
transform 1 0 3924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1680363874
transform 1 0 3940 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1680363874
transform 1 0 3956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1680363874
transform 1 0 3948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1680363874
transform 1 0 3956 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4794
timestamp 1680363874
transform 1 0 4028 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1680363874
transform 1 0 4020 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1680363874
transform 1 0 4060 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5307
timestamp 1680363874
transform 1 0 4020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1680363874
transform 1 0 4028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1680363874
transform 1 0 4060 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4857
timestamp 1680363874
transform 1 0 4036 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5392
timestamp 1680363874
transform 1 0 4108 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4880
timestamp 1680363874
transform 1 0 4108 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5310
timestamp 1680363874
transform 1 0 4124 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4858
timestamp 1680363874
transform 1 0 4124 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5411
timestamp 1680363874
transform 1 0 4124 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1680363874
transform 1 0 4140 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4795
timestamp 1680363874
transform 1 0 4300 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1680363874
transform 1 0 4292 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5311
timestamp 1680363874
transform 1 0 4252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1680363874
transform 1 0 4292 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4881
timestamp 1680363874
transform 1 0 4292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1680363874
transform 1 0 4316 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5312
timestamp 1680363874
transform 1 0 4316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1680363874
transform 1 0 4348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1680363874
transform 1 0 4340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1680363874
transform 1 0 4356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1680363874
transform 1 0 4364 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4882
timestamp 1680363874
transform 1 0 4340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1680363874
transform 1 0 4364 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1680363874
transform 1 0 4332 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1680363874
transform 1 0 4356 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5314
timestamp 1680363874
transform 1 0 4388 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4859
timestamp 1680363874
transform 1 0 4412 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5413
timestamp 1680363874
transform 1 0 4412 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4893
timestamp 1680363874
transform 1 0 4412 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5315
timestamp 1680363874
transform 1 0 4444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1680363874
transform 1 0 4460 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4839
timestamp 1680363874
transform 1 0 4468 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5317
timestamp 1680363874
transform 1 0 4476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1680363874
transform 1 0 4492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1680363874
transform 1 0 4468 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4860
timestamp 1680363874
transform 1 0 4484 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1680363874
transform 1 0 4508 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1680363874
transform 1 0 4508 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1680363874
transform 1 0 4532 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5414
timestamp 1680363874
transform 1 0 4532 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4771
timestamp 1680363874
transform 1 0 4556 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5398
timestamp 1680363874
transform 1 0 4548 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4840
timestamp 1680363874
transform 1 0 4572 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1680363874
transform 1 0 4604 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5319
timestamp 1680363874
transform 1 0 4580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1680363874
transform 1 0 4604 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4862
timestamp 1680363874
transform 1 0 4564 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5399
timestamp 1680363874
transform 1 0 4572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1680363874
transform 1 0 4588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4884
timestamp 1680363874
transform 1 0 4588 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5401
timestamp 1680363874
transform 1 0 4612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1680363874
transform 1 0 4628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1680363874
transform 1 0 4644 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4841
timestamp 1680363874
transform 1 0 4652 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5323
timestamp 1680363874
transform 1 0 4660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1680363874
transform 1 0 4636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1680363874
transform 1 0 4652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1680363874
transform 1 0 4660 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4842
timestamp 1680363874
transform 1 0 4708 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5405
timestamp 1680363874
transform 1 0 4756 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4760
timestamp 1680363874
transform 1 0 4788 0 1 2255
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_50
timestamp 1680363874
transform 1 0 48 0 1 2170
box -10 -3 10 3
use FILL  FILL_5866
timestamp 1680363874
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_5868
timestamp 1680363874
transform 1 0 80 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4894
timestamp 1680363874
transform 1 0 100 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_376
timestamp 1680363874
transform 1 0 88 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_377
timestamp 1680363874
transform 1 0 104 0 1 2170
box -9 -3 26 105
use FILL  FILL_5870
timestamp 1680363874
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_5876
timestamp 1680363874
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_5877
timestamp 1680363874
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_5878
timestamp 1680363874
transform 1 0 144 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_27
timestamp 1680363874
transform 1 0 152 0 1 2170
box -8 -3 40 105
use FILL  FILL_5879
timestamp 1680363874
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_5880
timestamp 1680363874
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_5881
timestamp 1680363874
transform 1 0 200 0 1 2170
box -8 -3 16 105
use FILL  FILL_5886
timestamp 1680363874
transform 1 0 208 0 1 2170
box -8 -3 16 105
use FILL  FILL_5888
timestamp 1680363874
transform 1 0 216 0 1 2170
box -8 -3 16 105
use FILL  FILL_5890
timestamp 1680363874
transform 1 0 224 0 1 2170
box -8 -3 16 105
use FILL  FILL_5891
timestamp 1680363874
transform 1 0 232 0 1 2170
box -8 -3 16 105
use FILL  FILL_5892
timestamp 1680363874
transform 1 0 240 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_29
timestamp 1680363874
transform 1 0 248 0 1 2170
box -8 -3 40 105
use FILL  FILL_5893
timestamp 1680363874
transform 1 0 280 0 1 2170
box -8 -3 16 105
use FILL  FILL_5894
timestamp 1680363874
transform 1 0 288 0 1 2170
box -8 -3 16 105
use FILL  FILL_5897
timestamp 1680363874
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_5899
timestamp 1680363874
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_5901
timestamp 1680363874
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_5902
timestamp 1680363874
transform 1 0 320 0 1 2170
box -8 -3 16 105
use AOI21X1  AOI21X1_12
timestamp 1680363874
transform -1 0 360 0 1 2170
box -7 -3 39 105
use FILL  FILL_5903
timestamp 1680363874
transform 1 0 360 0 1 2170
box -8 -3 16 105
use FILL  FILL_5907
timestamp 1680363874
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_5908
timestamp 1680363874
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_5909
timestamp 1680363874
transform 1 0 384 0 1 2170
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1680363874
transform -1 0 424 0 1 2170
box -8 -3 40 105
use FILL  FILL_5910
timestamp 1680363874
transform 1 0 424 0 1 2170
box -8 -3 16 105
use FILL  FILL_5911
timestamp 1680363874
transform 1 0 432 0 1 2170
box -8 -3 16 105
use FILL  FILL_5912
timestamp 1680363874
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_5913
timestamp 1680363874
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_5914
timestamp 1680363874
transform 1 0 456 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_136
timestamp 1680363874
transform -1 0 496 0 1 2170
box -8 -3 34 105
use FILL  FILL_5915
timestamp 1680363874
transform 1 0 496 0 1 2170
box -8 -3 16 105
use FILL  FILL_5916
timestamp 1680363874
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_5917
timestamp 1680363874
transform 1 0 512 0 1 2170
box -8 -3 16 105
use FILL  FILL_5918
timestamp 1680363874
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_5919
timestamp 1680363874
transform 1 0 528 0 1 2170
box -8 -3 16 105
use FILL  FILL_5920
timestamp 1680363874
transform 1 0 536 0 1 2170
box -8 -3 16 105
use FILL  FILL_5921
timestamp 1680363874
transform 1 0 544 0 1 2170
box -8 -3 16 105
use FILL  FILL_5922
timestamp 1680363874
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_5923
timestamp 1680363874
transform 1 0 560 0 1 2170
box -8 -3 16 105
use FILL  FILL_5924
timestamp 1680363874
transform 1 0 568 0 1 2170
box -8 -3 16 105
use FILL  FILL_5930
timestamp 1680363874
transform 1 0 576 0 1 2170
box -8 -3 16 105
use FILL  FILL_5932
timestamp 1680363874
transform 1 0 584 0 1 2170
box -8 -3 16 105
use FILL  FILL_5934
timestamp 1680363874
transform 1 0 592 0 1 2170
box -8 -3 16 105
use FILL  FILL_5936
timestamp 1680363874
transform 1 0 600 0 1 2170
box -8 -3 16 105
use FILL  FILL_5938
timestamp 1680363874
transform 1 0 608 0 1 2170
box -8 -3 16 105
use FILL  FILL_5939
timestamp 1680363874
transform 1 0 616 0 1 2170
box -8 -3 16 105
use FILL  FILL_5940
timestamp 1680363874
transform 1 0 624 0 1 2170
box -8 -3 16 105
use FILL  FILL_5941
timestamp 1680363874
transform 1 0 632 0 1 2170
box -8 -3 16 105
use FILL  FILL_5943
timestamp 1680363874
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_5945
timestamp 1680363874
transform 1 0 648 0 1 2170
box -8 -3 16 105
use FILL  FILL_5947
timestamp 1680363874
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_5949
timestamp 1680363874
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_5951
timestamp 1680363874
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_5953
timestamp 1680363874
transform 1 0 680 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4895
timestamp 1680363874
transform 1 0 700 0 1 2175
box -3 -3 3 3
use FILL  FILL_5954
timestamp 1680363874
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_5955
timestamp 1680363874
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_5956
timestamp 1680363874
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_5958
timestamp 1680363874
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_5960
timestamp 1680363874
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_5962
timestamp 1680363874
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_5964
timestamp 1680363874
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FAX1  FAX1_14
timestamp 1680363874
transform -1 0 864 0 1 2170
box -5 -3 126 105
use FILL  FILL_5965
timestamp 1680363874
transform 1 0 864 0 1 2170
box -8 -3 16 105
use FILL  FILL_5966
timestamp 1680363874
transform 1 0 872 0 1 2170
box -8 -3 16 105
use XOR2X1  XOR2X1_2
timestamp 1680363874
transform -1 0 936 0 1 2170
box -8 -3 64 105
use FILL  FILL_5967
timestamp 1680363874
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_5968
timestamp 1680363874
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_5978
timestamp 1680363874
transform 1 0 952 0 1 2170
box -8 -3 16 105
use FILL  FILL_5980
timestamp 1680363874
transform 1 0 960 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_45
timestamp 1680363874
transform 1 0 968 0 1 2170
box -8 -3 32 105
use FILL  FILL_5982
timestamp 1680363874
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_5984
timestamp 1680363874
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_5986
timestamp 1680363874
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use FILL  FILL_5988
timestamp 1680363874
transform 1 0 1016 0 1 2170
box -8 -3 16 105
use FILL  FILL_5989
timestamp 1680363874
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_5990
timestamp 1680363874
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_5991
timestamp 1680363874
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_31
timestamp 1680363874
transform -1 0 1080 0 1 2170
box -8 -3 40 105
use FILL  FILL_5992
timestamp 1680363874
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_5998
timestamp 1680363874
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6000
timestamp 1680363874
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6002
timestamp 1680363874
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6004
timestamp 1680363874
transform 1 0 1112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6006
timestamp 1680363874
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_33
timestamp 1680363874
transform -1 0 1160 0 1 2170
box -8 -3 40 105
use FILL  FILL_6007
timestamp 1680363874
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_6012
timestamp 1680363874
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_6014
timestamp 1680363874
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6016
timestamp 1680363874
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_6018
timestamp 1680363874
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6020
timestamp 1680363874
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6022
timestamp 1680363874
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6023
timestamp 1680363874
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6024
timestamp 1680363874
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6025
timestamp 1680363874
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6026
timestamp 1680363874
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_6028
timestamp 1680363874
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_6030
timestamp 1680363874
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_6032
timestamp 1680363874
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_6034
timestamp 1680363874
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_6036
timestamp 1680363874
transform 1 0 1280 0 1 2170
box -8 -3 16 105
use FILL  FILL_6037
timestamp 1680363874
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6038
timestamp 1680363874
transform 1 0 1296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6040
timestamp 1680363874
transform 1 0 1304 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4896
timestamp 1680363874
transform 1 0 1348 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_196
timestamp 1680363874
transform 1 0 1312 0 1 2170
box -8 -3 46 105
use FILL  FILL_6042
timestamp 1680363874
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6043
timestamp 1680363874
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_6044
timestamp 1680363874
transform 1 0 1368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6045
timestamp 1680363874
transform 1 0 1376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6046
timestamp 1680363874
transform 1 0 1384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6052
timestamp 1680363874
transform 1 0 1392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6054
timestamp 1680363874
transform 1 0 1400 0 1 2170
box -8 -3 16 105
use FILL  FILL_6056
timestamp 1680363874
transform 1 0 1408 0 1 2170
box -8 -3 16 105
use FILL  FILL_6058
timestamp 1680363874
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_6060
timestamp 1680363874
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4897
timestamp 1680363874
transform 1 0 1468 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_256
timestamp 1680363874
transform 1 0 1432 0 1 2170
box -8 -3 46 105
use FILL  FILL_6062
timestamp 1680363874
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_6063
timestamp 1680363874
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_6064
timestamp 1680363874
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_6065
timestamp 1680363874
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_6066
timestamp 1680363874
transform 1 0 1504 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_382
timestamp 1680363874
transform -1 0 1528 0 1 2170
box -9 -3 26 105
use FILL  FILL_6067
timestamp 1680363874
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6069
timestamp 1680363874
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6070
timestamp 1680363874
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_6071
timestamp 1680363874
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6072
timestamp 1680363874
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_257
timestamp 1680363874
transform 1 0 1568 0 1 2170
box -8 -3 46 105
use FILL  FILL_6073
timestamp 1680363874
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6074
timestamp 1680363874
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_6075
timestamp 1680363874
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_383
timestamp 1680363874
transform -1 0 1648 0 1 2170
box -9 -3 26 105
use FILL  FILL_6076
timestamp 1680363874
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_6080
timestamp 1680363874
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_6082
timestamp 1680363874
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_6084
timestamp 1680363874
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4898
timestamp 1680363874
transform 1 0 1716 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_258
timestamp 1680363874
transform 1 0 1680 0 1 2170
box -8 -3 46 105
use FILL  FILL_6085
timestamp 1680363874
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6088
timestamp 1680363874
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_384
timestamp 1680363874
transform -1 0 1752 0 1 2170
box -9 -3 26 105
use FILL  FILL_6089
timestamp 1680363874
transform 1 0 1752 0 1 2170
box -8 -3 16 105
use FILL  FILL_6094
timestamp 1680363874
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_6096
timestamp 1680363874
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_6098
timestamp 1680363874
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6099
timestamp 1680363874
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4899
timestamp 1680363874
transform 1 0 1812 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_260
timestamp 1680363874
transform 1 0 1792 0 1 2170
box -8 -3 46 105
use FILL  FILL_6100
timestamp 1680363874
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_6104
timestamp 1680363874
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_6105
timestamp 1680363874
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6106
timestamp 1680363874
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6107
timestamp 1680363874
transform 1 0 1864 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_385
timestamp 1680363874
transform -1 0 1888 0 1 2170
box -9 -3 26 105
use FILL  FILL_6108
timestamp 1680363874
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6109
timestamp 1680363874
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_327
timestamp 1680363874
transform -1 0 2000 0 1 2170
box -8 -3 104 105
use FILL  FILL_6110
timestamp 1680363874
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6111
timestamp 1680363874
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6112
timestamp 1680363874
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_6113
timestamp 1680363874
transform 1 0 2024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6114
timestamp 1680363874
transform 1 0 2032 0 1 2170
box -8 -3 16 105
use FILL  FILL_6115
timestamp 1680363874
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_386
timestamp 1680363874
transform 1 0 2048 0 1 2170
box -9 -3 26 105
use FILL  FILL_6116
timestamp 1680363874
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_6120
timestamp 1680363874
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4900
timestamp 1680363874
transform 1 0 2092 0 1 2175
box -3 -3 3 3
use FILL  FILL_6122
timestamp 1680363874
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_262
timestamp 1680363874
transform -1 0 2128 0 1 2170
box -8 -3 46 105
use FILL  FILL_6124
timestamp 1680363874
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6126
timestamp 1680363874
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4901
timestamp 1680363874
transform 1 0 2156 0 1 2175
box -3 -3 3 3
use FILL  FILL_6128
timestamp 1680363874
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_6130
timestamp 1680363874
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_6132
timestamp 1680363874
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_35
timestamp 1680363874
transform -1 0 2200 0 1 2170
box -8 -3 40 105
use FILL  FILL_6133
timestamp 1680363874
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6134
timestamp 1680363874
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6135
timestamp 1680363874
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6139
timestamp 1680363874
transform 1 0 2224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6141
timestamp 1680363874
transform 1 0 2232 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_197
timestamp 1680363874
transform -1 0 2280 0 1 2170
box -8 -3 46 105
use FILL  FILL_6142
timestamp 1680363874
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_6143
timestamp 1680363874
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6144
timestamp 1680363874
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4902
timestamp 1680363874
transform 1 0 2316 0 1 2175
box -3 -3 3 3
use FILL  FILL_6145
timestamp 1680363874
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_265
timestamp 1680363874
transform 1 0 2312 0 1 2170
box -8 -3 46 105
use FILL  FILL_6151
timestamp 1680363874
transform 1 0 2352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6152
timestamp 1680363874
transform 1 0 2360 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_388
timestamp 1680363874
transform -1 0 2384 0 1 2170
box -9 -3 26 105
use FILL  FILL_6153
timestamp 1680363874
transform 1 0 2384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6159
timestamp 1680363874
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6161
timestamp 1680363874
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_6163
timestamp 1680363874
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use AND2X2  AND2X2_19
timestamp 1680363874
transform -1 0 2448 0 1 2170
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_330
timestamp 1680363874
transform 1 0 2448 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_389
timestamp 1680363874
transform 1 0 2544 0 1 2170
box -9 -3 26 105
use FILL  FILL_6165
timestamp 1680363874
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_390
timestamp 1680363874
transform -1 0 2584 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_331
timestamp 1680363874
transform 1 0 2584 0 1 2170
box -8 -3 104 105
use FILL  FILL_6166
timestamp 1680363874
transform 1 0 2680 0 1 2170
box -8 -3 16 105
use FILL  FILL_6167
timestamp 1680363874
transform 1 0 2688 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_391
timestamp 1680363874
transform -1 0 2712 0 1 2170
box -9 -3 26 105
use FILL  FILL_6168
timestamp 1680363874
transform 1 0 2712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6187
timestamp 1680363874
transform 1 0 2720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6189
timestamp 1680363874
transform 1 0 2728 0 1 2170
box -8 -3 16 105
use FILL  FILL_6191
timestamp 1680363874
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_394
timestamp 1680363874
transform -1 0 2760 0 1 2170
box -9 -3 26 105
use FILL  FILL_6192
timestamp 1680363874
transform 1 0 2760 0 1 2170
box -8 -3 16 105
use FILL  FILL_6193
timestamp 1680363874
transform 1 0 2768 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_266
timestamp 1680363874
transform 1 0 2776 0 1 2170
box -8 -3 46 105
use FILL  FILL_6194
timestamp 1680363874
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use FILL  FILL_6195
timestamp 1680363874
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_6196
timestamp 1680363874
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_6197
timestamp 1680363874
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_6200
timestamp 1680363874
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6202
timestamp 1680363874
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6204
timestamp 1680363874
transform 1 0 2864 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_137
timestamp 1680363874
transform 1 0 2872 0 1 2170
box -8 -3 34 105
use FILL  FILL_6206
timestamp 1680363874
transform 1 0 2904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6207
timestamp 1680363874
transform 1 0 2912 0 1 2170
box -8 -3 16 105
use FILL  FILL_6208
timestamp 1680363874
transform 1 0 2920 0 1 2170
box -8 -3 16 105
use FILL  FILL_6209
timestamp 1680363874
transform 1 0 2928 0 1 2170
box -8 -3 16 105
use FILL  FILL_6214
timestamp 1680363874
transform 1 0 2936 0 1 2170
box -8 -3 16 105
use FILL  FILL_6216
timestamp 1680363874
transform 1 0 2944 0 1 2170
box -8 -3 16 105
use FILL  FILL_6218
timestamp 1680363874
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_139
timestamp 1680363874
transform 1 0 2960 0 1 2170
box -8 -3 34 105
use FILL  FILL_6220
timestamp 1680363874
transform 1 0 2992 0 1 2170
box -8 -3 16 105
use FILL  FILL_6221
timestamp 1680363874
transform 1 0 3000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6222
timestamp 1680363874
transform 1 0 3008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6223
timestamp 1680363874
transform 1 0 3016 0 1 2170
box -8 -3 16 105
use FILL  FILL_6224
timestamp 1680363874
transform 1 0 3024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6225
timestamp 1680363874
transform 1 0 3032 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_140
timestamp 1680363874
transform 1 0 3040 0 1 2170
box -8 -3 34 105
use FILL  FILL_6226
timestamp 1680363874
transform 1 0 3072 0 1 2170
box -8 -3 16 105
use FILL  FILL_6230
timestamp 1680363874
transform 1 0 3080 0 1 2170
box -8 -3 16 105
use FILL  FILL_6232
timestamp 1680363874
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6234
timestamp 1680363874
transform 1 0 3096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6236
timestamp 1680363874
transform 1 0 3104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6237
timestamp 1680363874
transform 1 0 3112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6238
timestamp 1680363874
transform 1 0 3120 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_141
timestamp 1680363874
transform -1 0 3160 0 1 2170
box -8 -3 34 105
use FILL  FILL_6239
timestamp 1680363874
transform 1 0 3160 0 1 2170
box -8 -3 16 105
use FILL  FILL_6243
timestamp 1680363874
transform 1 0 3168 0 1 2170
box -8 -3 16 105
use FILL  FILL_6245
timestamp 1680363874
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6247
timestamp 1680363874
transform 1 0 3184 0 1 2170
box -8 -3 16 105
use FILL  FILL_6249
timestamp 1680363874
transform 1 0 3192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6250
timestamp 1680363874
transform 1 0 3200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6251
timestamp 1680363874
transform 1 0 3208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6252
timestamp 1680363874
transform 1 0 3216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6253
timestamp 1680363874
transform 1 0 3224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6256
timestamp 1680363874
transform 1 0 3232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6258
timestamp 1680363874
transform 1 0 3240 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_201
timestamp 1680363874
transform -1 0 3288 0 1 2170
box -8 -3 46 105
use FILL  FILL_6259
timestamp 1680363874
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6260
timestamp 1680363874
transform 1 0 3296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6265
timestamp 1680363874
transform 1 0 3304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6267
timestamp 1680363874
transform 1 0 3312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6269
timestamp 1680363874
transform 1 0 3320 0 1 2170
box -8 -3 16 105
use FILL  FILL_6271
timestamp 1680363874
transform 1 0 3328 0 1 2170
box -8 -3 16 105
use FILL  FILL_6273
timestamp 1680363874
transform 1 0 3336 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_202
timestamp 1680363874
transform 1 0 3344 0 1 2170
box -8 -3 46 105
use FILL  FILL_6275
timestamp 1680363874
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6276
timestamp 1680363874
transform 1 0 3392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6277
timestamp 1680363874
transform 1 0 3400 0 1 2170
box -8 -3 16 105
use AND2X2  AND2X2_22
timestamp 1680363874
transform 1 0 3408 0 1 2170
box -8 -3 40 105
use FILL  FILL_6278
timestamp 1680363874
transform 1 0 3440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6288
timestamp 1680363874
transform 1 0 3448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6290
timestamp 1680363874
transform 1 0 3456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6291
timestamp 1680363874
transform 1 0 3464 0 1 2170
box -8 -3 16 105
use FILL  FILL_6292
timestamp 1680363874
transform 1 0 3472 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_267
timestamp 1680363874
transform 1 0 3480 0 1 2170
box -8 -3 46 105
use FILL  FILL_6293
timestamp 1680363874
transform 1 0 3520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6294
timestamp 1680363874
transform 1 0 3528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6295
timestamp 1680363874
transform 1 0 3536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6296
timestamp 1680363874
transform 1 0 3544 0 1 2170
box -8 -3 16 105
use FILL  FILL_6301
timestamp 1680363874
transform 1 0 3552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6303
timestamp 1680363874
transform 1 0 3560 0 1 2170
box -8 -3 16 105
use FILL  FILL_6305
timestamp 1680363874
transform 1 0 3568 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_203
timestamp 1680363874
transform 1 0 3576 0 1 2170
box -8 -3 46 105
use FILL  FILL_6307
timestamp 1680363874
transform 1 0 3616 0 1 2170
box -8 -3 16 105
use FILL  FILL_6308
timestamp 1680363874
transform 1 0 3624 0 1 2170
box -8 -3 16 105
use FILL  FILL_6309
timestamp 1680363874
transform 1 0 3632 0 1 2170
box -8 -3 16 105
use FILL  FILL_6310
timestamp 1680363874
transform 1 0 3640 0 1 2170
box -8 -3 16 105
use FILL  FILL_6315
timestamp 1680363874
transform 1 0 3648 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_334
timestamp 1680363874
transform -1 0 3752 0 1 2170
box -8 -3 104 105
use FILL  FILL_6316
timestamp 1680363874
transform 1 0 3752 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_395
timestamp 1680363874
transform 1 0 3760 0 1 2170
box -9 -3 26 105
use FILL  FILL_6317
timestamp 1680363874
transform 1 0 3776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6318
timestamp 1680363874
transform 1 0 3784 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_335
timestamp 1680363874
transform 1 0 3792 0 1 2170
box -8 -3 104 105
use FILL  FILL_6319
timestamp 1680363874
transform 1 0 3888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6337
timestamp 1680363874
transform 1 0 3896 0 1 2170
box -8 -3 16 105
use FILL  FILL_6339
timestamp 1680363874
transform 1 0 3904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6341
timestamp 1680363874
transform 1 0 3912 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_205
timestamp 1680363874
transform 1 0 3920 0 1 2170
box -8 -3 46 105
use FILL  FILL_6343
timestamp 1680363874
transform 1 0 3960 0 1 2170
box -8 -3 16 105
use FILL  FILL_6344
timestamp 1680363874
transform 1 0 3968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6345
timestamp 1680363874
transform 1 0 3976 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_397
timestamp 1680363874
transform 1 0 3984 0 1 2170
box -9 -3 26 105
use FILL  FILL_6346
timestamp 1680363874
transform 1 0 4000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6353
timestamp 1680363874
transform 1 0 4008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6355
timestamp 1680363874
transform 1 0 4016 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_337
timestamp 1680363874
transform -1 0 4120 0 1 2170
box -8 -3 104 105
use FILL  FILL_6356
timestamp 1680363874
transform 1 0 4120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6357
timestamp 1680363874
transform 1 0 4128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6358
timestamp 1680363874
transform 1 0 4136 0 1 2170
box -8 -3 16 105
use FILL  FILL_6359
timestamp 1680363874
transform 1 0 4144 0 1 2170
box -8 -3 16 105
use FILL  FILL_6360
timestamp 1680363874
transform 1 0 4152 0 1 2170
box -8 -3 16 105
use FILL  FILL_6361
timestamp 1680363874
transform 1 0 4160 0 1 2170
box -8 -3 16 105
use FILL  FILL_6362
timestamp 1680363874
transform 1 0 4168 0 1 2170
box -8 -3 16 105
use FILL  FILL_6363
timestamp 1680363874
transform 1 0 4176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6368
timestamp 1680363874
transform 1 0 4184 0 1 2170
box -8 -3 16 105
use FILL  FILL_6370
timestamp 1680363874
transform 1 0 4192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6372
timestamp 1680363874
transform 1 0 4200 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_339
timestamp 1680363874
transform -1 0 4304 0 1 2170
box -8 -3 104 105
use FILL  FILL_6373
timestamp 1680363874
transform 1 0 4304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6376
timestamp 1680363874
transform 1 0 4312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6378
timestamp 1680363874
transform 1 0 4320 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4903
timestamp 1680363874
transform 1 0 4348 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_206
timestamp 1680363874
transform 1 0 4328 0 1 2170
box -8 -3 46 105
use FILL  FILL_6380
timestamp 1680363874
transform 1 0 4368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6381
timestamp 1680363874
transform 1 0 4376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6382
timestamp 1680363874
transform 1 0 4384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6383
timestamp 1680363874
transform 1 0 4392 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4904
timestamp 1680363874
transform 1 0 4412 0 1 2175
box -3 -3 3 3
use FILL  FILL_6384
timestamp 1680363874
transform 1 0 4400 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_61
timestamp 1680363874
transform 1 0 4408 0 1 2170
box -8 -3 32 105
use FILL  FILL_6385
timestamp 1680363874
transform 1 0 4432 0 1 2170
box -8 -3 16 105
use FILL  FILL_6386
timestamp 1680363874
transform 1 0 4440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6387
timestamp 1680363874
transform 1 0 4448 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_207
timestamp 1680363874
transform -1 0 4496 0 1 2170
box -8 -3 46 105
use FILL  FILL_6388
timestamp 1680363874
transform 1 0 4496 0 1 2170
box -8 -3 16 105
use FILL  FILL_6397
timestamp 1680363874
transform 1 0 4504 0 1 2170
box -8 -3 16 105
use FILL  FILL_6399
timestamp 1680363874
transform 1 0 4512 0 1 2170
box -8 -3 16 105
use FILL  FILL_6401
timestamp 1680363874
transform 1 0 4520 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_62
timestamp 1680363874
transform 1 0 4528 0 1 2170
box -8 -3 32 105
use FILL  FILL_6402
timestamp 1680363874
transform 1 0 4552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6403
timestamp 1680363874
transform 1 0 4560 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_271
timestamp 1680363874
transform -1 0 4608 0 1 2170
box -8 -3 46 105
use FILL  FILL_6404
timestamp 1680363874
transform 1 0 4608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6409
timestamp 1680363874
transform 1 0 4616 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_208
timestamp 1680363874
transform 1 0 4624 0 1 2170
box -8 -3 46 105
use FILL  FILL_6411
timestamp 1680363874
transform 1 0 4664 0 1 2170
box -8 -3 16 105
use FILL  FILL_6413
timestamp 1680363874
transform 1 0 4672 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_399
timestamp 1680363874
transform 1 0 4680 0 1 2170
box -9 -3 26 105
use FILL  FILL_6415
timestamp 1680363874
transform 1 0 4696 0 1 2170
box -8 -3 16 105
use FILL  FILL_6416
timestamp 1680363874
transform 1 0 4704 0 1 2170
box -8 -3 16 105
use FILL  FILL_6417
timestamp 1680363874
transform 1 0 4712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6418
timestamp 1680363874
transform 1 0 4720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6419
timestamp 1680363874
transform 1 0 4728 0 1 2170
box -8 -3 16 105
use FILL  FILL_6420
timestamp 1680363874
transform 1 0 4736 0 1 2170
box -8 -3 16 105
use FILL  FILL_6421
timestamp 1680363874
transform 1 0 4744 0 1 2170
box -8 -3 16 105
use FILL  FILL_6422
timestamp 1680363874
transform 1 0 4752 0 1 2170
box -8 -3 16 105
use FILL  FILL_6423
timestamp 1680363874
transform 1 0 4760 0 1 2170
box -8 -3 16 105
use FILL  FILL_6424
timestamp 1680363874
transform 1 0 4768 0 1 2170
box -8 -3 16 105
use FILL  FILL_6425
timestamp 1680363874
transform 1 0 4776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6426
timestamp 1680363874
transform 1 0 4784 0 1 2170
box -8 -3 16 105
use FILL  FILL_6427
timestamp 1680363874
transform 1 0 4792 0 1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_51
timestamp 1680363874
transform 1 0 4827 0 1 2170
box -10 -3 10 3
use M2_M1  M2_M1_5591
timestamp 1680363874
transform 1 0 92 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4932
timestamp 1680363874
transform 1 0 116 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5497
timestamp 1680363874
transform 1 0 156 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1680363874
transform 1 0 164 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1680363874
transform 1 0 156 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4933
timestamp 1680363874
transform 1 0 188 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5423
timestamp 1680363874
transform 1 0 188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1680363874
transform 1 0 180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5010
timestamp 1680363874
transform 1 0 180 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1680363874
transform 1 0 204 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5499
timestamp 1680363874
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4914
timestamp 1680363874
transform 1 0 236 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1680363874
transform 1 0 252 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5416
timestamp 1680363874
transform 1 0 252 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1680363874
transform 1 0 252 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4993
timestamp 1680363874
transform 1 0 244 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5500
timestamp 1680363874
transform 1 0 268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1680363874
transform 1 0 260 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5011
timestamp 1680363874
transform 1 0 268 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5612
timestamp 1680363874
transform 1 0 260 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_5042
timestamp 1680363874
transform 1 0 284 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1680363874
transform 1 0 300 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5594
timestamp 1680363874
transform 1 0 300 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5056
timestamp 1680363874
transform 1 0 292 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1680363874
transform 1 0 316 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5425
timestamp 1680363874
transform 1 0 324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1680363874
transform 1 0 316 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1680363874
transform 1 0 348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1680363874
transform 1 0 340 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5043
timestamp 1680363874
transform 1 0 348 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1680363874
transform 1 0 348 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1680363874
transform 1 0 364 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1680363874
transform 1 0 380 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5502
timestamp 1680363874
transform 1 0 372 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4936
timestamp 1680363874
transform 1 0 420 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1680363874
transform 1 0 412 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5427
timestamp 1680363874
transform 1 0 420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1680363874
transform 1 0 412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1680363874
transform 1 0 444 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1680363874
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5012
timestamp 1680363874
transform 1 0 420 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1680363874
transform 1 0 516 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1680363874
transform 1 0 564 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5418
timestamp 1680363874
transform 1 0 460 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1680363874
transform 1 0 452 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4969
timestamp 1680363874
transform 1 0 460 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1680363874
transform 1 0 572 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5429
timestamp 1680363874
transform 1 0 564 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4994
timestamp 1680363874
transform 1 0 524 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5505
timestamp 1680363874
transform 1 0 548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1680363874
transform 1 0 556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5044
timestamp 1680363874
transform 1 0 564 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1680363874
transform 1 0 532 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1680363874
transform 1 0 564 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1680363874
transform 1 0 588 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5430
timestamp 1680363874
transform 1 0 596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1680363874
transform 1 0 588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4920
timestamp 1680363874
transform 1 0 628 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1680363874
transform 1 0 628 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5431
timestamp 1680363874
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_5013
timestamp 1680363874
transform 1 0 620 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5596
timestamp 1680363874
transform 1 0 628 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4921
timestamp 1680363874
transform 1 0 676 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5597
timestamp 1680363874
transform 1 0 700 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1680363874
transform 1 0 724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1680363874
transform 1 0 716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1680363874
transform 1 0 740 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5014
timestamp 1680363874
transform 1 0 764 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5433
timestamp 1680363874
transform 1 0 780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1680363874
transform 1 0 772 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5074
timestamp 1680363874
transform 1 0 772 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1680363874
transform 1 0 804 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1680363874
transform 1 0 796 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1680363874
transform 1 0 812 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5419
timestamp 1680363874
transform 1 0 932 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_4971
timestamp 1680363874
transform 1 0 860 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1680363874
transform 1 0 948 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5434
timestamp 1680363874
transform 1 0 940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1680363874
transform 1 0 948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1680363874
transform 1 0 828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1680363874
transform 1 0 836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1680363874
transform 1 0 844 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4996
timestamp 1680363874
transform 1 0 868 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1680363874
transform 1 0 940 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5513
timestamp 1680363874
transform 1 0 956 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5058
timestamp 1680363874
transform 1 0 948 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1680363874
transform 1 0 972 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5599
timestamp 1680363874
transform 1 0 988 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1680363874
transform 1 0 996 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5075
timestamp 1680363874
transform 1 0 988 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1680363874
transform 1 0 1004 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1680363874
transform 1 0 1020 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5601
timestamp 1680363874
transform 1 0 1052 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1680363874
transform 1 0 1036 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_5077
timestamp 1680363874
transform 1 0 1044 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5436
timestamp 1680363874
transform 1 0 1068 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4972
timestamp 1680363874
transform 1 0 1100 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1680363874
transform 1 0 1116 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5614
timestamp 1680363874
transform 1 0 1116 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4973
timestamp 1680363874
transform 1 0 1140 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5514
timestamp 1680363874
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1680363874
transform 1 0 1148 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5060
timestamp 1680363874
transform 1 0 1196 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5515
timestamp 1680363874
transform 1 0 1220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1680363874
transform 1 0 1212 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4998
timestamp 1680363874
transform 1 0 1236 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5603
timestamp 1680363874
transform 1 0 1236 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5061
timestamp 1680363874
transform 1 0 1228 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5437
timestamp 1680363874
transform 1 0 1284 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4939
timestamp 1680363874
transform 1 0 1308 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5516
timestamp 1680363874
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5017
timestamp 1680363874
transform 1 0 1300 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1680363874
transform 1 0 1340 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1680363874
transform 1 0 1364 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1680363874
transform 1 0 1380 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5438
timestamp 1680363874
transform 1 0 1348 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4999
timestamp 1680363874
transform 1 0 1332 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1680363874
transform 1 0 1356 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5439
timestamp 1680363874
transform 1 0 1364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1680363874
transform 1 0 1380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1680363874
transform 1 0 1356 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5000
timestamp 1680363874
transform 1 0 1380 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5518
timestamp 1680363874
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5018
timestamp 1680363874
transform 1 0 1356 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1680363874
transform 1 0 1388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1680363874
transform 1 0 1444 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5441
timestamp 1680363874
transform 1 0 1444 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4942
timestamp 1680363874
transform 1 0 1532 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5519
timestamp 1680363874
transform 1 0 1468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1680363874
transform 1 0 1524 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5062
timestamp 1680363874
transform 1 0 1492 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1680363874
transform 1 0 1508 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5442
timestamp 1680363874
transform 1 0 1548 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4976
timestamp 1680363874
transform 1 0 1596 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1680363874
transform 1 0 1644 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5521
timestamp 1680363874
transform 1 0 1596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1680363874
transform 1 0 1628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1680363874
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5063
timestamp 1680363874
transform 1 0 1564 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1680363874
transform 1 0 1636 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5443
timestamp 1680363874
transform 1 0 1652 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_5079
timestamp 1680363874
transform 1 0 1660 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1680363874
transform 1 0 1676 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1680363874
transform 1 0 1684 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5444
timestamp 1680363874
transform 1 0 1692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1680363874
transform 1 0 1700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1680363874
transform 1 0 1716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1680363874
transform 1 0 1716 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5021
timestamp 1680363874
transform 1 0 1716 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5415
timestamp 1680363874
transform 1 0 1772 0 1 2155
box -2 -2 2 2
use M3_M2  M3_M2_4924
timestamp 1680363874
transform 1 0 1788 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5446
timestamp 1680363874
transform 1 0 1780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1680363874
transform 1 0 1796 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4978
timestamp 1680363874
transform 1 0 1804 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5448
timestamp 1680363874
transform 1 0 1812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1680363874
transform 1 0 1788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1680363874
transform 1 0 1804 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4906
timestamp 1680363874
transform 1 0 1932 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1680363874
transform 1 0 1884 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5449
timestamp 1680363874
transform 1 0 1932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1680363874
transform 1 0 1852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1680363874
transform 1 0 1884 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5080
timestamp 1680363874
transform 1 0 1852 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1680363874
transform 1 0 1876 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1680363874
transform 1 0 1892 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1680363874
transform 1 0 1924 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1680363874
transform 1 0 1972 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5450
timestamp 1680363874
transform 1 0 1956 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4980
timestamp 1680363874
transform 1 0 2004 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1680363874
transform 1 0 1956 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5530
timestamp 1680363874
transform 1 0 2004 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4925
timestamp 1680363874
transform 1 0 2116 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1680363874
transform 1 0 2092 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5451
timestamp 1680363874
transform 1 0 2092 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4981
timestamp 1680363874
transform 1 0 2100 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5452
timestamp 1680363874
transform 1 0 2108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1680363874
transform 1 0 2084 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5002
timestamp 1680363874
transform 1 0 2092 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5532
timestamp 1680363874
transform 1 0 2100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1680363874
transform 1 0 2116 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5022
timestamp 1680363874
transform 1 0 2084 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1680363874
transform 1 0 2132 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5453
timestamp 1680363874
transform 1 0 2156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1680363874
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4947
timestamp 1680363874
transform 1 0 2212 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5455
timestamp 1680363874
transform 1 0 2196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1680363874
transform 1 0 2212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1680363874
transform 1 0 2220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1680363874
transform 1 0 2204 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5024
timestamp 1680363874
transform 1 0 2204 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1680363874
transform 1 0 2220 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1680363874
transform 1 0 2228 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1680363874
transform 1 0 2244 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5535
timestamp 1680363874
transform 1 0 2252 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4926
timestamp 1680363874
transform 1 0 2300 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1680363874
transform 1 0 2300 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5536
timestamp 1680363874
transform 1 0 2284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1680363874
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1680363874
transform 1 0 2308 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5064
timestamp 1680363874
transform 1 0 2276 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1680363874
transform 1 0 2316 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5458
timestamp 1680363874
transform 1 0 2340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1680363874
transform 1 0 2348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1680363874
transform 1 0 2364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1680363874
transform 1 0 2332 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4984
timestamp 1680363874
transform 1 0 2372 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5540
timestamp 1680363874
transform 1 0 2356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1680363874
transform 1 0 2372 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5026
timestamp 1680363874
transform 1 0 2348 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1680363874
transform 1 0 2348 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1680363874
transform 1 0 2404 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5542
timestamp 1680363874
transform 1 0 2420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1680363874
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5084
timestamp 1680363874
transform 1 0 2412 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5461
timestamp 1680363874
transform 1 0 2452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1680363874
transform 1 0 2484 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1680363874
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5027
timestamp 1680363874
transform 1 0 2516 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1680363874
transform 1 0 2500 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5616
timestamp 1680363874
transform 1 0 2508 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1680363874
transform 1 0 2516 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4985
timestamp 1680363874
transform 1 0 2548 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1680363874
transform 1 0 2540 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5545
timestamp 1680363874
transform 1 0 2572 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5085
timestamp 1680363874
transform 1 0 2572 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1680363874
transform 1 0 2580 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5462
timestamp 1680363874
transform 1 0 2588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1680363874
transform 1 0 2588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5046
timestamp 1680363874
transform 1 0 2588 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1680363874
transform 1 0 2604 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5547
timestamp 1680363874
transform 1 0 2652 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1680363874
transform 1 0 2644 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5029
timestamp 1680363874
transform 1 0 2652 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5606
timestamp 1680363874
transform 1 0 2668 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1680363874
transform 1 0 2676 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5047
timestamp 1680363874
transform 1 0 2644 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5618
timestamp 1680363874
transform 1 0 2660 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1680363874
transform 1 0 2692 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5030
timestamp 1680363874
transform 1 0 2692 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5619
timestamp 1680363874
transform 1 0 2684 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_5086
timestamp 1680363874
transform 1 0 2684 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5608
timestamp 1680363874
transform 1 0 2740 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5048
timestamp 1680363874
transform 1 0 2740 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1680363874
transform 1 0 2804 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5463
timestamp 1680363874
transform 1 0 2756 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4951
timestamp 1680363874
transform 1 0 2844 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5464
timestamp 1680363874
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1680363874
transform 1 0 2796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1680363874
transform 1 0 2836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1680363874
transform 1 0 2852 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5049
timestamp 1680363874
transform 1 0 2852 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5552
timestamp 1680363874
transform 1 0 2876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1680363874
transform 1 0 2932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1680363874
transform 1 0 2948 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4907
timestamp 1680363874
transform 1 0 2972 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1680363874
transform 1 0 3044 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1680363874
transform 1 0 3052 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5466
timestamp 1680363874
transform 1 0 3052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1680363874
transform 1 0 2972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1680363874
transform 1 0 3028 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5067
timestamp 1680363874
transform 1 0 3076 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1680363874
transform 1 0 3092 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1680363874
transform 1 0 3116 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5467
timestamp 1680363874
transform 1 0 3116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1680363874
transform 1 0 3108 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4986
timestamp 1680363874
transform 1 0 3132 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1680363874
transform 1 0 3156 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5556
timestamp 1680363874
transform 1 0 3132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1680363874
transform 1 0 3148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1680363874
transform 1 0 3156 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5068
timestamp 1680363874
transform 1 0 3148 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1680363874
transform 1 0 3196 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5468
timestamp 1680363874
transform 1 0 3188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1680363874
transform 1 0 3196 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_5031
timestamp 1680363874
transform 1 0 3188 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5559
timestamp 1680363874
transform 1 0 3220 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5032
timestamp 1680363874
transform 1 0 3220 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5420
timestamp 1680363874
transform 1 0 3244 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_5004
timestamp 1680363874
transform 1 0 3236 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1680363874
transform 1 0 3260 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1680363874
transform 1 0 3284 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5470
timestamp 1680363874
transform 1 0 3292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1680363874
transform 1 0 3284 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5033
timestamp 1680363874
transform 1 0 3276 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1680363874
transform 1 0 3324 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1680363874
transform 1 0 3356 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5561
timestamp 1680363874
transform 1 0 3388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5034
timestamp 1680363874
transform 1 0 3380 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1680363874
transform 1 0 3412 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5471
timestamp 1680363874
transform 1 0 3412 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4990
timestamp 1680363874
transform 1 0 3420 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1680363874
transform 1 0 3444 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5562
timestamp 1680363874
transform 1 0 3444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1680363874
transform 1 0 3460 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1680363874
transform 1 0 3476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1680363874
transform 1 0 3476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1680363874
transform 1 0 3484 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5050
timestamp 1680363874
transform 1 0 3500 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5473
timestamp 1680363874
transform 1 0 3524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1680363874
transform 1 0 3532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1680363874
transform 1 0 3556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5035
timestamp 1680363874
transform 1 0 3556 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1680363874
transform 1 0 3548 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1680363874
transform 1 0 3588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1680363874
transform 1 0 3612 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1680363874
transform 1 0 3644 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5474
timestamp 1680363874
transform 1 0 3604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1680363874
transform 1 0 3612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1680363874
transform 1 0 3628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1680363874
transform 1 0 3636 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_5005
timestamp 1680363874
transform 1 0 3596 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5567
timestamp 1680363874
transform 1 0 3620 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5052
timestamp 1680363874
transform 1 0 3628 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1680363874
transform 1 0 3644 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5568
timestamp 1680363874
transform 1 0 3652 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5069
timestamp 1680363874
transform 1 0 3668 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5478
timestamp 1680363874
transform 1 0 3812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1680363874
transform 1 0 3724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1680363874
transform 1 0 3732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1680363874
transform 1 0 3764 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5036
timestamp 1680363874
transform 1 0 3724 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1680363874
transform 1 0 3764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1680363874
transform 1 0 3732 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5572
timestamp 1680363874
transform 1 0 3844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1680363874
transform 1 0 3916 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4991
timestamp 1680363874
transform 1 0 3972 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5480
timestamp 1680363874
transform 1 0 3980 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4992
timestamp 1680363874
transform 1 0 3996 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5573
timestamp 1680363874
transform 1 0 3988 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1680363874
transform 1 0 4028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1680363874
transform 1 0 4036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1680363874
transform 1 0 4052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1680363874
transform 1 0 4068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1680363874
transform 1 0 4044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1680363874
transform 1 0 4060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1680363874
transform 1 0 4068 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5087
timestamp 1680363874
transform 1 0 4076 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1680363874
transform 1 0 4164 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5485
timestamp 1680363874
transform 1 0 4164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1680363874
transform 1 0 4140 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5088
timestamp 1680363874
transform 1 0 4156 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1680363874
transform 1 0 4212 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5486
timestamp 1680363874
transform 1 0 4212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1680363874
transform 1 0 4236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1680363874
transform 1 0 4324 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4910
timestamp 1680363874
transform 1 0 4348 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1680363874
transform 1 0 4372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1680363874
transform 1 0 4436 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1680363874
transform 1 0 4476 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1680363874
transform 1 0 4380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1680363874
transform 1 0 4468 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5487
timestamp 1680363874
transform 1 0 4380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1680363874
transform 1 0 4468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1680363874
transform 1 0 4428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1680363874
transform 1 0 4460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1680363874
transform 1 0 4468 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5038
timestamp 1680363874
transform 1 0 4428 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1680363874
transform 1 0 4468 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1680363874
transform 1 0 4460 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1680363874
transform 1 0 4508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1680363874
transform 1 0 4500 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1680363874
transform 1 0 4492 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1680363874
transform 1 0 4524 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5422
timestamp 1680363874
transform 1 0 4524 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1680363874
transform 1 0 4540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1680363874
transform 1 0 4540 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4931
timestamp 1680363874
transform 1 0 4580 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5490
timestamp 1680363874
transform 1 0 4564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1680363874
transform 1 0 4580 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1680363874
transform 1 0 4572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1680363874
transform 1 0 4604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1680363874
transform 1 0 4620 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_5007
timestamp 1680363874
transform 1 0 4620 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5610
timestamp 1680363874
transform 1 0 4620 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_5054
timestamp 1680363874
transform 1 0 4620 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5493
timestamp 1680363874
transform 1 0 4636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1680363874
transform 1 0 4652 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1680363874
transform 1 0 4660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1680363874
transform 1 0 4644 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5008
timestamp 1680363874
transform 1 0 4652 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5587
timestamp 1680363874
transform 1 0 4660 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5055
timestamp 1680363874
transform 1 0 4676 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5496
timestamp 1680363874
transform 1 0 4788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1680363874
transform 1 0 4700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1680363874
transform 1 0 4708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1680363874
transform 1 0 4756 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_5040
timestamp 1680363874
transform 1 0 4700 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1680363874
transform 1 0 4788 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1680363874
transform 1 0 4756 0 1 2115
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_52
timestamp 1680363874
transform 1 0 24 0 1 2070
box -10 -3 10 3
use FILL  FILL_5867
timestamp 1680363874
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5869
timestamp 1680363874
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5871
timestamp 1680363874
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5872
timestamp 1680363874
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5873
timestamp 1680363874
transform 1 0 104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5874
timestamp 1680363874
transform 1 0 112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5875
timestamp 1680363874
transform 1 0 120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5882
timestamp 1680363874
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_28
timestamp 1680363874
transform -1 0 168 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5883
timestamp 1680363874
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5884
timestamp 1680363874
transform 1 0 176 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_378
timestamp 1680363874
transform 1 0 184 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5885
timestamp 1680363874
transform 1 0 200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5887
timestamp 1680363874
transform 1 0 208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5889
timestamp 1680363874
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5895
timestamp 1680363874
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_58
timestamp 1680363874
transform -1 0 256 0 -1 2170
box -8 -3 32 105
use NAND3X1  NAND3X1_30
timestamp 1680363874
transform 1 0 256 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5896
timestamp 1680363874
transform 1 0 288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5898
timestamp 1680363874
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5900
timestamp 1680363874
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5904
timestamp 1680363874
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_135
timestamp 1680363874
transform -1 0 352 0 -1 2170
box -8 -3 34 105
use FILL  FILL_5905
timestamp 1680363874
transform 1 0 352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5906
timestamp 1680363874
transform 1 0 360 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_379
timestamp 1680363874
transform 1 0 368 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5925
timestamp 1680363874
transform 1 0 384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5926
timestamp 1680363874
transform 1 0 392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5927
timestamp 1680363874
transform 1 0 400 0 -1 2170
box -8 -3 16 105
use AOI21X1  AOI21X1_13
timestamp 1680363874
transform 1 0 408 0 -1 2170
box -7 -3 39 105
use FILL  FILL_5928
timestamp 1680363874
transform 1 0 440 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5089
timestamp 1680363874
transform 1 0 564 0 1 2075
box -3 -3 3 3
use FAX1  FAX1_13
timestamp 1680363874
transform -1 0 568 0 -1 2170
box -5 -3 126 105
use FILL  FILL_5929
timestamp 1680363874
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5931
timestamp 1680363874
transform 1 0 576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5933
timestamp 1680363874
transform 1 0 584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5935
timestamp 1680363874
transform 1 0 592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5937
timestamp 1680363874
transform 1 0 600 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_42
timestamp 1680363874
transform 1 0 608 0 -1 2170
box -8 -3 32 105
use FILL  FILL_5942
timestamp 1680363874
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5944
timestamp 1680363874
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5946
timestamp 1680363874
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5948
timestamp 1680363874
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5950
timestamp 1680363874
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5952
timestamp 1680363874
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_43
timestamp 1680363874
transform 1 0 680 0 -1 2170
box -8 -3 32 105
use FILL  FILL_5957
timestamp 1680363874
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5959
timestamp 1680363874
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5961
timestamp 1680363874
transform 1 0 720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5963
timestamp 1680363874
transform 1 0 728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5969
timestamp 1680363874
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5970
timestamp 1680363874
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_44
timestamp 1680363874
transform 1 0 752 0 -1 2170
box -8 -3 32 105
use FILL  FILL_5971
timestamp 1680363874
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5972
timestamp 1680363874
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5973
timestamp 1680363874
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5974
timestamp 1680363874
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5975
timestamp 1680363874
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5976
timestamp 1680363874
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FAX1  FAX1_15
timestamp 1680363874
transform 1 0 824 0 -1 2170
box -5 -3 126 105
use FILL  FILL_5977
timestamp 1680363874
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5979
timestamp 1680363874
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5981
timestamp 1680363874
transform 1 0 960 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1680363874
transform 1 0 968 0 -1 2170
box -8 -3 32 105
use FILL  FILL_5983
timestamp 1680363874
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5985
timestamp 1680363874
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5987
timestamp 1680363874
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5993
timestamp 1680363874
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_32
timestamp 1680363874
transform -1 0 1056 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5994
timestamp 1680363874
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5995
timestamp 1680363874
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5090
timestamp 1680363874
transform 1 0 1084 0 1 2075
box -3 -3 3 3
use FILL  FILL_5996
timestamp 1680363874
transform 1 0 1072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5997
timestamp 1680363874
transform 1 0 1080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5999
timestamp 1680363874
transform 1 0 1088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6001
timestamp 1680363874
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6003
timestamp 1680363874
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6005
timestamp 1680363874
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_380
timestamp 1680363874
transform 1 0 1120 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6008
timestamp 1680363874
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6009
timestamp 1680363874
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6010
timestamp 1680363874
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6011
timestamp 1680363874
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6013
timestamp 1680363874
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6015
timestamp 1680363874
transform 1 0 1176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6017
timestamp 1680363874
transform 1 0 1184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6019
timestamp 1680363874
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6021
timestamp 1680363874
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_34
timestamp 1680363874
transform 1 0 1208 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6027
timestamp 1680363874
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6029
timestamp 1680363874
transform 1 0 1248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6031
timestamp 1680363874
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6033
timestamp 1680363874
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6035
timestamp 1680363874
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_381
timestamp 1680363874
transform 1 0 1280 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6039
timestamp 1680363874
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6041
timestamp 1680363874
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6047
timestamp 1680363874
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6048
timestamp 1680363874
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6049
timestamp 1680363874
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6050
timestamp 1680363874
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_255
timestamp 1680363874
transform -1 0 1384 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6051
timestamp 1680363874
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6053
timestamp 1680363874
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6055
timestamp 1680363874
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6057
timestamp 1680363874
transform 1 0 1408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6059
timestamp 1680363874
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6061
timestamp 1680363874
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_325
timestamp 1680363874
transform 1 0 1432 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6068
timestamp 1680363874
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5091
timestamp 1680363874
transform 1 0 1548 0 1 2075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_326
timestamp 1680363874
transform 1 0 1536 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6077
timestamp 1680363874
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6078
timestamp 1680363874
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6079
timestamp 1680363874
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6081
timestamp 1680363874
transform 1 0 1656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6083
timestamp 1680363874
transform 1 0 1664 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_259
timestamp 1680363874
transform 1 0 1672 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6086
timestamp 1680363874
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6087
timestamp 1680363874
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6090
timestamp 1680363874
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6091
timestamp 1680363874
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6092
timestamp 1680363874
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6093
timestamp 1680363874
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6095
timestamp 1680363874
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6097
timestamp 1680363874
transform 1 0 1768 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_261
timestamp 1680363874
transform 1 0 1776 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6101
timestamp 1680363874
transform 1 0 1816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6102
timestamp 1680363874
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6103
timestamp 1680363874
transform 1 0 1832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6117
timestamp 1680363874
transform 1 0 1840 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_328
timestamp 1680363874
transform -1 0 1944 0 -1 2170
box -8 -3 104 105
use M3_M2  M3_M2_5092
timestamp 1680363874
transform 1 0 2004 0 1 2075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_329
timestamp 1680363874
transform 1 0 1944 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_387
timestamp 1680363874
transform 1 0 2040 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6118
timestamp 1680363874
transform 1 0 2056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6119
timestamp 1680363874
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6121
timestamp 1680363874
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6123
timestamp 1680363874
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_263
timestamp 1680363874
transform -1 0 2128 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6125
timestamp 1680363874
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6127
timestamp 1680363874
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6129
timestamp 1680363874
transform 1 0 2144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6131
timestamp 1680363874
transform 1 0 2152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6136
timestamp 1680363874
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6137
timestamp 1680363874
transform 1 0 2168 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_264
timestamp 1680363874
transform 1 0 2176 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6138
timestamp 1680363874
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6140
timestamp 1680363874
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6146
timestamp 1680363874
transform 1 0 2232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6147
timestamp 1680363874
transform 1 0 2240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6148
timestamp 1680363874
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6149
timestamp 1680363874
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_198
timestamp 1680363874
transform 1 0 2264 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6150
timestamp 1680363874
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6154
timestamp 1680363874
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6155
timestamp 1680363874
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6156
timestamp 1680363874
transform 1 0 2328 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_199
timestamp 1680363874
transform 1 0 2336 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6157
timestamp 1680363874
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6158
timestamp 1680363874
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6160
timestamp 1680363874
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6162
timestamp 1680363874
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6164
timestamp 1680363874
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_20
timestamp 1680363874
transform -1 0 2448 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6169
timestamp 1680363874
transform 1 0 2448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6170
timestamp 1680363874
transform 1 0 2456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6171
timestamp 1680363874
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6172
timestamp 1680363874
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6173
timestamp 1680363874
transform 1 0 2480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6174
timestamp 1680363874
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_36
timestamp 1680363874
transform -1 0 2528 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6175
timestamp 1680363874
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6176
timestamp 1680363874
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6177
timestamp 1680363874
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6178
timestamp 1680363874
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5093
timestamp 1680363874
transform 1 0 2572 0 1 2075
box -3 -3 3 3
use FILL  FILL_6179
timestamp 1680363874
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_392
timestamp 1680363874
transform 1 0 2568 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_393
timestamp 1680363874
transform 1 0 2584 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6180
timestamp 1680363874
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6181
timestamp 1680363874
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6182
timestamp 1680363874
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5094
timestamp 1680363874
transform 1 0 2636 0 1 2075
box -3 -3 3 3
use FILL  FILL_6183
timestamp 1680363874
transform 1 0 2624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6184
timestamp 1680363874
transform 1 0 2632 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_37
timestamp 1680363874
transform 1 0 2640 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6185
timestamp 1680363874
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_38
timestamp 1680363874
transform 1 0 2680 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6186
timestamp 1680363874
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6188
timestamp 1680363874
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6190
timestamp 1680363874
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6198
timestamp 1680363874
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_332
timestamp 1680363874
transform 1 0 2744 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6199
timestamp 1680363874
transform 1 0 2840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6201
timestamp 1680363874
transform 1 0 2848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6203
timestamp 1680363874
transform 1 0 2856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6205
timestamp 1680363874
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6210
timestamp 1680363874
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6211
timestamp 1680363874
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6212
timestamp 1680363874
transform 1 0 2888 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_138
timestamp 1680363874
transform 1 0 2896 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6213
timestamp 1680363874
transform 1 0 2928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6215
timestamp 1680363874
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6217
timestamp 1680363874
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6219
timestamp 1680363874
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6227
timestamp 1680363874
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_333
timestamp 1680363874
transform -1 0 3064 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6228
timestamp 1680363874
transform 1 0 3064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6229
timestamp 1680363874
transform 1 0 3072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6231
timestamp 1680363874
transform 1 0 3080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6233
timestamp 1680363874
transform 1 0 3088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6235
timestamp 1680363874
transform 1 0 3096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6240
timestamp 1680363874
transform 1 0 3104 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5095
timestamp 1680363874
transform 1 0 3156 0 1 2075
box -3 -3 3 3
use AOI22X1  AOI22X1_200
timestamp 1680363874
transform -1 0 3152 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6241
timestamp 1680363874
transform 1 0 3152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6242
timestamp 1680363874
transform 1 0 3160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6244
timestamp 1680363874
transform 1 0 3168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6246
timestamp 1680363874
transform 1 0 3176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6248
timestamp 1680363874
transform 1 0 3184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6254
timestamp 1680363874
transform 1 0 3192 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_59
timestamp 1680363874
transform -1 0 3224 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6255
timestamp 1680363874
transform 1 0 3224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6257
timestamp 1680363874
transform 1 0 3232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6261
timestamp 1680363874
transform 1 0 3240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6262
timestamp 1680363874
transform 1 0 3248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6263
timestamp 1680363874
transform 1 0 3256 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_21
timestamp 1680363874
transform -1 0 3296 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6264
timestamp 1680363874
transform 1 0 3296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6266
timestamp 1680363874
transform 1 0 3304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6268
timestamp 1680363874
transform 1 0 3312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6270
timestamp 1680363874
transform 1 0 3320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6272
timestamp 1680363874
transform 1 0 3328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6274
timestamp 1680363874
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6279
timestamp 1680363874
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6280
timestamp 1680363874
transform 1 0 3352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6281
timestamp 1680363874
transform 1 0 3360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6282
timestamp 1680363874
transform 1 0 3368 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1680363874
transform 1 0 3376 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6283
timestamp 1680363874
transform 1 0 3408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6284
timestamp 1680363874
transform 1 0 3416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6285
timestamp 1680363874
transform 1 0 3424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6286
timestamp 1680363874
transform 1 0 3432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6287
timestamp 1680363874
transform 1 0 3440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6289
timestamp 1680363874
transform 1 0 3448 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1680363874
transform 1 0 3456 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6297
timestamp 1680363874
transform 1 0 3480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6298
timestamp 1680363874
transform 1 0 3488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6299
timestamp 1680363874
transform 1 0 3496 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_268
timestamp 1680363874
transform 1 0 3504 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6300
timestamp 1680363874
transform 1 0 3544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6302
timestamp 1680363874
transform 1 0 3552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6304
timestamp 1680363874
transform 1 0 3560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6306
timestamp 1680363874
transform 1 0 3568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6311
timestamp 1680363874
transform 1 0 3576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6312
timestamp 1680363874
transform 1 0 3584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6313
timestamp 1680363874
transform 1 0 3592 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_204
timestamp 1680363874
transform 1 0 3600 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6314
timestamp 1680363874
transform 1 0 3640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6320
timestamp 1680363874
transform 1 0 3648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6321
timestamp 1680363874
transform 1 0 3656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6322
timestamp 1680363874
transform 1 0 3664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6323
timestamp 1680363874
transform 1 0 3672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6324
timestamp 1680363874
transform 1 0 3680 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_396
timestamp 1680363874
transform 1 0 3688 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6325
timestamp 1680363874
transform 1 0 3704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6326
timestamp 1680363874
transform 1 0 3712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6327
timestamp 1680363874
transform 1 0 3720 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_336
timestamp 1680363874
transform -1 0 3824 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6328
timestamp 1680363874
transform 1 0 3824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6329
timestamp 1680363874
transform 1 0 3832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6330
timestamp 1680363874
transform 1 0 3840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6331
timestamp 1680363874
transform 1 0 3848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6332
timestamp 1680363874
transform 1 0 3856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6333
timestamp 1680363874
transform 1 0 3864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6334
timestamp 1680363874
transform 1 0 3872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6335
timestamp 1680363874
transform 1 0 3880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6336
timestamp 1680363874
transform 1 0 3888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6338
timestamp 1680363874
transform 1 0 3896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6340
timestamp 1680363874
transform 1 0 3904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6342
timestamp 1680363874
transform 1 0 3912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6347
timestamp 1680363874
transform 1 0 3920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6348
timestamp 1680363874
transform 1 0 3928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6349
timestamp 1680363874
transform 1 0 3936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6350
timestamp 1680363874
transform 1 0 3944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6351
timestamp 1680363874
transform 1 0 3952 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_269
timestamp 1680363874
transform 1 0 3960 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6352
timestamp 1680363874
transform 1 0 4000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6354
timestamp 1680363874
transform 1 0 4008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6364
timestamp 1680363874
transform 1 0 4016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6365
timestamp 1680363874
transform 1 0 4024 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5096
timestamp 1680363874
transform 1 0 4076 0 1 2075
box -3 -3 3 3
use OAI22X1  OAI22X1_270
timestamp 1680363874
transform -1 0 4072 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6366
timestamp 1680363874
transform 1 0 4072 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5097
timestamp 1680363874
transform 1 0 4124 0 1 2075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_338
timestamp 1680363874
transform -1 0 4176 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6367
timestamp 1680363874
transform 1 0 4176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6369
timestamp 1680363874
transform 1 0 4184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6371
timestamp 1680363874
transform 1 0 4192 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_340
timestamp 1680363874
transform 1 0 4200 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6374
timestamp 1680363874
transform 1 0 4296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6375
timestamp 1680363874
transform 1 0 4304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6377
timestamp 1680363874
transform 1 0 4312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6379
timestamp 1680363874
transform 1 0 4320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6389
timestamp 1680363874
transform 1 0 4328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6390
timestamp 1680363874
transform 1 0 4336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6391
timestamp 1680363874
transform 1 0 4344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6392
timestamp 1680363874
transform 1 0 4352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6393
timestamp 1680363874
transform 1 0 4360 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_341
timestamp 1680363874
transform 1 0 4368 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_398
timestamp 1680363874
transform 1 0 4464 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6394
timestamp 1680363874
transform 1 0 4480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6395
timestamp 1680363874
transform 1 0 4488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6396
timestamp 1680363874
transform 1 0 4496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6398
timestamp 1680363874
transform 1 0 4504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6400
timestamp 1680363874
transform 1 0 4512 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_63
timestamp 1680363874
transform 1 0 4520 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6405
timestamp 1680363874
transform 1 0 4544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6406
timestamp 1680363874
transform 1 0 4552 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_272
timestamp 1680363874
transform -1 0 4600 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6407
timestamp 1680363874
transform 1 0 4600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6408
timestamp 1680363874
transform 1 0 4608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6410
timestamp 1680363874
transform 1 0 4616 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_209
timestamp 1680363874
transform 1 0 4624 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6412
timestamp 1680363874
transform 1 0 4664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6414
timestamp 1680363874
transform 1 0 4672 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_400
timestamp 1680363874
transform 1 0 4680 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6428
timestamp 1680363874
transform 1 0 4696 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_342
timestamp 1680363874
transform -1 0 4800 0 -1 2170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_53
timestamp 1680363874
transform 1 0 4851 0 1 2070
box -10 -3 10 3
use M2_M1  M2_M1_5811
timestamp 1680363874
transform 1 0 100 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1680363874
transform 1 0 116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1680363874
transform 1 0 124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1680363874
transform 1 0 156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1680363874
transform 1 0 172 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1680363874
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1680363874
transform 1 0 236 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1680363874
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1680363874
transform 1 0 260 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5125
timestamp 1680363874
transform 1 0 292 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1680363874
transform 1 0 324 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5749
timestamp 1680363874
transform 1 0 324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1680363874
transform 1 0 340 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5098
timestamp 1680363874
transform 1 0 460 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1680363874
transform 1 0 380 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1680363874
transform 1 0 460 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5650
timestamp 1680363874
transform 1 0 452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1680363874
transform 1 0 460 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5109
timestamp 1680363874
transform 1 0 508 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1680363874
transform 1 0 516 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1680363874
transform 1 0 580 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1680363874
transform 1 0 596 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1680363874
transform 1 0 668 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5652
timestamp 1680363874
transform 1 0 508 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5173
timestamp 1680363874
transform 1 0 548 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5653
timestamp 1680363874
transform 1 0 564 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5174
timestamp 1680363874
transform 1 0 572 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5654
timestamp 1680363874
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1680363874
transform 1 0 676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1680363874
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1680363874
transform 1 0 484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1680363874
transform 1 0 572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1680363874
transform 1 0 364 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5206
timestamp 1680363874
transform 1 0 484 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1680363874
transform 1 0 548 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1680363874
transform 1 0 580 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1680363874
transform 1 0 628 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5815
timestamp 1680363874
transform 1 0 580 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5228
timestamp 1680363874
transform 1 0 612 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1680363874
transform 1 0 708 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5753
timestamp 1680363874
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1680363874
transform 1 0 708 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5112
timestamp 1680363874
transform 1 0 796 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1680363874
transform 1 0 780 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1680363874
transform 1 0 804 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1680363874
transform 1 0 828 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5656
timestamp 1680363874
transform 1 0 812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1680363874
transform 1 0 820 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5193
timestamp 1680363874
transform 1 0 772 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1680363874
transform 1 0 860 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1680363874
transform 1 0 852 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5658
timestamp 1680363874
transform 1 0 836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1680363874
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1680363874
transform 1 0 860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1680363874
transform 1 0 828 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1680363874
transform 1 0 724 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5133
timestamp 1680363874
transform 1 0 876 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1680363874
transform 1 0 868 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5756
timestamp 1680363874
transform 1 0 876 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5229
timestamp 1680363874
transform 1 0 860 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1680363874
transform 1 0 996 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1680363874
transform 1 0 1044 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1680363874
transform 1 0 972 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1680363874
transform 1 0 1012 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1680363874
transform 1 0 1060 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5661
timestamp 1680363874
transform 1 0 1012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1680363874
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5195
timestamp 1680363874
transform 1 0 1004 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5662
timestamp 1680363874
transform 1 0 1068 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5115
timestamp 1680363874
transform 1 0 1124 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1680363874
transform 1 0 1132 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5663
timestamp 1680363874
transform 1 0 1116 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5175
timestamp 1680363874
transform 1 0 1124 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5664
timestamp 1680363874
transform 1 0 1132 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5155
timestamp 1680363874
transform 1 0 1148 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5758
timestamp 1680363874
transform 1 0 1108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1680363874
transform 1 0 1124 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1680363874
transform 1 0 1140 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1680363874
transform 1 0 1148 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5136
timestamp 1680363874
transform 1 0 1172 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5665
timestamp 1680363874
transform 1 0 1188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1680363874
transform 1 0 1228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1680363874
transform 1 0 1244 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5137
timestamp 1680363874
transform 1 0 1364 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5668
timestamp 1680363874
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1680363874
transform 1 0 1340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1680363874
transform 1 0 1276 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5208
timestamp 1680363874
transform 1 0 1276 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5745
timestamp 1680363874
transform 1 0 1364 0 1 2007
box -2 -2 2 2
use M3_M2  M3_M2_5230
timestamp 1680363874
transform 1 0 1292 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1680363874
transform 1 0 1364 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1680363874
transform 1 0 1380 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1680363874
transform 1 0 1444 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1680363874
transform 1 0 1404 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5670
timestamp 1680363874
transform 1 0 1428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1680363874
transform 1 0 1404 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5209
timestamp 1680363874
transform 1 0 1436 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5629
timestamp 1680363874
transform 1 0 1532 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1680363874
transform 1 0 1524 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5210
timestamp 1680363874
transform 1 0 1524 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1680363874
transform 1 0 1572 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5622
timestamp 1680363874
transform 1 0 1564 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1680363874
transform 1 0 1572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1680363874
transform 1 0 1596 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1680363874
transform 1 0 1620 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5110
timestamp 1680363874
transform 1 0 1660 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1680363874
transform 1 0 1668 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5673
timestamp 1680363874
transform 1 0 1668 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5140
timestamp 1680363874
transform 1 0 1700 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5674
timestamp 1680363874
transform 1 0 1692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1680363874
transform 1 0 1708 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5211
timestamp 1680363874
transform 1 0 1684 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5765
timestamp 1680363874
transform 1 0 1716 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5212
timestamp 1680363874
transform 1 0 1716 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1680363874
transform 1 0 1740 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5631
timestamp 1680363874
transform 1 0 1748 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1680363874
transform 1 0 1740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1680363874
transform 1 0 1748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1680363874
transform 1 0 1772 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5232
timestamp 1680363874
transform 1 0 1772 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1680363874
transform 1 0 1812 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1680363874
transform 1 0 1804 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5678
timestamp 1680363874
transform 1 0 1812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1680363874
transform 1 0 1804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1680363874
transform 1 0 1820 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5213
timestamp 1680363874
transform 1 0 1804 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5620
timestamp 1680363874
transform 1 0 1844 0 1 2045
box -2 -2 2 2
use M3_M2  M3_M2_5160
timestamp 1680363874
transform 1 0 1836 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5679
timestamp 1680363874
transform 1 0 1836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1680363874
transform 1 0 1860 0 1 2045
box -2 -2 2 2
use M3_M2  M3_M2_5176
timestamp 1680363874
transform 1 0 1852 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5768
timestamp 1680363874
transform 1 0 1852 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5233
timestamp 1680363874
transform 1 0 1844 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5680
timestamp 1680363874
transform 1 0 1876 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5214
timestamp 1680363874
transform 1 0 1868 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1680363874
transform 1 0 1868 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1680363874
transform 1 0 1932 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5633
timestamp 1680363874
transform 1 0 1980 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1680363874
transform 1 0 1940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1680363874
transform 1 0 1972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1680363874
transform 1 0 1892 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5196
timestamp 1680363874
transform 1 0 1940 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1680363874
transform 1 0 1916 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1680363874
transform 1 0 1988 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5683
timestamp 1680363874
transform 1 0 2036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1680363874
transform 1 0 2068 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1680363874
transform 1 0 2052 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1680363874
transform 1 0 2060 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5161
timestamp 1680363874
transform 1 0 2068 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1680363874
transform 1 0 2100 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5624
timestamp 1680363874
transform 1 0 2092 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1680363874
transform 1 0 2100 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1680363874
transform 1 0 2084 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5198
timestamp 1680363874
transform 1 0 2092 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1680363874
transform 1 0 2196 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1680363874
transform 1 0 2132 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5685
timestamp 1680363874
transform 1 0 2180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1680363874
transform 1 0 2132 0 1 2007
box -2 -2 2 2
use M3_M2  M3_M2_5119
timestamp 1680363874
transform 1 0 2236 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5637
timestamp 1680363874
transform 1 0 2236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1680363874
transform 1 0 2228 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5179
timestamp 1680363874
transform 1 0 2276 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1680363874
transform 1 0 2300 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5625
timestamp 1680363874
transform 1 0 2300 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1680363874
transform 1 0 2308 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1680363874
transform 1 0 2292 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5180
timestamp 1680363874
transform 1 0 2308 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5626
timestamp 1680363874
transform 1 0 2356 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1680363874
transform 1 0 2356 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1680363874
transform 1 0 2380 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1680363874
transform 1 0 2396 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1680363874
transform 1 0 2404 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5102
timestamp 1680363874
transform 1 0 2428 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5689
timestamp 1680363874
transform 1 0 2444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1680363874
transform 1 0 2460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1680363874
transform 1 0 2452 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5103
timestamp 1680363874
transform 1 0 2516 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5691
timestamp 1680363874
transform 1 0 2500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1680363874
transform 1 0 2516 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1680363874
transform 1 0 2524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1680363874
transform 1 0 2532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1680363874
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5215
timestamp 1680363874
transform 1 0 2508 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5772
timestamp 1680363874
transform 1 0 2540 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5104
timestamp 1680363874
transform 1 0 2588 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5628
timestamp 1680363874
transform 1 0 2588 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1680363874
transform 1 0 2580 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1680363874
transform 1 0 2596 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1680363874
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1680363874
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1680363874
transform 1 0 2612 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5236
timestamp 1680363874
transform 1 0 2604 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5774
timestamp 1680363874
transform 1 0 2628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1680363874
transform 1 0 2692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1680363874
transform 1 0 2668 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5120
timestamp 1680363874
transform 1 0 2772 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5698
timestamp 1680363874
transform 1 0 2764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1680363874
transform 1 0 2756 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5216
timestamp 1680363874
transform 1 0 2756 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5699
timestamp 1680363874
transform 1 0 2804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1680363874
transform 1 0 2820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1680363874
transform 1 0 2836 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5217
timestamp 1680363874
transform 1 0 2828 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5701
timestamp 1680363874
transform 1 0 2844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1680363874
transform 1 0 2876 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5181
timestamp 1680363874
transform 1 0 2884 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1680363874
transform 1 0 2900 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5703
timestamp 1680363874
transform 1 0 2892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1680363874
transform 1 0 2908 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5218
timestamp 1680363874
transform 1 0 2908 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5643
timestamp 1680363874
transform 1 0 2932 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5237
timestamp 1680363874
transform 1 0 2972 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1680363874
transform 1 0 2988 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5779
timestamp 1680363874
transform 1 0 2996 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5219
timestamp 1680363874
transform 1 0 2988 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5817
timestamp 1680363874
transform 1 0 3012 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1680363874
transform 1 0 3028 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5141
timestamp 1680363874
transform 1 0 3108 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5704
timestamp 1680363874
transform 1 0 3108 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5183
timestamp 1680363874
transform 1 0 3116 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5780
timestamp 1680363874
transform 1 0 3116 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5184
timestamp 1680363874
transform 1 0 3132 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1680363874
transform 1 0 3164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1680363874
transform 1 0 3164 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5705
timestamp 1680363874
transform 1 0 3140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1680363874
transform 1 0 3156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1680363874
transform 1 0 3164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1680363874
transform 1 0 3132 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5220
timestamp 1680363874
transform 1 0 3132 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5782
timestamp 1680363874
transform 1 0 3172 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5185
timestamp 1680363874
transform 1 0 3188 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5818
timestamp 1680363874
transform 1 0 3188 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5106
timestamp 1680363874
transform 1 0 3228 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5708
timestamp 1680363874
transform 1 0 3220 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5186
timestamp 1680363874
transform 1 0 3228 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5709
timestamp 1680363874
transform 1 0 3236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1680363874
transform 1 0 3244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1680363874
transform 1 0 3212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1680363874
transform 1 0 3228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1680363874
transform 1 0 3308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1680363874
transform 1 0 3324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1680363874
transform 1 0 3300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1680363874
transform 1 0 3324 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5221
timestamp 1680363874
transform 1 0 3300 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5713
timestamp 1680363874
transform 1 0 3348 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5162
timestamp 1680363874
transform 1 0 3364 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1680363874
transform 1 0 3364 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5714
timestamp 1680363874
transform 1 0 3388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1680363874
transform 1 0 3396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1680363874
transform 1 0 3412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1680363874
transform 1 0 3404 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5199
timestamp 1680363874
transform 1 0 3412 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5788
timestamp 1680363874
transform 1 0 3420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1680363874
transform 1 0 3428 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5222
timestamp 1680363874
transform 1 0 3428 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5717
timestamp 1680363874
transform 1 0 3452 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5200
timestamp 1680363874
transform 1 0 3492 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5819
timestamp 1680363874
transform 1 0 3492 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5239
timestamp 1680363874
transform 1 0 3484 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1680363874
transform 1 0 3516 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1680363874
transform 1 0 3532 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5718
timestamp 1680363874
transform 1 0 3532 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5201
timestamp 1680363874
transform 1 0 3524 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1680363874
transform 1 0 3580 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1680363874
transform 1 0 3620 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5719
timestamp 1680363874
transform 1 0 3580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1680363874
transform 1 0 3620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1680363874
transform 1 0 3676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1680363874
transform 1 0 3572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5223
timestamp 1680363874
transform 1 0 3572 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5791
timestamp 1680363874
transform 1 0 3596 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5224
timestamp 1680363874
transform 1 0 3620 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1680363874
transform 1 0 3772 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5722
timestamp 1680363874
transform 1 0 3756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1680363874
transform 1 0 3772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1680363874
transform 1 0 3788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1680363874
transform 1 0 3764 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5240
timestamp 1680363874
transform 1 0 3756 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5725
timestamp 1680363874
transform 1 0 3844 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5167
timestamp 1680363874
transform 1 0 3884 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5726
timestamp 1680363874
transform 1 0 3884 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1680363874
transform 1 0 3852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1680363874
transform 1 0 3860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1680363874
transform 1 0 3876 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1680363874
transform 1 0 3892 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5241
timestamp 1680363874
transform 1 0 3884 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1680363874
transform 1 0 3908 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1680363874
transform 1 0 3972 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1680363874
transform 1 0 3988 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1680363874
transform 1 0 3980 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5797
timestamp 1680363874
transform 1 0 3972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1680363874
transform 1 0 3996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1680363874
transform 1 0 4068 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5225
timestamp 1680363874
transform 1 0 4060 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1680363874
transform 1 0 4092 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1680363874
transform 1 0 4108 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5728
timestamp 1680363874
transform 1 0 4092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1680363874
transform 1 0 4108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1680363874
transform 1 0 4124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1680363874
transform 1 0 4140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1680363874
transform 1 0 4148 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5242
timestamp 1680363874
transform 1 0 4148 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1680363874
transform 1 0 4164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1680363874
transform 1 0 4172 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5800
timestamp 1680363874
transform 1 0 4172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1680363874
transform 1 0 4180 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5226
timestamp 1680363874
transform 1 0 4180 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1680363874
transform 1 0 4228 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1680363874
transform 1 0 4220 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1680363874
transform 1 0 4244 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5732
timestamp 1680363874
transform 1 0 4228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1680363874
transform 1 0 4236 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5144
timestamp 1680363874
transform 1 0 4276 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5734
timestamp 1680363874
transform 1 0 4276 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5190
timestamp 1680363874
transform 1 0 4324 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5735
timestamp 1680363874
transform 1 0 4332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1680363874
transform 1 0 4348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1680363874
transform 1 0 4316 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1680363874
transform 1 0 4324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1680363874
transform 1 0 4340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1680363874
transform 1 0 4348 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5227
timestamp 1680363874
transform 1 0 4340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1680363874
transform 1 0 4332 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1680363874
transform 1 0 4364 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5737
timestamp 1680363874
transform 1 0 4364 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5244
timestamp 1680363874
transform 1 0 4404 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5738
timestamp 1680363874
transform 1 0 4436 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5107
timestamp 1680363874
transform 1 0 4452 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1680363874
transform 1 0 4476 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1680363874
transform 1 0 4484 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5739
timestamp 1680363874
transform 1 0 4452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1680363874
transform 1 0 4468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1680363874
transform 1 0 4484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1680363874
transform 1 0 4452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1680363874
transform 1 0 4460 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5202
timestamp 1680363874
transform 1 0 4468 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5808
timestamp 1680363874
transform 1 0 4492 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5146
timestamp 1680363874
transform 1 0 4660 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1680363874
transform 1 0 4652 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5809
timestamp 1680363874
transform 1 0 4660 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5147
timestamp 1680363874
transform 1 0 4692 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5742
timestamp 1680363874
transform 1 0 4700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1680363874
transform 1 0 4756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1680363874
transform 1 0 4796 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5204
timestamp 1680363874
transform 1 0 4700 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5810
timestamp 1680363874
transform 1 0 4716 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5205
timestamp 1680363874
transform 1 0 4756 0 1 2005
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_54
timestamp 1680363874
transform 1 0 48 0 1 1970
box -10 -3 10 3
use FILL  FILL_6429
timestamp 1680363874
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_6430
timestamp 1680363874
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_6431
timestamp 1680363874
transform 1 0 88 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_64
timestamp 1680363874
transform 1 0 96 0 1 1970
box -8 -3 32 105
use FILL  FILL_6432
timestamp 1680363874
transform 1 0 120 0 1 1970
box -8 -3 16 105
use FILL  FILL_6433
timestamp 1680363874
transform 1 0 128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6434
timestamp 1680363874
transform 1 0 136 0 1 1970
box -8 -3 16 105
use FILL  FILL_6435
timestamp 1680363874
transform 1 0 144 0 1 1970
box -8 -3 16 105
use FILL  FILL_6436
timestamp 1680363874
transform 1 0 152 0 1 1970
box -8 -3 16 105
use FILL  FILL_6437
timestamp 1680363874
transform 1 0 160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6440
timestamp 1680363874
transform 1 0 168 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_65
timestamp 1680363874
transform 1 0 176 0 1 1970
box -8 -3 32 105
use FILL  FILL_6442
timestamp 1680363874
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_6443
timestamp 1680363874
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_6444
timestamp 1680363874
transform 1 0 216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6445
timestamp 1680363874
transform 1 0 224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6446
timestamp 1680363874
transform 1 0 232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6451
timestamp 1680363874
transform 1 0 240 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_66
timestamp 1680363874
transform 1 0 248 0 1 1970
box -8 -3 32 105
use FILL  FILL_6452
timestamp 1680363874
transform 1 0 272 0 1 1970
box -8 -3 16 105
use FILL  FILL_6454
timestamp 1680363874
transform 1 0 280 0 1 1970
box -8 -3 16 105
use FILL  FILL_6456
timestamp 1680363874
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6458
timestamp 1680363874
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6459
timestamp 1680363874
transform 1 0 304 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5245
timestamp 1680363874
transform 1 0 324 0 1 1975
box -3 -3 3 3
use FILL  FILL_6460
timestamp 1680363874
transform 1 0 312 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_403
timestamp 1680363874
transform 1 0 320 0 1 1970
box -9 -3 26 105
use FILL  FILL_6461
timestamp 1680363874
transform 1 0 336 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5246
timestamp 1680363874
transform 1 0 356 0 1 1975
box -3 -3 3 3
use FILL  FILL_6464
timestamp 1680363874
transform 1 0 344 0 1 1970
box -8 -3 16 105
use FAX1  FAX1_16
timestamp 1680363874
transform -1 0 472 0 1 1970
box -5 -3 126 105
use DFFNEGX1  DFFNEGX1_343
timestamp 1680363874
transform 1 0 472 0 1 1970
box -8 -3 104 105
use FAX1  FAX1_17
timestamp 1680363874
transform -1 0 688 0 1 1970
box -5 -3 126 105
use FILL  FILL_6465
timestamp 1680363874
transform 1 0 688 0 1 1970
box -8 -3 16 105
use FILL  FILL_6486
timestamp 1680363874
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_6488
timestamp 1680363874
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FAX1  FAX1_18
timestamp 1680363874
transform -1 0 832 0 1 1970
box -5 -3 126 105
use FILL  FILL_6489
timestamp 1680363874
transform 1 0 832 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_24
timestamp 1680363874
transform -1 0 872 0 1 1970
box -8 -3 40 105
use FILL  FILL_6490
timestamp 1680363874
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6491
timestamp 1680363874
transform 1 0 880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6492
timestamp 1680363874
transform 1 0 888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6493
timestamp 1680363874
transform 1 0 896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6494
timestamp 1680363874
transform 1 0 904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6495
timestamp 1680363874
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6496
timestamp 1680363874
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6497
timestamp 1680363874
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6498
timestamp 1680363874
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6499
timestamp 1680363874
transform 1 0 944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6500
timestamp 1680363874
transform 1 0 952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6501
timestamp 1680363874
transform 1 0 960 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_346
timestamp 1680363874
transform 1 0 968 0 1 1970
box -8 -3 104 105
use FILL  FILL_6502
timestamp 1680363874
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_6503
timestamp 1680363874
transform 1 0 1072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6504
timestamp 1680363874
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_6505
timestamp 1680363874
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5247
timestamp 1680363874
transform 1 0 1108 0 1 1975
box -3 -3 3 3
use FILL  FILL_6506
timestamp 1680363874
transform 1 0 1096 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_273
timestamp 1680363874
transform 1 0 1104 0 1 1970
box -8 -3 46 105
use FILL  FILL_6507
timestamp 1680363874
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_6521
timestamp 1680363874
transform 1 0 1152 0 1 1970
box -8 -3 16 105
use FILL  FILL_6523
timestamp 1680363874
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6525
timestamp 1680363874
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6527
timestamp 1680363874
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6528
timestamp 1680363874
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6529
timestamp 1680363874
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6530
timestamp 1680363874
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_210
timestamp 1680363874
transform -1 0 1248 0 1 1970
box -8 -3 46 105
use FILL  FILL_6531
timestamp 1680363874
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6532
timestamp 1680363874
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6533
timestamp 1680363874
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use FILL  FILL_6534
timestamp 1680363874
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5248
timestamp 1680363874
transform 1 0 1332 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1680363874
transform 1 0 1356 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1680363874
transform 1 0 1380 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_350
timestamp 1680363874
transform -1 0 1376 0 1 1970
box -8 -3 104 105
use FILL  FILL_6535
timestamp 1680363874
transform 1 0 1376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6545
timestamp 1680363874
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5251
timestamp 1680363874
transform 1 0 1444 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1680363874
transform 1 0 1460 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_352
timestamp 1680363874
transform 1 0 1392 0 1 1970
box -8 -3 104 105
use FILL  FILL_6547
timestamp 1680363874
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_6556
timestamp 1680363874
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6558
timestamp 1680363874
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5253
timestamp 1680363874
transform 1 0 1532 0 1 1975
box -3 -3 3 3
use INVX2  INVX2_405
timestamp 1680363874
transform 1 0 1512 0 1 1970
box -9 -3 26 105
use FILL  FILL_6560
timestamp 1680363874
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6561
timestamp 1680363874
transform 1 0 1536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6562
timestamp 1680363874
transform 1 0 1544 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_40
timestamp 1680363874
transform -1 0 1584 0 1 1970
box -8 -3 40 105
use FILL  FILL_6563
timestamp 1680363874
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_6569
timestamp 1680363874
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_6571
timestamp 1680363874
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5254
timestamp 1680363874
transform 1 0 1620 0 1 1975
box -3 -3 3 3
use FILL  FILL_6573
timestamp 1680363874
transform 1 0 1608 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_406
timestamp 1680363874
transform 1 0 1616 0 1 1970
box -9 -3 26 105
use FILL  FILL_6575
timestamp 1680363874
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6576
timestamp 1680363874
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6577
timestamp 1680363874
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_6578
timestamp 1680363874
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_6581
timestamp 1680363874
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_6583
timestamp 1680363874
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use FILL  FILL_6585
timestamp 1680363874
transform 1 0 1680 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_212
timestamp 1680363874
transform 1 0 1688 0 1 1970
box -8 -3 46 105
use FILL  FILL_6587
timestamp 1680363874
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_6588
timestamp 1680363874
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use FILL  FILL_6592
timestamp 1680363874
transform 1 0 1744 0 1 1970
box -8 -3 16 105
use FILL  FILL_6594
timestamp 1680363874
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6596
timestamp 1680363874
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5255
timestamp 1680363874
transform 1 0 1780 0 1 1975
box -3 -3 3 3
use FILL  FILL_6598
timestamp 1680363874
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_6599
timestamp 1680363874
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_6600
timestamp 1680363874
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_213
timestamp 1680363874
transform 1 0 1792 0 1 1970
box -8 -3 46 105
use FILL  FILL_6601
timestamp 1680363874
transform 1 0 1832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6602
timestamp 1680363874
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6603
timestamp 1680363874
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6604
timestamp 1680363874
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5256
timestamp 1680363874
transform 1 0 1884 0 1 1975
box -3 -3 3 3
use INVX2  INVX2_407
timestamp 1680363874
transform -1 0 1880 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_353
timestamp 1680363874
transform 1 0 1880 0 1 1970
box -8 -3 104 105
use FILL  FILL_6605
timestamp 1680363874
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_6606
timestamp 1680363874
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_6607
timestamp 1680363874
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6608
timestamp 1680363874
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_6609
timestamp 1680363874
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1680363874
transform -1 0 2048 0 1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5257
timestamp 1680363874
transform 1 0 2060 0 1 1975
box -3 -3 3 3
use FILL  FILL_6610
timestamp 1680363874
transform 1 0 2048 0 1 1970
box -8 -3 16 105
use FILL  FILL_6626
timestamp 1680363874
transform 1 0 2056 0 1 1970
box -8 -3 16 105
use FILL  FILL_6627
timestamp 1680363874
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_44
timestamp 1680363874
transform 1 0 2072 0 1 1970
box -8 -3 40 105
use FILL  FILL_6628
timestamp 1680363874
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6629
timestamp 1680363874
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_355
timestamp 1680363874
transform 1 0 2120 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_410
timestamp 1680363874
transform 1 0 2216 0 1 1970
box -9 -3 26 105
use FILL  FILL_6630
timestamp 1680363874
transform 1 0 2232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6640
timestamp 1680363874
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6642
timestamp 1680363874
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6643
timestamp 1680363874
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6644
timestamp 1680363874
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use FILL  FILL_6645
timestamp 1680363874
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_45
timestamp 1680363874
transform 1 0 2280 0 1 1970
box -8 -3 40 105
use FILL  FILL_6646
timestamp 1680363874
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6652
timestamp 1680363874
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5258
timestamp 1680363874
transform 1 0 2340 0 1 1975
box -3 -3 3 3
use FILL  FILL_6654
timestamp 1680363874
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_6656
timestamp 1680363874
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use FILL  FILL_6658
timestamp 1680363874
transform 1 0 2344 0 1 1970
box -8 -3 16 105
use FILL  FILL_6659
timestamp 1680363874
transform 1 0 2352 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_47
timestamp 1680363874
transform 1 0 2360 0 1 1970
box -8 -3 40 105
use FILL  FILL_6660
timestamp 1680363874
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6665
timestamp 1680363874
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_6666
timestamp 1680363874
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6667
timestamp 1680363874
transform 1 0 2416 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1680363874
transform -1 0 2456 0 1 1970
box -8 -3 40 105
use FILL  FILL_6668
timestamp 1680363874
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_6669
timestamp 1680363874
transform 1 0 2464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6670
timestamp 1680363874
transform 1 0 2472 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_26
timestamp 1680363874
transform -1 0 2512 0 1 1970
box -8 -3 40 105
use INVX2  INVX2_412
timestamp 1680363874
transform -1 0 2528 0 1 1970
box -9 -3 26 105
use FILL  FILL_6671
timestamp 1680363874
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6672
timestamp 1680363874
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6673
timestamp 1680363874
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_43
timestamp 1680363874
transform 1 0 2552 0 1 1970
box -5 -3 28 105
use NAND3X1  NAND3X1_48
timestamp 1680363874
transform -1 0 2608 0 1 1970
box -8 -3 40 105
use FILL  FILL_6681
timestamp 1680363874
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_6682
timestamp 1680363874
transform 1 0 2616 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_413
timestamp 1680363874
transform 1 0 2624 0 1 1970
box -9 -3 26 105
use FILL  FILL_6683
timestamp 1680363874
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6684
timestamp 1680363874
transform 1 0 2648 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_357
timestamp 1680363874
transform 1 0 2656 0 1 1970
box -8 -3 104 105
use FILL  FILL_6685
timestamp 1680363874
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6686
timestamp 1680363874
transform 1 0 2760 0 1 1970
box -8 -3 16 105
use FILL  FILL_6687
timestamp 1680363874
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_6697
timestamp 1680363874
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_6699
timestamp 1680363874
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_30
timestamp 1680363874
transform 1 0 2792 0 1 1970
box -8 -3 40 105
use FILL  FILL_6700
timestamp 1680363874
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_6703
timestamp 1680363874
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6704
timestamp 1680363874
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_416
timestamp 1680363874
transform 1 0 2848 0 1 1970
box -9 -3 26 105
use FILL  FILL_6705
timestamp 1680363874
transform 1 0 2864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6707
timestamp 1680363874
transform 1 0 2872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6709
timestamp 1680363874
transform 1 0 2880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6711
timestamp 1680363874
transform 1 0 2888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6713
timestamp 1680363874
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_143
timestamp 1680363874
transform 1 0 2904 0 1 1970
box -8 -3 34 105
use FILL  FILL_6714
timestamp 1680363874
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6717
timestamp 1680363874
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6719
timestamp 1680363874
transform 1 0 2952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6720
timestamp 1680363874
transform 1 0 2960 0 1 1970
box -8 -3 16 105
use FILL  FILL_6721
timestamp 1680363874
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use FILL  FILL_6722
timestamp 1680363874
transform 1 0 2976 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_68
timestamp 1680363874
transform -1 0 3008 0 1 1970
box -8 -3 32 105
use FILL  FILL_6723
timestamp 1680363874
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_6724
timestamp 1680363874
transform 1 0 3016 0 1 1970
box -8 -3 16 105
use FILL  FILL_6725
timestamp 1680363874
transform 1 0 3024 0 1 1970
box -8 -3 16 105
use FILL  FILL_6726
timestamp 1680363874
transform 1 0 3032 0 1 1970
box -8 -3 16 105
use FILL  FILL_6727
timestamp 1680363874
transform 1 0 3040 0 1 1970
box -8 -3 16 105
use FILL  FILL_6728
timestamp 1680363874
transform 1 0 3048 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_417
timestamp 1680363874
transform -1 0 3072 0 1 1970
box -9 -3 26 105
use FILL  FILL_6729
timestamp 1680363874
transform 1 0 3072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6730
timestamp 1680363874
transform 1 0 3080 0 1 1970
box -8 -3 16 105
use FILL  FILL_6731
timestamp 1680363874
transform 1 0 3088 0 1 1970
box -8 -3 16 105
use FILL  FILL_6733
timestamp 1680363874
transform 1 0 3096 0 1 1970
box -8 -3 16 105
use FILL  FILL_6735
timestamp 1680363874
transform 1 0 3104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6736
timestamp 1680363874
transform 1 0 3112 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_214
timestamp 1680363874
transform -1 0 3160 0 1 1970
box -8 -3 46 105
use FILL  FILL_6737
timestamp 1680363874
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6738
timestamp 1680363874
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6739
timestamp 1680363874
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6740
timestamp 1680363874
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6741
timestamp 1680363874
transform 1 0 3192 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_215
timestamp 1680363874
transform -1 0 3240 0 1 1970
box -8 -3 46 105
use FILL  FILL_6742
timestamp 1680363874
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6747
timestamp 1680363874
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6749
timestamp 1680363874
transform 1 0 3256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6751
timestamp 1680363874
transform 1 0 3264 0 1 1970
box -8 -3 16 105
use FILL  FILL_6752
timestamp 1680363874
transform 1 0 3272 0 1 1970
box -8 -3 16 105
use FILL  FILL_6753
timestamp 1680363874
transform 1 0 3280 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5259
timestamp 1680363874
transform 1 0 3308 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_216
timestamp 1680363874
transform 1 0 3288 0 1 1970
box -8 -3 46 105
use FILL  FILL_6754
timestamp 1680363874
transform 1 0 3328 0 1 1970
box -8 -3 16 105
use FILL  FILL_6755
timestamp 1680363874
transform 1 0 3336 0 1 1970
box -8 -3 16 105
use FILL  FILL_6758
timestamp 1680363874
transform 1 0 3344 0 1 1970
box -8 -3 16 105
use FILL  FILL_6760
timestamp 1680363874
transform 1 0 3352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6762
timestamp 1680363874
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6764
timestamp 1680363874
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6766
timestamp 1680363874
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6768
timestamp 1680363874
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_217
timestamp 1680363874
transform 1 0 3392 0 1 1970
box -8 -3 46 105
use FILL  FILL_6769
timestamp 1680363874
transform 1 0 3432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6772
timestamp 1680363874
transform 1 0 3440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6774
timestamp 1680363874
transform 1 0 3448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6776
timestamp 1680363874
transform 1 0 3456 0 1 1970
box -8 -3 16 105
use FILL  FILL_6778
timestamp 1680363874
transform 1 0 3464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6780
timestamp 1680363874
transform 1 0 3472 0 1 1970
box -8 -3 16 105
use FILL  FILL_6782
timestamp 1680363874
transform 1 0 3480 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_69
timestamp 1680363874
transform 1 0 3488 0 1 1970
box -8 -3 32 105
use FILL  FILL_6784
timestamp 1680363874
transform 1 0 3512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6785
timestamp 1680363874
transform 1 0 3520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6786
timestamp 1680363874
transform 1 0 3528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6787
timestamp 1680363874
transform 1 0 3536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6790
timestamp 1680363874
transform 1 0 3544 0 1 1970
box -8 -3 16 105
use FILL  FILL_6792
timestamp 1680363874
transform 1 0 3552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6794
timestamp 1680363874
transform 1 0 3560 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_420
timestamp 1680363874
transform 1 0 3568 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_5260
timestamp 1680363874
transform 1 0 3652 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_361
timestamp 1680363874
transform 1 0 3584 0 1 1970
box -8 -3 104 105
use FILL  FILL_6796
timestamp 1680363874
transform 1 0 3680 0 1 1970
box -8 -3 16 105
use FILL  FILL_6797
timestamp 1680363874
transform 1 0 3688 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5261
timestamp 1680363874
transform 1 0 3708 0 1 1975
box -3 -3 3 3
use FILL  FILL_6798
timestamp 1680363874
transform 1 0 3696 0 1 1970
box -8 -3 16 105
use FILL  FILL_6799
timestamp 1680363874
transform 1 0 3704 0 1 1970
box -8 -3 16 105
use FILL  FILL_6810
timestamp 1680363874
transform 1 0 3712 0 1 1970
box -8 -3 16 105
use FILL  FILL_6812
timestamp 1680363874
transform 1 0 3720 0 1 1970
box -8 -3 16 105
use FILL  FILL_6814
timestamp 1680363874
transform 1 0 3728 0 1 1970
box -8 -3 16 105
use FILL  FILL_6816
timestamp 1680363874
transform 1 0 3736 0 1 1970
box -8 -3 16 105
use FILL  FILL_6818
timestamp 1680363874
transform 1 0 3744 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_219
timestamp 1680363874
transform -1 0 3792 0 1 1970
box -8 -3 46 105
use FILL  FILL_6819
timestamp 1680363874
transform 1 0 3792 0 1 1970
box -8 -3 16 105
use FILL  FILL_6824
timestamp 1680363874
transform 1 0 3800 0 1 1970
box -8 -3 16 105
use FILL  FILL_6826
timestamp 1680363874
transform 1 0 3808 0 1 1970
box -8 -3 16 105
use FILL  FILL_6828
timestamp 1680363874
transform 1 0 3816 0 1 1970
box -8 -3 16 105
use FILL  FILL_6830
timestamp 1680363874
transform 1 0 3824 0 1 1970
box -8 -3 16 105
use FILL  FILL_6831
timestamp 1680363874
transform 1 0 3832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6832
timestamp 1680363874
transform 1 0 3840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6833
timestamp 1680363874
transform 1 0 3848 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_280
timestamp 1680363874
transform 1 0 3856 0 1 1970
box -8 -3 46 105
use FILL  FILL_6835
timestamp 1680363874
transform 1 0 3896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6836
timestamp 1680363874
transform 1 0 3904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6841
timestamp 1680363874
transform 1 0 3912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6842
timestamp 1680363874
transform 1 0 3920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6843
timestamp 1680363874
transform 1 0 3928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6844
timestamp 1680363874
transform 1 0 3936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6846
timestamp 1680363874
transform 1 0 3944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6848
timestamp 1680363874
transform 1 0 3952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6850
timestamp 1680363874
transform 1 0 3960 0 1 1970
box -8 -3 16 105
use FILL  FILL_6852
timestamp 1680363874
transform 1 0 3968 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_47
timestamp 1680363874
transform -1 0 4000 0 1 1970
box -5 -3 28 105
use FILL  FILL_6853
timestamp 1680363874
transform 1 0 4000 0 1 1970
box -8 -3 16 105
use FILL  FILL_6856
timestamp 1680363874
transform 1 0 4008 0 1 1970
box -8 -3 16 105
use FILL  FILL_6858
timestamp 1680363874
transform 1 0 4016 0 1 1970
box -8 -3 16 105
use FILL  FILL_6859
timestamp 1680363874
transform 1 0 4024 0 1 1970
box -8 -3 16 105
use FILL  FILL_6860
timestamp 1680363874
transform 1 0 4032 0 1 1970
box -8 -3 16 105
use FILL  FILL_6861
timestamp 1680363874
transform 1 0 4040 0 1 1970
box -8 -3 16 105
use FILL  FILL_6862
timestamp 1680363874
transform 1 0 4048 0 1 1970
box -8 -3 16 105
use FILL  FILL_6863
timestamp 1680363874
transform 1 0 4056 0 1 1970
box -8 -3 16 105
use FILL  FILL_6864
timestamp 1680363874
transform 1 0 4064 0 1 1970
box -8 -3 16 105
use FILL  FILL_6867
timestamp 1680363874
transform 1 0 4072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6869
timestamp 1680363874
transform 1 0 4080 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_220
timestamp 1680363874
transform -1 0 4128 0 1 1970
box -8 -3 46 105
use FILL  FILL_6870
timestamp 1680363874
transform 1 0 4128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6878
timestamp 1680363874
transform 1 0 4136 0 1 1970
box -8 -3 16 105
use FILL  FILL_6879
timestamp 1680363874
transform 1 0 4144 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_421
timestamp 1680363874
transform -1 0 4168 0 1 1970
box -9 -3 26 105
use FILL  FILL_6880
timestamp 1680363874
transform 1 0 4168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6883
timestamp 1680363874
transform 1 0 4176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6885
timestamp 1680363874
transform 1 0 4184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6887
timestamp 1680363874
transform 1 0 4192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6889
timestamp 1680363874
transform 1 0 4200 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_49
timestamp 1680363874
transform -1 0 4232 0 1 1970
box -5 -3 28 105
use FILL  FILL_6890
timestamp 1680363874
transform 1 0 4232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6891
timestamp 1680363874
transform 1 0 4240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6892
timestamp 1680363874
transform 1 0 4248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6893
timestamp 1680363874
transform 1 0 4256 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_422
timestamp 1680363874
transform -1 0 4280 0 1 1970
box -9 -3 26 105
use FILL  FILL_6894
timestamp 1680363874
transform 1 0 4280 0 1 1970
box -8 -3 16 105
use FILL  FILL_6901
timestamp 1680363874
transform 1 0 4288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6903
timestamp 1680363874
transform 1 0 4296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6905
timestamp 1680363874
transform 1 0 4304 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_221
timestamp 1680363874
transform -1 0 4352 0 1 1970
box -8 -3 46 105
use FILL  FILL_6906
timestamp 1680363874
transform 1 0 4352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6911
timestamp 1680363874
transform 1 0 4360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6913
timestamp 1680363874
transform 1 0 4368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6915
timestamp 1680363874
transform 1 0 4376 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_51
timestamp 1680363874
transform 1 0 4384 0 1 1970
box -5 -3 28 105
use FILL  FILL_6916
timestamp 1680363874
transform 1 0 4408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6919
timestamp 1680363874
transform 1 0 4416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6921
timestamp 1680363874
transform 1 0 4424 0 1 1970
box -8 -3 16 105
use FILL  FILL_6923
timestamp 1680363874
transform 1 0 4432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6924
timestamp 1680363874
transform 1 0 4440 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_222
timestamp 1680363874
transform 1 0 4448 0 1 1970
box -8 -3 46 105
use FILL  FILL_6925
timestamp 1680363874
transform 1 0 4488 0 1 1970
box -8 -3 16 105
use FILL  FILL_6929
timestamp 1680363874
transform 1 0 4496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6931
timestamp 1680363874
transform 1 0 4504 0 1 1970
box -8 -3 16 105
use FILL  FILL_6933
timestamp 1680363874
transform 1 0 4512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6935
timestamp 1680363874
transform 1 0 4520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6937
timestamp 1680363874
transform 1 0 4528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6938
timestamp 1680363874
transform 1 0 4536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6939
timestamp 1680363874
transform 1 0 4544 0 1 1970
box -8 -3 16 105
use FILL  FILL_6940
timestamp 1680363874
transform 1 0 4552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6942
timestamp 1680363874
transform 1 0 4560 0 1 1970
box -8 -3 16 105
use FILL  FILL_6943
timestamp 1680363874
transform 1 0 4568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6944
timestamp 1680363874
transform 1 0 4576 0 1 1970
box -8 -3 16 105
use FILL  FILL_6945
timestamp 1680363874
transform 1 0 4584 0 1 1970
box -8 -3 16 105
use FILL  FILL_6946
timestamp 1680363874
transform 1 0 4592 0 1 1970
box -8 -3 16 105
use FILL  FILL_6947
timestamp 1680363874
transform 1 0 4600 0 1 1970
box -8 -3 16 105
use FILL  FILL_6948
timestamp 1680363874
transform 1 0 4608 0 1 1970
box -8 -3 16 105
use FILL  FILL_6951
timestamp 1680363874
transform 1 0 4616 0 1 1970
box -8 -3 16 105
use FILL  FILL_6953
timestamp 1680363874
transform 1 0 4624 0 1 1970
box -8 -3 16 105
use FILL  FILL_6955
timestamp 1680363874
transform 1 0 4632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6957
timestamp 1680363874
transform 1 0 4640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6958
timestamp 1680363874
transform 1 0 4648 0 1 1970
box -8 -3 16 105
use FILL  FILL_6959
timestamp 1680363874
transform 1 0 4656 0 1 1970
box -8 -3 16 105
use FILL  FILL_6960
timestamp 1680363874
transform 1 0 4664 0 1 1970
box -8 -3 16 105
use FILL  FILL_6961
timestamp 1680363874
transform 1 0 4672 0 1 1970
box -8 -3 16 105
use FILL  FILL_6962
timestamp 1680363874
transform 1 0 4680 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_423
timestamp 1680363874
transform 1 0 4688 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_362
timestamp 1680363874
transform 1 0 4704 0 1 1970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_55
timestamp 1680363874
transform 1 0 4827 0 1 1970
box -10 -3 10 3
use M3_M2  M3_M2_5273
timestamp 1680363874
transform 1 0 100 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5828
timestamp 1680363874
transform 1 0 124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1680363874
transform 1 0 92 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5274
timestamp 1680363874
transform 1 0 156 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5829
timestamp 1680363874
transform 1 0 156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1680363874
transform 1 0 164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1680363874
transform 1 0 148 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5328
timestamp 1680363874
transform 1 0 172 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1680363874
transform 1 0 220 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5910
timestamp 1680363874
transform 1 0 212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1680363874
transform 1 0 220 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5314
timestamp 1680363874
transform 1 0 236 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5831
timestamp 1680363874
transform 1 0 236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1680363874
transform 1 0 236 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5275
timestamp 1680363874
transform 1 0 252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1680363874
transform 1 0 276 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5832
timestamp 1680363874
transform 1 0 276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1680363874
transform 1 0 252 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5351
timestamp 1680363874
transform 1 0 268 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_6016
timestamp 1680363874
transform 1 0 260 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1680363874
transform 1 0 284 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1680363874
transform 1 0 300 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5316
timestamp 1680363874
transform 1 0 332 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5833
timestamp 1680363874
transform 1 0 332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1680363874
transform 1 0 324 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5352
timestamp 1680363874
transform 1 0 332 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5914
timestamp 1680363874
transform 1 0 348 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5276
timestamp 1680363874
transform 1 0 404 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1680363874
transform 1 0 532 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1680363874
transform 1 0 564 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1680363874
transform 1 0 556 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5834
timestamp 1680363874
transform 1 0 548 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1680363874
transform 1 0 524 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5353
timestamp 1680363874
transform 1 0 548 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1680363874
transform 1 0 652 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1680363874
transform 1 0 676 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5835
timestamp 1680363874
transform 1 0 676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1680363874
transform 1 0 596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1680363874
transform 1 0 652 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5354
timestamp 1680363874
transform 1 0 676 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1680363874
transform 1 0 636 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1680363874
transform 1 0 692 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5918
timestamp 1680363874
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5378
timestamp 1680363874
transform 1 0 692 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1680363874
transform 1 0 700 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1680363874
transform 1 0 748 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5836
timestamp 1680363874
transform 1 0 796 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5355
timestamp 1680363874
transform 1 0 764 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5919
timestamp 1680363874
transform 1 0 772 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5356
timestamp 1680363874
transform 1 0 796 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1680363874
transform 1 0 876 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1680363874
transform 1 0 876 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5837
timestamp 1680363874
transform 1 0 892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1680363874
transform 1 0 812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1680363874
transform 1 0 844 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5357
timestamp 1680363874
transform 1 0 892 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1680363874
transform 1 0 964 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5838
timestamp 1680363874
transform 1 0 988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1680363874
transform 1 0 1004 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1680363874
transform 1 0 908 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5379
timestamp 1680363874
transform 1 0 828 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1680363874
transform 1 0 916 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5923
timestamp 1680363874
transform 1 0 964 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5359
timestamp 1680363874
transform 1 0 1004 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1680363874
transform 1 0 916 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5840
timestamp 1680363874
transform 1 0 1020 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5282
timestamp 1680363874
transform 1 0 1036 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1680363874
transform 1 0 1076 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1680363874
transform 1 0 1076 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5841
timestamp 1680363874
transform 1 0 1084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1680363874
transform 1 0 1068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1680363874
transform 1 0 1076 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5360
timestamp 1680363874
transform 1 0 1084 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5926
timestamp 1680363874
transform 1 0 1092 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5381
timestamp 1680363874
transform 1 0 1068 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1680363874
transform 1 0 1092 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1680363874
transform 1 0 1116 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5842
timestamp 1680363874
transform 1 0 1140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1680363874
transform 1 0 1148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1680363874
transform 1 0 1132 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5383
timestamp 1680363874
transform 1 0 1148 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1680363874
transform 1 0 1204 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5820
timestamp 1680363874
transform 1 0 1228 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1680363874
transform 1 0 1188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1680363874
transform 1 0 1204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1680363874
transform 1 0 1220 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5384
timestamp 1680363874
transform 1 0 1204 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1680363874
transform 1 0 1220 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1680363874
transform 1 0 1188 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5821
timestamp 1680363874
transform 1 0 1252 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1680363874
transform 1 0 1252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1680363874
transform 1 0 1244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1680363874
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5284
timestamp 1680363874
transform 1 0 1308 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1680363874
transform 1 0 1324 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1680363874
transform 1 0 1340 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5845
timestamp 1680363874
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1680363874
transform 1 0 1292 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5406
timestamp 1680363874
transform 1 0 1260 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1680363874
transform 1 0 1292 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5846
timestamp 1680363874
transform 1 0 1356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1680363874
transform 1 0 1356 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5386
timestamp 1680363874
transform 1 0 1356 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1680363874
transform 1 0 1404 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5847
timestamp 1680363874
transform 1 0 1428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1680363874
transform 1 0 1444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1680363874
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5362
timestamp 1680363874
transform 1 0 1444 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5936
timestamp 1680363874
transform 1 0 1452 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5387
timestamp 1680363874
transform 1 0 1452 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5849
timestamp 1680363874
transform 1 0 1508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1680363874
transform 1 0 1516 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5265
timestamp 1680363874
transform 1 0 1564 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5850
timestamp 1680363874
transform 1 0 1540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1680363874
transform 1 0 1556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1680363874
transform 1 0 1548 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5363
timestamp 1680363874
transform 1 0 1556 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_6010
timestamp 1680363874
transform 1 0 1564 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5266
timestamp 1680363874
transform 1 0 1652 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5939
timestamp 1680363874
transform 1 0 1644 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5408
timestamp 1680363874
transform 1 0 1644 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_6017
timestamp 1680363874
transform 1 0 1660 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5420
timestamp 1680363874
transform 1 0 1668 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_6011
timestamp 1680363874
transform 1 0 1692 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1680363874
transform 1 0 1700 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1680363874
transform 1 0 1716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1680363874
transform 1 0 1732 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1680363874
transform 1 0 1724 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5409
timestamp 1680363874
transform 1 0 1732 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1680363874
transform 1 0 1732 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1680363874
transform 1 0 1756 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1680363874
transform 1 0 1780 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5852
timestamp 1680363874
transform 1 0 1780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1680363874
transform 1 0 1820 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5364
timestamp 1680363874
transform 1 0 1852 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1680363874
transform 1 0 1820 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1680363874
transform 1 0 1852 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1680363874
transform 1 0 1892 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5942
timestamp 1680363874
transform 1 0 1892 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5334
timestamp 1680363874
transform 1 0 1908 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1680363874
transform 1 0 1940 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5853
timestamp 1680363874
transform 1 0 1940 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5365
timestamp 1680363874
transform 1 0 1940 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5854
timestamp 1680363874
transform 1 0 1956 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5291
timestamp 1680363874
transform 1 0 1972 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5943
timestamp 1680363874
transform 1 0 1964 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5317
timestamp 1680363874
transform 1 0 1980 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5855
timestamp 1680363874
transform 1 0 1988 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5335
timestamp 1680363874
transform 1 0 1996 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5944
timestamp 1680363874
transform 1 0 1980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1680363874
transform 1 0 1996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1680363874
transform 1 0 2012 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5366
timestamp 1680363874
transform 1 0 2012 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5857
timestamp 1680363874
transform 1 0 2068 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5336
timestamp 1680363874
transform 1 0 2092 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1680363874
transform 1 0 2116 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5946
timestamp 1680363874
transform 1 0 2116 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5423
timestamp 1680363874
transform 1 0 2060 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1680363874
transform 1 0 2156 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5947
timestamp 1680363874
transform 1 0 2188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1680363874
transform 1 0 2204 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1680363874
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1680363874
transform 1 0 2300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1680363874
transform 1 0 2348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1680363874
transform 1 0 2340 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1680363874
transform 1 0 2372 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5318
timestamp 1680363874
transform 1 0 2404 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5858
timestamp 1680363874
transform 1 0 2404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1680363874
transform 1 0 2428 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5390
timestamp 1680363874
transform 1 0 2428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1680363874
transform 1 0 2444 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5952
timestamp 1680363874
transform 1 0 2452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1680363874
transform 1 0 2468 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5293
timestamp 1680363874
transform 1 0 2484 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1680363874
transform 1 0 2500 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1680363874
transform 1 0 2492 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1680363874
transform 1 0 2540 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1680363874
transform 1 0 2532 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5859
timestamp 1680363874
transform 1 0 2508 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5338
timestamp 1680363874
transform 1 0 2516 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5860
timestamp 1680363874
transform 1 0 2540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1680363874
transform 1 0 2516 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1680363874
transform 1 0 2532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1680363874
transform 1 0 2548 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5392
timestamp 1680363874
transform 1 0 2540 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1680363874
transform 1 0 2532 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1680363874
transform 1 0 2564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1680363874
transform 1 0 2580 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1680363874
transform 1 0 2596 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5861
timestamp 1680363874
transform 1 0 2604 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5368
timestamp 1680363874
transform 1 0 2604 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1680363874
transform 1 0 2620 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1680363874
transform 1 0 2668 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5862
timestamp 1680363874
transform 1 0 2620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1680363874
transform 1 0 2652 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5393
timestamp 1680363874
transform 1 0 2644 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1680363874
transform 1 0 2628 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5958
timestamp 1680363874
transform 1 0 2716 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5394
timestamp 1680363874
transform 1 0 2716 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5863
timestamp 1680363874
transform 1 0 2756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1680363874
transform 1 0 2764 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5426
timestamp 1680363874
transform 1 0 2756 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1680363874
transform 1 0 2828 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5865
timestamp 1680363874
transform 1 0 2820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1680363874
transform 1 0 2796 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5369
timestamp 1680363874
transform 1 0 2812 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1680363874
transform 1 0 2796 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5960
timestamp 1680363874
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5267
timestamp 1680363874
transform 1 0 2860 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5961
timestamp 1680363874
transform 1 0 2844 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5427
timestamp 1680363874
transform 1 0 2844 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1680363874
transform 1 0 2868 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5866
timestamp 1680363874
transform 1 0 2868 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5370
timestamp 1680363874
transform 1 0 2876 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1680363874
transform 1 0 2892 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5962
timestamp 1680363874
transform 1 0 2892 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5428
timestamp 1680363874
transform 1 0 2892 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5963
timestamp 1680363874
transform 1 0 2908 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5429
timestamp 1680363874
transform 1 0 2916 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1680363874
transform 1 0 2948 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5964
timestamp 1680363874
transform 1 0 2940 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5410
timestamp 1680363874
transform 1 0 2940 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_6020
timestamp 1680363874
transform 1 0 2948 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1680363874
transform 1 0 2972 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5340
timestamp 1680363874
transform 1 0 2980 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5868
timestamp 1680363874
transform 1 0 3060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1680363874
transform 1 0 2980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1680363874
transform 1 0 3036 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5371
timestamp 1680363874
transform 1 0 3060 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5967
timestamp 1680363874
transform 1 0 3076 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5396
timestamp 1680363874
transform 1 0 2972 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1680363874
transform 1 0 2996 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1680363874
transform 1 0 3036 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1680363874
transform 1 0 3076 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1680363874
transform 1 0 3004 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1680363874
transform 1 0 3020 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1680363874
transform 1 0 3100 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5869
timestamp 1680363874
transform 1 0 3100 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5400
timestamp 1680363874
transform 1 0 3100 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1680363874
transform 1 0 3100 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1680363874
transform 1 0 3124 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1680363874
transform 1 0 3140 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5870
timestamp 1680363874
transform 1 0 3116 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5341
timestamp 1680363874
transform 1 0 3164 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1680363874
transform 1 0 3116 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1680363874
transform 1 0 3140 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1680363874
transform 1 0 3204 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5968
timestamp 1680363874
transform 1 0 3164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1680363874
transform 1 0 3196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1680363874
transform 1 0 3204 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5437
timestamp 1680363874
transform 1 0 3156 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5871
timestamp 1680363874
transform 1 0 3220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1680363874
transform 1 0 3228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1680363874
transform 1 0 3260 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5270
timestamp 1680363874
transform 1 0 3300 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5874
timestamp 1680363874
transform 1 0 3300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1680363874
transform 1 0 3276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1680363874
transform 1 0 3292 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5411
timestamp 1680363874
transform 1 0 3284 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1680363874
transform 1 0 3292 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5973
timestamp 1680363874
transform 1 0 3316 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5320
timestamp 1680363874
transform 1 0 3356 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5974
timestamp 1680363874
transform 1 0 3356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1680363874
transform 1 0 3364 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5304
timestamp 1680363874
transform 1 0 3404 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5875
timestamp 1680363874
transform 1 0 3388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1680363874
transform 1 0 3404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1680363874
transform 1 0 3412 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5412
timestamp 1680363874
transform 1 0 3412 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5977
timestamp 1680363874
transform 1 0 3452 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5413
timestamp 1680363874
transform 1 0 3444 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5877
timestamp 1680363874
transform 1 0 3492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1680363874
transform 1 0 3500 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1680363874
transform 1 0 3516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1680363874
transform 1 0 3524 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5414
timestamp 1680363874
transform 1 0 3524 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1680363874
transform 1 0 3516 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1680363874
transform 1 0 3548 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5979
timestamp 1680363874
transform 1 0 3556 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5401
timestamp 1680363874
transform 1 0 3556 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1680363874
transform 1 0 3604 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1680363874
transform 1 0 3628 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1680363874
transform 1 0 3612 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5880
timestamp 1680363874
transform 1 0 3604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1680363874
transform 1 0 3612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1680363874
transform 1 0 3604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1680363874
transform 1 0 3620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1680363874
transform 1 0 3636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1680363874
transform 1 0 3644 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5305
timestamp 1680363874
transform 1 0 3684 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5882
timestamp 1680363874
transform 1 0 3676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1680363874
transform 1 0 3684 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5374
timestamp 1680363874
transform 1 0 3716 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1680363874
transform 1 0 3732 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5822
timestamp 1680363874
transform 1 0 3732 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1680363874
transform 1 0 3748 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1680363874
transform 1 0 3764 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5415
timestamp 1680363874
transform 1 0 3756 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5984
timestamp 1680363874
transform 1 0 3820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1680363874
transform 1 0 3828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1680363874
transform 1 0 3844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1680363874
transform 1 0 3852 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5307
timestamp 1680363874
transform 1 0 3876 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5986
timestamp 1680363874
transform 1 0 3884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1680363874
transform 1 0 3908 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5343
timestamp 1680363874
transform 1 0 3908 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5987
timestamp 1680363874
transform 1 0 3908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1680363874
transform 1 0 3932 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5344
timestamp 1680363874
transform 1 0 3940 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5988
timestamp 1680363874
transform 1 0 3940 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1680363874
transform 1 0 3996 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5375
timestamp 1680363874
transform 1 0 3988 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5889
timestamp 1680363874
transform 1 0 4028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1680363874
transform 1 0 4044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1680363874
transform 1 0 4036 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5376
timestamp 1680363874
transform 1 0 4044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1680363874
transform 1 0 4028 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5891
timestamp 1680363874
transform 1 0 4068 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5439
timestamp 1680363874
transform 1 0 4116 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1680363874
transform 1 0 4140 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5825
timestamp 1680363874
transform 1 0 4140 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5345
timestamp 1680363874
transform 1 0 4140 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5990
timestamp 1680363874
transform 1 0 4140 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5346
timestamp 1680363874
transform 1 0 4180 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5892
timestamp 1680363874
transform 1 0 4188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1680363874
transform 1 0 4172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1680363874
transform 1 0 4196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1680363874
transform 1 0 4220 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5309
timestamp 1680363874
transform 1 0 4252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1680363874
transform 1 0 4260 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5894
timestamp 1680363874
transform 1 0 4252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1680363874
transform 1 0 4260 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5402
timestamp 1680363874
transform 1 0 4260 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5994
timestamp 1680363874
transform 1 0 4276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1680363874
transform 1 0 4300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1680363874
transform 1 0 4332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1680363874
transform 1 0 4356 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5310
timestamp 1680363874
transform 1 0 4380 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5826
timestamp 1680363874
transform 1 0 4380 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5347
timestamp 1680363874
transform 1 0 4380 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5898
timestamp 1680363874
transform 1 0 4420 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5348
timestamp 1680363874
transform 1 0 4436 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5995
timestamp 1680363874
transform 1 0 4436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5311
timestamp 1680363874
transform 1 0 4460 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5899
timestamp 1680363874
transform 1 0 4460 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5349
timestamp 1680363874
transform 1 0 4468 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5996
timestamp 1680363874
transform 1 0 4452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1680363874
transform 1 0 4468 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5403
timestamp 1680363874
transform 1 0 4452 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5900
timestamp 1680363874
transform 1 0 4484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1680363874
transform 1 0 4500 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5312
timestamp 1680363874
transform 1 0 4532 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1680363874
transform 1 0 4524 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5827
timestamp 1680363874
transform 1 0 4532 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1680363874
transform 1 0 4556 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5313
timestamp 1680363874
transform 1 0 4588 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5902
timestamp 1680363874
transform 1 0 4572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1680363874
transform 1 0 4588 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5350
timestamp 1680363874
transform 1 0 4604 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5999
timestamp 1680363874
transform 1 0 4580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1680363874
transform 1 0 4604 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5404
timestamp 1680363874
transform 1 0 4572 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1680363874
transform 1 0 4580 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1680363874
transform 1 0 4644 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1680363874
transform 1 0 4676 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5904
timestamp 1680363874
transform 1 0 4644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1680363874
transform 1 0 4652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1680363874
transform 1 0 4676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1680363874
transform 1 0 4636 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5417
timestamp 1680363874
transform 1 0 4628 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_6002
timestamp 1680363874
transform 1 0 4660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1680363874
transform 1 0 4676 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5405
timestamp 1680363874
transform 1 0 4660 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1680363874
transform 1 0 4676 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_6004
timestamp 1680363874
transform 1 0 4692 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5327
timestamp 1680363874
transform 1 0 4796 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5907
timestamp 1680363874
transform 1 0 4716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1680363874
transform 1 0 4756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1680363874
transform 1 0 4796 0 1 1925
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_56
timestamp 1680363874
transform 1 0 24 0 1 1870
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1680363874
transform -1 0 128 0 -1 1970
box -8 -3 64 105
use FILL  FILL_6438
timestamp 1680363874
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1680363874
transform -1 0 160 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6439
timestamp 1680363874
transform 1 0 160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6441
timestamp 1680363874
transform 1 0 168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6447
timestamp 1680363874
transform 1 0 176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6448
timestamp 1680363874
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6449
timestamp 1680363874
transform 1 0 192 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_401
timestamp 1680363874
transform 1 0 200 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_402
timestamp 1680363874
transform -1 0 232 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6450
timestamp 1680363874
transform 1 0 232 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_39
timestamp 1680363874
transform 1 0 240 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6453
timestamp 1680363874
transform 1 0 272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6455
timestamp 1680363874
transform 1 0 280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6457
timestamp 1680363874
transform 1 0 288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6462
timestamp 1680363874
transform 1 0 296 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_142
timestamp 1680363874
transform -1 0 336 0 -1 1970
box -8 -3 34 105
use FILL  FILL_6463
timestamp 1680363874
transform 1 0 336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6466
timestamp 1680363874
transform 1 0 344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6467
timestamp 1680363874
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6468
timestamp 1680363874
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6469
timestamp 1680363874
transform 1 0 368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6470
timestamp 1680363874
transform 1 0 376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6471
timestamp 1680363874
transform 1 0 384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6472
timestamp 1680363874
transform 1 0 392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6473
timestamp 1680363874
transform 1 0 400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6474
timestamp 1680363874
transform 1 0 408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6475
timestamp 1680363874
transform 1 0 416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6476
timestamp 1680363874
transform 1 0 424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6477
timestamp 1680363874
transform 1 0 432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6478
timestamp 1680363874
transform 1 0 440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6479
timestamp 1680363874
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6480
timestamp 1680363874
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_344
timestamp 1680363874
transform -1 0 560 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6481
timestamp 1680363874
transform 1 0 560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6482
timestamp 1680363874
transform 1 0 568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6483
timestamp 1680363874
transform 1 0 576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6484
timestamp 1680363874
transform 1 0 584 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_345
timestamp 1680363874
transform -1 0 688 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6485
timestamp 1680363874
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6487
timestamp 1680363874
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6508
timestamp 1680363874
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_347
timestamp 1680363874
transform -1 0 808 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_348
timestamp 1680363874
transform -1 0 904 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_349
timestamp 1680363874
transform -1 0 1000 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_404
timestamp 1680363874
transform 1 0 1000 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6509
timestamp 1680363874
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6510
timestamp 1680363874
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6511
timestamp 1680363874
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6512
timestamp 1680363874
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6513
timestamp 1680363874
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6514
timestamp 1680363874
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_274
timestamp 1680363874
transform 1 0 1064 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6515
timestamp 1680363874
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6516
timestamp 1680363874
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6517
timestamp 1680363874
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6518
timestamp 1680363874
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6519
timestamp 1680363874
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6520
timestamp 1680363874
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6522
timestamp 1680363874
transform 1 0 1152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6524
timestamp 1680363874
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6526
timestamp 1680363874
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6536
timestamp 1680363874
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_211
timestamp 1680363874
transform -1 0 1224 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6537
timestamp 1680363874
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5440
timestamp 1680363874
transform 1 0 1244 0 1 1875
box -3 -3 3 3
use FILL  FILL_6538
timestamp 1680363874
transform 1 0 1232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6539
timestamp 1680363874
transform 1 0 1240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6540
timestamp 1680363874
transform 1 0 1248 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_351
timestamp 1680363874
transform -1 0 1352 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6541
timestamp 1680363874
transform 1 0 1352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6542
timestamp 1680363874
transform 1 0 1360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6543
timestamp 1680363874
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6544
timestamp 1680363874
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6546
timestamp 1680363874
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6548
timestamp 1680363874
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6549
timestamp 1680363874
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_275
timestamp 1680363874
transform 1 0 1408 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6550
timestamp 1680363874
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6551
timestamp 1680363874
transform 1 0 1456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6552
timestamp 1680363874
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5441
timestamp 1680363874
transform 1 0 1484 0 1 1875
box -3 -3 3 3
use FILL  FILL_6553
timestamp 1680363874
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6554
timestamp 1680363874
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6555
timestamp 1680363874
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6557
timestamp 1680363874
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6559
timestamp 1680363874
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6564
timestamp 1680363874
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5442
timestamp 1680363874
transform 1 0 1548 0 1 1875
box -3 -3 3 3
use OAI22X1  OAI22X1_276
timestamp 1680363874
transform 1 0 1520 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6565
timestamp 1680363874
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6566
timestamp 1680363874
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6567
timestamp 1680363874
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6568
timestamp 1680363874
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6570
timestamp 1680363874
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6572
timestamp 1680363874
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6574
timestamp 1680363874
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6579
timestamp 1680363874
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5443
timestamp 1680363874
transform 1 0 1660 0 1 1875
box -3 -3 3 3
use NAND3X1  NAND3X1_41
timestamp 1680363874
transform -1 0 1656 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6580
timestamp 1680363874
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6582
timestamp 1680363874
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6584
timestamp 1680363874
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6586
timestamp 1680363874
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6589
timestamp 1680363874
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6590
timestamp 1680363874
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_42
timestamp 1680363874
transform 1 0 1704 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6591
timestamp 1680363874
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5444
timestamp 1680363874
transform 1 0 1756 0 1 1875
box -3 -3 3 3
use FILL  FILL_6593
timestamp 1680363874
transform 1 0 1744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6595
timestamp 1680363874
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6597
timestamp 1680363874
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5445
timestamp 1680363874
transform 1 0 1860 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_354
timestamp 1680363874
transform 1 0 1768 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6611
timestamp 1680363874
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6612
timestamp 1680363874
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_408
timestamp 1680363874
transform 1 0 1880 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6613
timestamp 1680363874
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6614
timestamp 1680363874
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6615
timestamp 1680363874
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6616
timestamp 1680363874
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6617
timestamp 1680363874
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_409
timestamp 1680363874
transform 1 0 1936 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6618
timestamp 1680363874
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6619
timestamp 1680363874
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5446
timestamp 1680363874
transform 1 0 1980 0 1 1875
box -3 -3 3 3
use OAI22X1  OAI22X1_277
timestamp 1680363874
transform -1 0 2008 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6620
timestamp 1680363874
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6621
timestamp 1680363874
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5447
timestamp 1680363874
transform 1 0 2036 0 1 1875
box -3 -3 3 3
use FILL  FILL_6622
timestamp 1680363874
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6623
timestamp 1680363874
transform 1 0 2032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6624
timestamp 1680363874
transform 1 0 2040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6625
timestamp 1680363874
transform 1 0 2048 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_356
timestamp 1680363874
transform 1 0 2056 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5448
timestamp 1680363874
transform 1 0 2164 0 1 1875
box -3 -3 3 3
use FILL  FILL_6631
timestamp 1680363874
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6632
timestamp 1680363874
transform 1 0 2160 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_411
timestamp 1680363874
transform 1 0 2168 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6633
timestamp 1680363874
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6634
timestamp 1680363874
transform 1 0 2192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6635
timestamp 1680363874
transform 1 0 2200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6636
timestamp 1680363874
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6637
timestamp 1680363874
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6638
timestamp 1680363874
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5449
timestamp 1680363874
transform 1 0 2244 0 1 1875
box -3 -3 3 3
use FILL  FILL_6639
timestamp 1680363874
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6641
timestamp 1680363874
transform 1 0 2240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6647
timestamp 1680363874
transform 1 0 2248 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_46
timestamp 1680363874
transform -1 0 2288 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6648
timestamp 1680363874
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6649
timestamp 1680363874
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6650
timestamp 1680363874
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6651
timestamp 1680363874
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5450
timestamp 1680363874
transform 1 0 2332 0 1 1875
box -3 -3 3 3
use FILL  FILL_6653
timestamp 1680363874
transform 1 0 2320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6655
timestamp 1680363874
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6657
timestamp 1680363874
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5451
timestamp 1680363874
transform 1 0 2364 0 1 1875
box -3 -3 3 3
use BUFX2  BUFX2_42
timestamp 1680363874
transform 1 0 2344 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6661
timestamp 1680363874
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6662
timestamp 1680363874
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6663
timestamp 1680363874
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6664
timestamp 1680363874
transform 1 0 2392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6674
timestamp 1680363874
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_27
timestamp 1680363874
transform -1 0 2440 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6675
timestamp 1680363874
transform 1 0 2440 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_28
timestamp 1680363874
transform -1 0 2480 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6676
timestamp 1680363874
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6677
timestamp 1680363874
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6678
timestamp 1680363874
transform 1 0 2496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6679
timestamp 1680363874
transform 1 0 2504 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1680363874
transform -1 0 2544 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6680
timestamp 1680363874
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6688
timestamp 1680363874
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6689
timestamp 1680363874
transform 1 0 2560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6690
timestamp 1680363874
transform 1 0 2568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6691
timestamp 1680363874
transform 1 0 2576 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_414
timestamp 1680363874
transform -1 0 2600 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6692
timestamp 1680363874
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_358
timestamp 1680363874
transform 1 0 2608 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6693
timestamp 1680363874
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_415
timestamp 1680363874
transform 1 0 2712 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6694
timestamp 1680363874
transform 1 0 2728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6695
timestamp 1680363874
transform 1 0 2736 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_67
timestamp 1680363874
transform 1 0 2744 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6696
timestamp 1680363874
transform 1 0 2768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6698
timestamp 1680363874
transform 1 0 2776 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_31
timestamp 1680363874
transform 1 0 2784 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6701
timestamp 1680363874
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6702
timestamp 1680363874
transform 1 0 2824 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5452
timestamp 1680363874
transform 1 0 2852 0 1 1875
box -3 -3 3 3
use AND2X2  AND2X2_32
timestamp 1680363874
transform 1 0 2832 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6706
timestamp 1680363874
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6708
timestamp 1680363874
transform 1 0 2872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6710
timestamp 1680363874
transform 1 0 2880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6712
timestamp 1680363874
transform 1 0 2888 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_33
timestamp 1680363874
transform 1 0 2896 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6715
timestamp 1680363874
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6716
timestamp 1680363874
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6718
timestamp 1680363874
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_44
timestamp 1680363874
transform 1 0 2952 0 -1 1970
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_359
timestamp 1680363874
transform -1 0 3072 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5453
timestamp 1680363874
transform 1 0 3084 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_418
timestamp 1680363874
transform -1 0 3088 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6732
timestamp 1680363874
transform 1 0 3088 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5454
timestamp 1680363874
transform 1 0 3108 0 1 1875
box -3 -3 3 3
use FILL  FILL_6734
timestamp 1680363874
transform 1 0 3096 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_360
timestamp 1680363874
transform 1 0 3104 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5455
timestamp 1680363874
transform 1 0 3212 0 1 1875
box -3 -3 3 3
use FILL  FILL_6743
timestamp 1680363874
transform 1 0 3200 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_419
timestamp 1680363874
transform -1 0 3224 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6744
timestamp 1680363874
transform 1 0 3224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6745
timestamp 1680363874
transform 1 0 3232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6746
timestamp 1680363874
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6748
timestamp 1680363874
transform 1 0 3248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6750
timestamp 1680363874
transform 1 0 3256 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_34
timestamp 1680363874
transform 1 0 3264 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6756
timestamp 1680363874
transform 1 0 3296 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_35
timestamp 1680363874
transform 1 0 3304 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6757
timestamp 1680363874
transform 1 0 3336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6759
timestamp 1680363874
transform 1 0 3344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6761
timestamp 1680363874
transform 1 0 3352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6763
timestamp 1680363874
transform 1 0 3360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6765
timestamp 1680363874
transform 1 0 3368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6767
timestamp 1680363874
transform 1 0 3376 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_278
timestamp 1680363874
transform 1 0 3384 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6770
timestamp 1680363874
transform 1 0 3424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6771
timestamp 1680363874
transform 1 0 3432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6773
timestamp 1680363874
transform 1 0 3440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6775
timestamp 1680363874
transform 1 0 3448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6777
timestamp 1680363874
transform 1 0 3456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6779
timestamp 1680363874
transform 1 0 3464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6781
timestamp 1680363874
transform 1 0 3472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6783
timestamp 1680363874
transform 1 0 3480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6788
timestamp 1680363874
transform 1 0 3488 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_279
timestamp 1680363874
transform 1 0 3496 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6789
timestamp 1680363874
transform 1 0 3536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6791
timestamp 1680363874
transform 1 0 3544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6793
timestamp 1680363874
transform 1 0 3552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6795
timestamp 1680363874
transform 1 0 3560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6800
timestamp 1680363874
transform 1 0 3568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6801
timestamp 1680363874
transform 1 0 3576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6802
timestamp 1680363874
transform 1 0 3584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6803
timestamp 1680363874
transform 1 0 3592 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_218
timestamp 1680363874
transform 1 0 3600 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6804
timestamp 1680363874
transform 1 0 3640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6805
timestamp 1680363874
transform 1 0 3648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6806
timestamp 1680363874
transform 1 0 3656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6807
timestamp 1680363874
transform 1 0 3664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6808
timestamp 1680363874
transform 1 0 3672 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_70
timestamp 1680363874
transform -1 0 3704 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6809
timestamp 1680363874
transform 1 0 3704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6811
timestamp 1680363874
transform 1 0 3712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6813
timestamp 1680363874
transform 1 0 3720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6815
timestamp 1680363874
transform 1 0 3728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6817
timestamp 1680363874
transform 1 0 3736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6820
timestamp 1680363874
transform 1 0 3744 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_71
timestamp 1680363874
transform 1 0 3752 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6821
timestamp 1680363874
transform 1 0 3776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6822
timestamp 1680363874
transform 1 0 3784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6823
timestamp 1680363874
transform 1 0 3792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6825
timestamp 1680363874
transform 1 0 3800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6827
timestamp 1680363874
transform 1 0 3808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6829
timestamp 1680363874
transform 1 0 3816 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_45
timestamp 1680363874
transform 1 0 3824 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6834
timestamp 1680363874
transform 1 0 3848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6837
timestamp 1680363874
transform 1 0 3856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6838
timestamp 1680363874
transform 1 0 3864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6839
timestamp 1680363874
transform 1 0 3872 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_72
timestamp 1680363874
transform -1 0 3904 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6840
timestamp 1680363874
transform 1 0 3904 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_46
timestamp 1680363874
transform 1 0 3912 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6845
timestamp 1680363874
transform 1 0 3936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6847
timestamp 1680363874
transform 1 0 3944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6849
timestamp 1680363874
transform 1 0 3952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6851
timestamp 1680363874
transform 1 0 3960 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_48
timestamp 1680363874
transform 1 0 3968 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6854
timestamp 1680363874
transform 1 0 3992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6855
timestamp 1680363874
transform 1 0 4000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6857
timestamp 1680363874
transform 1 0 4008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6865
timestamp 1680363874
transform 1 0 4016 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_281
timestamp 1680363874
transform -1 0 4064 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6866
timestamp 1680363874
transform 1 0 4064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6868
timestamp 1680363874
transform 1 0 4072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6871
timestamp 1680363874
transform 1 0 4080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6872
timestamp 1680363874
transform 1 0 4088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6873
timestamp 1680363874
transform 1 0 4096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6874
timestamp 1680363874
transform 1 0 4104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6875
timestamp 1680363874
transform 1 0 4112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6876
timestamp 1680363874
transform 1 0 4120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6877
timestamp 1680363874
transform 1 0 4128 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_73
timestamp 1680363874
transform 1 0 4136 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6881
timestamp 1680363874
transform 1 0 4160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6882
timestamp 1680363874
transform 1 0 4168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6884
timestamp 1680363874
transform 1 0 4176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6886
timestamp 1680363874
transform 1 0 4184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6888
timestamp 1680363874
transform 1 0 4192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6895
timestamp 1680363874
transform 1 0 4200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6896
timestamp 1680363874
transform 1 0 4208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6897
timestamp 1680363874
transform 1 0 4216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6898
timestamp 1680363874
transform 1 0 4224 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_282
timestamp 1680363874
transform 1 0 4232 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6899
timestamp 1680363874
transform 1 0 4272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6900
timestamp 1680363874
transform 1 0 4280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6902
timestamp 1680363874
transform 1 0 4288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6904
timestamp 1680363874
transform 1 0 4296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6907
timestamp 1680363874
transform 1 0 4304 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_50
timestamp 1680363874
transform 1 0 4312 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6908
timestamp 1680363874
transform 1 0 4336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6909
timestamp 1680363874
transform 1 0 4344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6910
timestamp 1680363874
transform 1 0 4352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6912
timestamp 1680363874
transform 1 0 4360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6914
timestamp 1680363874
transform 1 0 4368 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_74
timestamp 1680363874
transform 1 0 4376 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6917
timestamp 1680363874
transform 1 0 4400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6918
timestamp 1680363874
transform 1 0 4408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6920
timestamp 1680363874
transform 1 0 4416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6922
timestamp 1680363874
transform 1 0 4424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6926
timestamp 1680363874
transform 1 0 4432 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_283
timestamp 1680363874
transform -1 0 4480 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6927
timestamp 1680363874
transform 1 0 4480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6928
timestamp 1680363874
transform 1 0 4488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6930
timestamp 1680363874
transform 1 0 4496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6932
timestamp 1680363874
transform 1 0 4504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6934
timestamp 1680363874
transform 1 0 4512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6936
timestamp 1680363874
transform 1 0 4520 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_75
timestamp 1680363874
transform 1 0 4528 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6941
timestamp 1680363874
transform 1 0 4552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6949
timestamp 1680363874
transform 1 0 4560 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_284
timestamp 1680363874
transform -1 0 4608 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6950
timestamp 1680363874
transform 1 0 4608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6952
timestamp 1680363874
transform 1 0 4616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6954
timestamp 1680363874
transform 1 0 4624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6956
timestamp 1680363874
transform 1 0 4632 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_223
timestamp 1680363874
transform 1 0 4640 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6963
timestamp 1680363874
transform 1 0 4680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6964
timestamp 1680363874
transform 1 0 4688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6965
timestamp 1680363874
transform 1 0 4696 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5456
timestamp 1680363874
transform 1 0 4748 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_363
timestamp 1680363874
transform 1 0 4704 0 -1 1970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_57
timestamp 1680363874
transform 1 0 4851 0 1 1870
box -10 -3 10 3
use M2_M1  M2_M1_6021
timestamp 1680363874
transform 1 0 108 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1680363874
transform 1 0 100 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5576
timestamp 1680363874
transform 1 0 100 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1680363874
transform 1 0 124 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6024
timestamp 1680363874
transform 1 0 124 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5500
timestamp 1680363874
transform 1 0 140 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1680363874
transform 1 0 156 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6031
timestamp 1680363874
transform 1 0 156 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5577
timestamp 1680363874
transform 1 0 148 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6137
timestamp 1680363874
transform 1 0 156 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5634
timestamp 1680363874
transform 1 0 156 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6032
timestamp 1680363874
transform 1 0 220 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5578
timestamp 1680363874
transform 1 0 220 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1680363874
transform 1 0 228 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6138
timestamp 1680363874
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5597
timestamp 1680363874
transform 1 0 244 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6025
timestamp 1680363874
transform 1 0 268 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5636
timestamp 1680363874
transform 1 0 268 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1680363874
transform 1 0 292 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6139
timestamp 1680363874
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1680363874
transform 1 0 340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1680363874
transform 1 0 316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1680363874
transform 1 0 332 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5580
timestamp 1680363874
transform 1 0 316 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1680363874
transform 1 0 340 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6140
timestamp 1680363874
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5598
timestamp 1680363874
transform 1 0 332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1680363874
transform 1 0 356 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6035
timestamp 1680363874
transform 1 0 412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1680363874
transform 1 0 436 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5637
timestamp 1680363874
transform 1 0 412 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1680363874
transform 1 0 468 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1680363874
transform 1 0 524 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1680363874
transform 1 0 620 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6036
timestamp 1680363874
transform 1 0 620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1680363874
transform 1 0 612 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5518
timestamp 1680363874
transform 1 0 652 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6037
timestamp 1680363874
transform 1 0 644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1680363874
transform 1 0 652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1680363874
transform 1 0 748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1680363874
transform 1 0 772 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5502
timestamp 1680363874
transform 1 0 940 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1680363874
transform 1 0 908 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6040
timestamp 1680363874
transform 1 0 900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1680363874
transform 1 0 948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1680363874
transform 1 0 988 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5599
timestamp 1680363874
transform 1 0 948 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1680363874
transform 1 0 1020 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6145
timestamp 1680363874
transform 1 0 1020 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5600
timestamp 1680363874
transform 1 0 1108 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6217
timestamp 1680363874
transform 1 0 1124 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1680363874
transform 1 0 1132 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5469
timestamp 1680363874
transform 1 0 1148 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1680363874
transform 1 0 1172 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1680363874
transform 1 0 1156 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6043
timestamp 1680363874
transform 1 0 1156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1680363874
transform 1 0 1172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1680363874
transform 1 0 1212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1680363874
transform 1 0 1220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1680363874
transform 1 0 1212 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5457
timestamp 1680363874
transform 1 0 1276 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1680363874
transform 1 0 1244 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1680363874
transform 1 0 1268 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1680363874
transform 1 0 1252 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6047
timestamp 1680363874
transform 1 0 1268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1680363874
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1680363874
transform 1 0 1236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1680363874
transform 1 0 1244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1680363874
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1680363874
transform 1 0 1276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1680363874
transform 1 0 1228 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5601
timestamp 1680363874
transform 1 0 1236 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1680363874
transform 1 0 1284 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6150
timestamp 1680363874
transform 1 0 1324 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5522
timestamp 1680363874
transform 1 0 1332 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6151
timestamp 1680363874
transform 1 0 1332 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5506
timestamp 1680363874
transform 1 0 1356 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6049
timestamp 1680363874
transform 1 0 1356 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5603
timestamp 1680363874
transform 1 0 1396 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1680363874
transform 1 0 1444 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6022
timestamp 1680363874
transform 1 0 1468 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1680363874
transform 1 0 1452 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5507
timestamp 1680363874
transform 1 0 1476 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6028
timestamp 1680363874
transform 1 0 1476 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1680363874
transform 1 0 1460 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5582
timestamp 1680363874
transform 1 0 1476 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6051
timestamp 1680363874
transform 1 0 1556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1680363874
transform 1 0 1532 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5604
timestamp 1680363874
transform 1 0 1532 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1680363874
transform 1 0 1660 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6052
timestamp 1680363874
transform 1 0 1660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1680363874
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1680363874
transform 1 0 1676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1680363874
transform 1 0 1684 0 1 1785
box -2 -2 2 2
use M3_M2  M3_M2_5471
timestamp 1680363874
transform 1 0 1748 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1680363874
transform 1 0 1740 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6055
timestamp 1680363874
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1680363874
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1680363874
transform 1 0 1740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1680363874
transform 1 0 1708 0 1 1785
box -2 -2 2 2
use M3_M2  M3_M2_5472
timestamp 1680363874
transform 1 0 1772 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6056
timestamp 1680363874
transform 1 0 1812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1680363874
transform 1 0 1820 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5583
timestamp 1680363874
transform 1 0 1812 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1680363874
transform 1 0 1804 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1680363874
transform 1 0 1844 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1680363874
transform 1 0 1860 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6058
timestamp 1680363874
transform 1 0 1844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1680363874
transform 1 0 1860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1680363874
transform 1 0 1836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1680363874
transform 1 0 1852 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5473
timestamp 1680363874
transform 1 0 1876 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6157
timestamp 1680363874
transform 1 0 1876 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5526
timestamp 1680363874
transform 1 0 1892 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6158
timestamp 1680363874
transform 1 0 1892 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5474
timestamp 1680363874
transform 1 0 1956 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1680363874
transform 1 0 1932 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6060
timestamp 1680363874
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1680363874
transform 1 0 1948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1680363874
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5584
timestamp 1680363874
transform 1 0 1924 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6159
timestamp 1680363874
transform 1 0 1956 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5585
timestamp 1680363874
transform 1 0 1964 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1680363874
transform 1 0 1996 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1680363874
transform 1 0 2044 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6063
timestamp 1680363874
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1680363874
transform 1 0 2044 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1680363874
transform 1 0 2020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1680363874
transform 1 0 2036 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5586
timestamp 1680363874
transform 1 0 2044 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1680363874
transform 1 0 2020 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1680363874
transform 1 0 2036 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6162
timestamp 1680363874
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5587
timestamp 1680363874
transform 1 0 2084 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1680363874
transform 1 0 2100 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1680363874
transform 1 0 2108 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1680363874
transform 1 0 2100 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6065
timestamp 1680363874
transform 1 0 2100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1680363874
transform 1 0 2124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1680363874
transform 1 0 2092 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5608
timestamp 1680363874
transform 1 0 2092 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6164
timestamp 1680363874
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1680363874
transform 1 0 2132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1680363874
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5530
timestamp 1680363874
transform 1 0 2148 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6067
timestamp 1680363874
transform 1 0 2156 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5588
timestamp 1680363874
transform 1 0 2156 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6068
timestamp 1680363874
transform 1 0 2196 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5557
timestamp 1680363874
transform 1 0 2204 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6167
timestamp 1680363874
transform 1 0 2188 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5531
timestamp 1680363874
transform 1 0 2228 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6069
timestamp 1680363874
transform 1 0 2220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1680363874
transform 1 0 2228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1680363874
transform 1 0 2228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1680363874
transform 1 0 2244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5476
timestamp 1680363874
transform 1 0 2268 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1680363874
transform 1 0 2284 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1680363874
transform 1 0 2268 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6071
timestamp 1680363874
transform 1 0 2284 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5559
timestamp 1680363874
transform 1 0 2292 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6170
timestamp 1680363874
transform 1 0 2276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1680363874
transform 1 0 2292 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5609
timestamp 1680363874
transform 1 0 2276 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1680363874
transform 1 0 2372 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6072
timestamp 1680363874
transform 1 0 2340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1680363874
transform 1 0 2316 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5610
timestamp 1680363874
transform 1 0 2340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1680363874
transform 1 0 2412 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1680363874
transform 1 0 2412 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6073
timestamp 1680363874
transform 1 0 2412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1680363874
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5638
timestamp 1680363874
transform 1 0 2404 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1680363874
transform 1 0 2436 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6075
timestamp 1680363874
transform 1 0 2444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1680363874
transform 1 0 2452 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5611
timestamp 1680363874
transform 1 0 2452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1680363874
transform 1 0 2468 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6076
timestamp 1680363874
transform 1 0 2476 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5492
timestamp 1680363874
transform 1 0 2516 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_6077
timestamp 1680363874
transform 1 0 2516 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5561
timestamp 1680363874
transform 1 0 2524 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6174
timestamp 1680363874
transform 1 0 2524 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5493
timestamp 1680363874
transform 1 0 2540 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1680363874
transform 1 0 2572 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1680363874
transform 1 0 2588 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1680363874
transform 1 0 2636 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1680363874
transform 1 0 2668 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6078
timestamp 1680363874
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1680363874
transform 1 0 2636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1680363874
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1680363874
transform 1 0 2660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1680363874
transform 1 0 2556 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5589
timestamp 1680363874
transform 1 0 2636 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1680363874
transform 1 0 2556 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6176
timestamp 1680363874
transform 1 0 2668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5613
timestamp 1680363874
transform 1 0 2668 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1680363874
transform 1 0 2660 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6082
timestamp 1680363874
transform 1 0 2684 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5562
timestamp 1680363874
transform 1 0 2692 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6083
timestamp 1680363874
transform 1 0 2700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1680363874
transform 1 0 2716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1680363874
transform 1 0 2708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1680363874
transform 1 0 2716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5614
timestamp 1680363874
transform 1 0 2708 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1680363874
transform 1 0 2716 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1680363874
transform 1 0 2732 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1680363874
transform 1 0 2732 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1680363874
transform 1 0 2780 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6085
timestamp 1680363874
transform 1 0 2780 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5615
timestamp 1680363874
transform 1 0 2780 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6179
timestamp 1680363874
transform 1 0 2804 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5537
timestamp 1680363874
transform 1 0 2820 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6086
timestamp 1680363874
transform 1 0 2820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1680363874
transform 1 0 2820 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5642
timestamp 1680363874
transform 1 0 2820 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1680363874
transform 1 0 2836 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6180
timestamp 1680363874
transform 1 0 2836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1680363874
transform 1 0 2860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1680363874
transform 1 0 2852 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5478
timestamp 1680363874
transform 1 0 2868 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1680363874
transform 1 0 2884 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6088
timestamp 1680363874
transform 1 0 2884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1680363874
transform 1 0 2892 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5509
timestamp 1680363874
transform 1 0 2916 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1680363874
transform 1 0 2908 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6089
timestamp 1680363874
transform 1 0 2908 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5563
timestamp 1680363874
transform 1 0 2924 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1680363874
transform 1 0 2948 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1680363874
transform 1 0 2940 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6090
timestamp 1680363874
transform 1 0 2940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1680363874
transform 1 0 2948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1680363874
transform 1 0 2932 0 1 1785
box -2 -2 2 2
use M3_M2  M3_M2_5496
timestamp 1680363874
transform 1 0 2988 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_6092
timestamp 1680363874
transform 1 0 2972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1680363874
transform 1 0 2988 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5591
timestamp 1680363874
transform 1 0 2964 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6183
timestamp 1680363874
transform 1 0 2972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5616
timestamp 1680363874
transform 1 0 2956 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1680363874
transform 1 0 2980 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6094
timestamp 1680363874
transform 1 0 3012 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5497
timestamp 1680363874
transform 1 0 3020 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1680363874
transform 1 0 3012 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1680363874
transform 1 0 3028 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1680363874
transform 1 0 3036 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6095
timestamp 1680363874
transform 1 0 3060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1680363874
transform 1 0 3052 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5643
timestamp 1680363874
transform 1 0 3052 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1680363874
transform 1 0 3076 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1680363874
transform 1 0 3068 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6185
timestamp 1680363874
transform 1 0 3076 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5541
timestamp 1680363874
transform 1 0 3124 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6096
timestamp 1680363874
transform 1 0 3124 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5542
timestamp 1680363874
transform 1 0 3156 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6097
timestamp 1680363874
transform 1 0 3156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1680363874
transform 1 0 3140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5594
timestamp 1680363874
transform 1 0 3148 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1680363874
transform 1 0 3156 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6098
timestamp 1680363874
transform 1 0 3188 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5463
timestamp 1680363874
transform 1 0 3228 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6099
timestamp 1680363874
transform 1 0 3228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1680363874
transform 1 0 3252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1680363874
transform 1 0 3212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1680363874
transform 1 0 3220 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1680363874
transform 1 0 3236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1680363874
transform 1 0 3244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5619
timestamp 1680363874
transform 1 0 3220 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1680363874
transform 1 0 3244 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1680363874
transform 1 0 3260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1680363874
transform 1 0 3276 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6221
timestamp 1680363874
transform 1 0 3292 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5464
timestamp 1680363874
transform 1 0 3316 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6029
timestamp 1680363874
transform 1 0 3316 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1680363874
transform 1 0 3308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1680363874
transform 1 0 3332 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1680363874
transform 1 0 3332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1680363874
transform 1 0 3324 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5512
timestamp 1680363874
transform 1 0 3356 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1680363874
transform 1 0 3388 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6222
timestamp 1680363874
transform 1 0 3396 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5480
timestamp 1680363874
transform 1 0 3420 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1680363874
transform 1 0 3460 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1680363874
transform 1 0 3436 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6103
timestamp 1680363874
transform 1 0 3436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1680363874
transform 1 0 3492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1680363874
transform 1 0 3412 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5622
timestamp 1680363874
transform 1 0 3412 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6105
timestamp 1680363874
transform 1 0 3508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1680363874
transform 1 0 3548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1680363874
transform 1 0 3572 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5567
timestamp 1680363874
transform 1 0 3580 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6107
timestamp 1680363874
transform 1 0 3596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1680363874
transform 1 0 3580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1680363874
transform 1 0 3588 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5568
timestamp 1680363874
transform 1 0 3612 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6108
timestamp 1680363874
transform 1 0 3636 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5569
timestamp 1680363874
transform 1 0 3676 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1680363874
transform 1 0 3692 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6109
timestamp 1680363874
transform 1 0 3684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1680363874
transform 1 0 3692 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5623
timestamp 1680363874
transform 1 0 3692 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1680363874
transform 1 0 3716 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6196
timestamp 1680363874
transform 1 0 3708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1680363874
transform 1 0 3716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5482
timestamp 1680363874
transform 1 0 3732 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6111
timestamp 1680363874
transform 1 0 3732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1680363874
transform 1 0 3756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1680363874
transform 1 0 3748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1680363874
transform 1 0 3764 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5624
timestamp 1680363874
transform 1 0 3764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1680363874
transform 1 0 3828 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1680363874
transform 1 0 3844 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6113
timestamp 1680363874
transform 1 0 3812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1680363874
transform 1 0 3788 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5625
timestamp 1680363874
transform 1 0 3860 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6114
timestamp 1680363874
transform 1 0 3876 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5626
timestamp 1680363874
transform 1 0 3876 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6201
timestamp 1680363874
transform 1 0 3892 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5513
timestamp 1680363874
transform 1 0 3924 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6202
timestamp 1680363874
transform 1 0 3916 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5627
timestamp 1680363874
transform 1 0 3916 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1680363874
transform 1 0 3932 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6115
timestamp 1680363874
transform 1 0 3932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1680363874
transform 1 0 3948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1680363874
transform 1 0 3940 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5644
timestamp 1680363874
transform 1 0 3940 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1680363874
transform 1 0 3980 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1680363874
transform 1 0 4004 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1680363874
transform 1 0 3996 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6117
timestamp 1680363874
transform 1 0 3996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1680363874
transform 1 0 3988 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5514
timestamp 1680363874
transform 1 0 4012 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1680363874
transform 1 0 4036 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_6118
timestamp 1680363874
transform 1 0 4020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1680363874
transform 1 0 4012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1680363874
transform 1 0 4020 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5466
timestamp 1680363874
transform 1 0 4068 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6119
timestamp 1680363874
transform 1 0 4068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1680363874
transform 1 0 4060 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5547
timestamp 1680363874
transform 1 0 4108 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1680363874
transform 1 0 4148 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6120
timestamp 1680363874
transform 1 0 4108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1680363874
transform 1 0 4116 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5571
timestamp 1680363874
transform 1 0 4124 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6122
timestamp 1680363874
transform 1 0 4148 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5572
timestamp 1680363874
transform 1 0 4196 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6206
timestamp 1680363874
transform 1 0 4092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1680363874
transform 1 0 4100 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5628
timestamp 1680363874
transform 1 0 4092 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6208
timestamp 1680363874
transform 1 0 4196 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5629
timestamp 1680363874
transform 1 0 4124 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1680363874
transform 1 0 4196 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1680363874
transform 1 0 4228 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1680363874
transform 1 0 4276 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1680363874
transform 1 0 4284 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6123
timestamp 1680363874
transform 1 0 4252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1680363874
transform 1 0 4300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1680363874
transform 1 0 4220 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5630
timestamp 1680363874
transform 1 0 4220 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1680363874
transform 1 0 4348 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6125
timestamp 1680363874
transform 1 0 4364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1680363874
transform 1 0 4420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1680363874
transform 1 0 4340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5631
timestamp 1680363874
transform 1 0 4340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1680363874
transform 1 0 4548 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1680363874
transform 1 0 4588 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1680363874
transform 1 0 4532 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1680363874
transform 1 0 4580 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6127
timestamp 1680363874
transform 1 0 4532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1680363874
transform 1 0 4572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1680363874
transform 1 0 4580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1680363874
transform 1 0 4492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1680363874
transform 1 0 4580 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5632
timestamp 1680363874
transform 1 0 4492 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6130
timestamp 1680363874
transform 1 0 4612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1680363874
transform 1 0 4604 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5515
timestamp 1680363874
transform 1 0 4660 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1680363874
transform 1 0 4652 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6131
timestamp 1680363874
transform 1 0 4636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1680363874
transform 1 0 4652 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5552
timestamp 1680363874
transform 1 0 4676 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6214
timestamp 1680363874
transform 1 0 4660 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5595
timestamp 1680363874
transform 1 0 4668 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6215
timestamp 1680363874
transform 1 0 4676 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5516
timestamp 1680363874
transform 1 0 4796 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1680363874
transform 1 0 4700 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1680363874
transform 1 0 4748 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6133
timestamp 1680363874
transform 1 0 4692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1680363874
transform 1 0 4700 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5573
timestamp 1680363874
transform 1 0 4716 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6135
timestamp 1680363874
transform 1 0 4748 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5574
timestamp 1680363874
transform 1 0 4780 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6136
timestamp 1680363874
transform 1 0 4796 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5575
timestamp 1680363874
transform 1 0 4812 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1680363874
transform 1 0 4700 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6216
timestamp 1680363874
transform 1 0 4716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5633
timestamp 1680363874
transform 1 0 4716 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1680363874
transform 1 0 4740 0 1 1785
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_58
timestamp 1680363874
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_6966
timestamp 1680363874
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_6968
timestamp 1680363874
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_6969
timestamp 1680363874
transform 1 0 88 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_49
timestamp 1680363874
transform -1 0 128 0 1 1770
box -8 -3 40 105
use FILL  FILL_6970
timestamp 1680363874
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_6971
timestamp 1680363874
transform 1 0 136 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_424
timestamp 1680363874
transform -1 0 160 0 1 1770
box -9 -3 26 105
use FILL  FILL_6972
timestamp 1680363874
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_6978
timestamp 1680363874
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_6980
timestamp 1680363874
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_6982
timestamp 1680363874
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_6984
timestamp 1680363874
transform 1 0 192 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_426
timestamp 1680363874
transform -1 0 216 0 1 1770
box -9 -3 26 105
use FILL  FILL_6985
timestamp 1680363874
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_6990
timestamp 1680363874
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_6992
timestamp 1680363874
transform 1 0 232 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_144
timestamp 1680363874
transform 1 0 240 0 1 1770
box -8 -3 34 105
use FILL  FILL_6994
timestamp 1680363874
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_6995
timestamp 1680363874
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_6996
timestamp 1680363874
transform 1 0 288 0 1 1770
box -8 -3 16 105
use FILL  FILL_6997
timestamp 1680363874
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_6998
timestamp 1680363874
transform 1 0 304 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_36
timestamp 1680363874
transform -1 0 344 0 1 1770
box -8 -3 40 105
use FILL  FILL_6999
timestamp 1680363874
transform 1 0 344 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_364
timestamp 1680363874
transform -1 0 448 0 1 1770
box -8 -3 104 105
use FILL  FILL_7000
timestamp 1680363874
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_7001
timestamp 1680363874
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_7002
timestamp 1680363874
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7008
timestamp 1680363874
transform 1 0 472 0 1 1770
box -8 -3 16 105
use FILL  FILL_7010
timestamp 1680363874
transform 1 0 480 0 1 1770
box -8 -3 16 105
use FILL  FILL_7011
timestamp 1680363874
transform 1 0 488 0 1 1770
box -8 -3 16 105
use FILL  FILL_7012
timestamp 1680363874
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7013
timestamp 1680363874
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7014
timestamp 1680363874
transform 1 0 512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7015
timestamp 1680363874
transform 1 0 520 0 1 1770
box -8 -3 16 105
use FILL  FILL_7016
timestamp 1680363874
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_7017
timestamp 1680363874
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_7018
timestamp 1680363874
transform 1 0 544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7019
timestamp 1680363874
transform 1 0 552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7020
timestamp 1680363874
transform 1 0 560 0 1 1770
box -8 -3 16 105
use FILL  FILL_7021
timestamp 1680363874
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_7022
timestamp 1680363874
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_7024
timestamp 1680363874
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7026
timestamp 1680363874
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7028
timestamp 1680363874
transform 1 0 600 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_37
timestamp 1680363874
transform 1 0 608 0 1 1770
box -8 -3 40 105
use FILL  FILL_7030
timestamp 1680363874
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_7031
timestamp 1680363874
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_7032
timestamp 1680363874
transform 1 0 656 0 1 1770
box -8 -3 16 105
use FILL  FILL_7033
timestamp 1680363874
transform 1 0 664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7034
timestamp 1680363874
transform 1 0 672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7035
timestamp 1680363874
transform 1 0 680 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_368
timestamp 1680363874
transform -1 0 784 0 1 1770
box -8 -3 104 105
use FILL  FILL_7036
timestamp 1680363874
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_7045
timestamp 1680363874
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_7046
timestamp 1680363874
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_7047
timestamp 1680363874
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_7048
timestamp 1680363874
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_7049
timestamp 1680363874
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_7050
timestamp 1680363874
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_7051
timestamp 1680363874
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_7052
timestamp 1680363874
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_7053
timestamp 1680363874
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_7054
timestamp 1680363874
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_7055
timestamp 1680363874
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7056
timestamp 1680363874
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_7057
timestamp 1680363874
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_7059
timestamp 1680363874
transform 1 0 896 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_370
timestamp 1680363874
transform -1 0 1000 0 1 1770
box -8 -3 104 105
use FILL  FILL_7060
timestamp 1680363874
transform 1 0 1000 0 1 1770
box -8 -3 16 105
use FILL  FILL_7061
timestamp 1680363874
transform 1 0 1008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7062
timestamp 1680363874
transform 1 0 1016 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5647
timestamp 1680363874
transform 1 0 1052 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_427
timestamp 1680363874
transform 1 0 1024 0 1 1770
box -9 -3 26 105
use FILL  FILL_7063
timestamp 1680363874
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7064
timestamp 1680363874
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5648
timestamp 1680363874
transform 1 0 1068 0 1 1775
box -3 -3 3 3
use FILL  FILL_7073
timestamp 1680363874
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_7075
timestamp 1680363874
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_7077
timestamp 1680363874
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_7079
timestamp 1680363874
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7081
timestamp 1680363874
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7083
timestamp 1680363874
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7084
timestamp 1680363874
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7085
timestamp 1680363874
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_7086
timestamp 1680363874
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_7087
timestamp 1680363874
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_224
timestamp 1680363874
transform -1 0 1176 0 1 1770
box -8 -3 46 105
use FILL  FILL_7088
timestamp 1680363874
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_7095
timestamp 1680363874
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_7097
timestamp 1680363874
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7099
timestamp 1680363874
transform 1 0 1200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7101
timestamp 1680363874
transform 1 0 1208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7102
timestamp 1680363874
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7103
timestamp 1680363874
transform 1 0 1224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7104
timestamp 1680363874
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_286
timestamp 1680363874
transform 1 0 1240 0 1 1770
box -8 -3 46 105
use FILL  FILL_7105
timestamp 1680363874
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_7111
timestamp 1680363874
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use FILL  FILL_7113
timestamp 1680363874
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_428
timestamp 1680363874
transform -1 0 1320 0 1 1770
box -9 -3 26 105
use FILL  FILL_7114
timestamp 1680363874
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_7115
timestamp 1680363874
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_7116
timestamp 1680363874
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_7117
timestamp 1680363874
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_7118
timestamp 1680363874
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_429
timestamp 1680363874
transform 1 0 1360 0 1 1770
box -9 -3 26 105
use FILL  FILL_7119
timestamp 1680363874
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_7120
timestamp 1680363874
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7121
timestamp 1680363874
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_7122
timestamp 1680363874
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_7123
timestamp 1680363874
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5649
timestamp 1680363874
transform 1 0 1428 0 1 1775
box -3 -3 3 3
use FILL  FILL_7127
timestamp 1680363874
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_7128
timestamp 1680363874
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7129
timestamp 1680363874
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7130
timestamp 1680363874
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1680363874
transform 1 0 1448 0 1 1770
box -8 -3 40 105
use FILL  FILL_7131
timestamp 1680363874
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_7132
timestamp 1680363874
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_7133
timestamp 1680363874
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7134
timestamp 1680363874
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7135
timestamp 1680363874
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_374
timestamp 1680363874
transform 1 0 1520 0 1 1770
box -8 -3 104 105
use FILL  FILL_7137
timestamp 1680363874
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_7146
timestamp 1680363874
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_7148
timestamp 1680363874
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_7150
timestamp 1680363874
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_430
timestamp 1680363874
transform 1 0 1648 0 1 1770
box -9 -3 26 105
use FILL  FILL_7152
timestamp 1680363874
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7154
timestamp 1680363874
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7156
timestamp 1680363874
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7158
timestamp 1680363874
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_7160
timestamp 1680363874
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_7162
timestamp 1680363874
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_225
timestamp 1680363874
transform -1 0 1752 0 1 1770
box -8 -3 46 105
use FILL  FILL_7163
timestamp 1680363874
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_7164
timestamp 1680363874
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_7165
timestamp 1680363874
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_7166
timestamp 1680363874
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_7167
timestamp 1680363874
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use FILL  FILL_7168
timestamp 1680363874
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_7169
timestamp 1680363874
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_7170
timestamp 1680363874
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_7171
timestamp 1680363874
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_7175
timestamp 1680363874
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_289
timestamp 1680363874
transform 1 0 1832 0 1 1770
box -8 -3 46 105
use FILL  FILL_7177
timestamp 1680363874
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7178
timestamp 1680363874
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_7179
timestamp 1680363874
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_7180
timestamp 1680363874
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_7181
timestamp 1680363874
transform 1 0 1904 0 1 1770
box -8 -3 16 105
use FILL  FILL_7182
timestamp 1680363874
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7183
timestamp 1680363874
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_226
timestamp 1680363874
transform -1 0 1968 0 1 1770
box -8 -3 46 105
use FILL  FILL_7184
timestamp 1680363874
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_7191
timestamp 1680363874
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_7193
timestamp 1680363874
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_7194
timestamp 1680363874
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_7195
timestamp 1680363874
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_227
timestamp 1680363874
transform 1 0 2008 0 1 1770
box -8 -3 46 105
use FILL  FILL_7196
timestamp 1680363874
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5650
timestamp 1680363874
transform 1 0 2068 0 1 1775
box -3 -3 3 3
use FILL  FILL_7197
timestamp 1680363874
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_7198
timestamp 1680363874
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_7199
timestamp 1680363874
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_7200
timestamp 1680363874
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7201
timestamp 1680363874
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_290
timestamp 1680363874
transform 1 0 2096 0 1 1770
box -8 -3 46 105
use FILL  FILL_7202
timestamp 1680363874
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use FILL  FILL_7203
timestamp 1680363874
transform 1 0 2144 0 1 1770
box -8 -3 16 105
use FILL  FILL_7204
timestamp 1680363874
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_7205
timestamp 1680363874
transform 1 0 2160 0 1 1770
box -8 -3 16 105
use FILL  FILL_7206
timestamp 1680363874
transform 1 0 2168 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_228
timestamp 1680363874
transform -1 0 2216 0 1 1770
box -8 -3 46 105
use FILL  FILL_7207
timestamp 1680363874
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7208
timestamp 1680363874
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7212
timestamp 1680363874
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_7214
timestamp 1680363874
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use FILL  FILL_7216
timestamp 1680363874
transform 1 0 2248 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_291
timestamp 1680363874
transform 1 0 2256 0 1 1770
box -8 -3 46 105
use FILL  FILL_7218
timestamp 1680363874
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5651
timestamp 1680363874
transform 1 0 2340 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1680363874
transform 1 0 2364 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_379
timestamp 1680363874
transform 1 0 2304 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_434
timestamp 1680363874
transform 1 0 2400 0 1 1770
box -9 -3 26 105
use FILL  FILL_7219
timestamp 1680363874
transform 1 0 2416 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_38
timestamp 1680363874
transform -1 0 2456 0 1 1770
box -8 -3 40 105
use FILL  FILL_7220
timestamp 1680363874
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_7221
timestamp 1680363874
transform 1 0 2464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7222
timestamp 1680363874
transform 1 0 2472 0 1 1770
box -8 -3 16 105
use FILL  FILL_7223
timestamp 1680363874
transform 1 0 2480 0 1 1770
box -8 -3 16 105
use FILL  FILL_7224
timestamp 1680363874
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_39
timestamp 1680363874
transform -1 0 2528 0 1 1770
box -8 -3 40 105
use FILL  FILL_7225
timestamp 1680363874
transform 1 0 2528 0 1 1770
box -8 -3 16 105
use FILL  FILL_7226
timestamp 1680363874
transform 1 0 2536 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_381
timestamp 1680363874
transform 1 0 2544 0 1 1770
box -8 -3 104 105
use AND2X2  AND2X2_40
timestamp 1680363874
transform -1 0 2672 0 1 1770
box -8 -3 40 105
use FILL  FILL_7242
timestamp 1680363874
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_41
timestamp 1680363874
transform -1 0 2712 0 1 1770
box -8 -3 40 105
use FILL  FILL_7243
timestamp 1680363874
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use FILL  FILL_7244
timestamp 1680363874
transform 1 0 2720 0 1 1770
box -8 -3 16 105
use FILL  FILL_7245
timestamp 1680363874
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_435
timestamp 1680363874
transform 1 0 2736 0 1 1770
box -9 -3 26 105
use FILL  FILL_7246
timestamp 1680363874
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_76
timestamp 1680363874
transform 1 0 2760 0 1 1770
box -8 -3 32 105
use FILL  FILL_7247
timestamp 1680363874
transform 1 0 2784 0 1 1770
box -8 -3 16 105
use FILL  FILL_7248
timestamp 1680363874
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_77
timestamp 1680363874
transform -1 0 2824 0 1 1770
box -8 -3 32 105
use FILL  FILL_7249
timestamp 1680363874
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_7250
timestamp 1680363874
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_436
timestamp 1680363874
transform -1 0 2856 0 1 1770
box -9 -3 26 105
use FILL  FILL_7251
timestamp 1680363874
transform 1 0 2856 0 1 1770
box -8 -3 16 105
use FILL  FILL_7252
timestamp 1680363874
transform 1 0 2864 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_437
timestamp 1680363874
transform -1 0 2888 0 1 1770
box -9 -3 26 105
use FILL  FILL_7253
timestamp 1680363874
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5653
timestamp 1680363874
transform 1 0 2932 0 1 1775
box -3 -3 3 3
use AND2X2  AND2X2_42
timestamp 1680363874
transform 1 0 2896 0 1 1770
box -8 -3 40 105
use FILL  FILL_7254
timestamp 1680363874
transform 1 0 2928 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_438
timestamp 1680363874
transform 1 0 2936 0 1 1770
box -9 -3 26 105
use FILL  FILL_7255
timestamp 1680363874
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5654
timestamp 1680363874
transform 1 0 2972 0 1 1775
box -3 -3 3 3
use FILL  FILL_7267
timestamp 1680363874
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_230
timestamp 1680363874
transform 1 0 2968 0 1 1770
box -8 -3 46 105
use FILL  FILL_7268
timestamp 1680363874
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7269
timestamp 1680363874
transform 1 0 3016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7270
timestamp 1680363874
transform 1 0 3024 0 1 1770
box -8 -3 16 105
use FILL  FILL_7271
timestamp 1680363874
transform 1 0 3032 0 1 1770
box -8 -3 16 105
use FILL  FILL_7272
timestamp 1680363874
transform 1 0 3040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7273
timestamp 1680363874
transform 1 0 3048 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_59
timestamp 1680363874
transform 1 0 3056 0 1 1770
box -5 -3 28 105
use FILL  FILL_7274
timestamp 1680363874
transform 1 0 3080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7275
timestamp 1680363874
transform 1 0 3088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7276
timestamp 1680363874
transform 1 0 3096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7280
timestamp 1680363874
transform 1 0 3104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7281
timestamp 1680363874
transform 1 0 3112 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_65
timestamp 1680363874
transform 1 0 3120 0 1 1770
box -5 -3 28 105
use FILL  FILL_7282
timestamp 1680363874
transform 1 0 3144 0 1 1770
box -8 -3 16 105
use FILL  FILL_7286
timestamp 1680363874
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_67
timestamp 1680363874
transform 1 0 3160 0 1 1770
box -5 -3 28 105
use FILL  FILL_7288
timestamp 1680363874
transform 1 0 3184 0 1 1770
box -8 -3 16 105
use FILL  FILL_7289
timestamp 1680363874
transform 1 0 3192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7290
timestamp 1680363874
transform 1 0 3200 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_231
timestamp 1680363874
transform 1 0 3208 0 1 1770
box -8 -3 46 105
use FILL  FILL_7291
timestamp 1680363874
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_7292
timestamp 1680363874
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use FILL  FILL_7293
timestamp 1680363874
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_7294
timestamp 1680363874
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_7295
timestamp 1680363874
transform 1 0 3280 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_78
timestamp 1680363874
transform 1 0 3288 0 1 1770
box -8 -3 32 105
use FILL  FILL_7296
timestamp 1680363874
transform 1 0 3312 0 1 1770
box -8 -3 16 105
use FILL  FILL_7303
timestamp 1680363874
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use FILL  FILL_7305
timestamp 1680363874
transform 1 0 3328 0 1 1770
box -8 -3 16 105
use FILL  FILL_7307
timestamp 1680363874
transform 1 0 3336 0 1 1770
box -8 -3 16 105
use FILL  FILL_7309
timestamp 1680363874
transform 1 0 3344 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_79
timestamp 1680363874
transform -1 0 3376 0 1 1770
box -8 -3 32 105
use FILL  FILL_7310
timestamp 1680363874
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_7312
timestamp 1680363874
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7314
timestamp 1680363874
transform 1 0 3392 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_384
timestamp 1680363874
transform 1 0 3400 0 1 1770
box -8 -3 104 105
use FILL  FILL_7316
timestamp 1680363874
transform 1 0 3496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7317
timestamp 1680363874
transform 1 0 3504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7318
timestamp 1680363874
transform 1 0 3512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7327
timestamp 1680363874
transform 1 0 3520 0 1 1770
box -8 -3 16 105
use FILL  FILL_7329
timestamp 1680363874
transform 1 0 3528 0 1 1770
box -8 -3 16 105
use FILL  FILL_7331
timestamp 1680363874
transform 1 0 3536 0 1 1770
box -8 -3 16 105
use FILL  FILL_7333
timestamp 1680363874
transform 1 0 3544 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_233
timestamp 1680363874
transform 1 0 3552 0 1 1770
box -8 -3 46 105
use FILL  FILL_7335
timestamp 1680363874
transform 1 0 3592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7342
timestamp 1680363874
transform 1 0 3600 0 1 1770
box -8 -3 16 105
use FILL  FILL_7344
timestamp 1680363874
transform 1 0 3608 0 1 1770
box -8 -3 16 105
use FILL  FILL_7346
timestamp 1680363874
transform 1 0 3616 0 1 1770
box -8 -3 16 105
use FILL  FILL_7348
timestamp 1680363874
transform 1 0 3624 0 1 1770
box -8 -3 16 105
use FILL  FILL_7350
timestamp 1680363874
transform 1 0 3632 0 1 1770
box -8 -3 16 105
use FILL  FILL_7352
timestamp 1680363874
transform 1 0 3640 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_441
timestamp 1680363874
transform 1 0 3648 0 1 1770
box -9 -3 26 105
use FILL  FILL_7353
timestamp 1680363874
transform 1 0 3664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7354
timestamp 1680363874
transform 1 0 3672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7355
timestamp 1680363874
transform 1 0 3680 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_68
timestamp 1680363874
transform 1 0 3688 0 1 1770
box -5 -3 28 105
use FILL  FILL_7356
timestamp 1680363874
transform 1 0 3712 0 1 1770
box -8 -3 16 105
use FILL  FILL_7357
timestamp 1680363874
transform 1 0 3720 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_292
timestamp 1680363874
transform 1 0 3728 0 1 1770
box -8 -3 46 105
use FILL  FILL_7358
timestamp 1680363874
transform 1 0 3768 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_386
timestamp 1680363874
transform 1 0 3776 0 1 1770
box -8 -3 104 105
use FILL  FILL_7364
timestamp 1680363874
transform 1 0 3872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7365
timestamp 1680363874
transform 1 0 3880 0 1 1770
box -8 -3 16 105
use FILL  FILL_7366
timestamp 1680363874
transform 1 0 3888 0 1 1770
box -8 -3 16 105
use FILL  FILL_7367
timestamp 1680363874
transform 1 0 3896 0 1 1770
box -8 -3 16 105
use FILL  FILL_7377
timestamp 1680363874
transform 1 0 3904 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_69
timestamp 1680363874
transform -1 0 3936 0 1 1770
box -5 -3 28 105
use FILL  FILL_7378
timestamp 1680363874
transform 1 0 3936 0 1 1770
box -8 -3 16 105
use FILL  FILL_7379
timestamp 1680363874
transform 1 0 3944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7380
timestamp 1680363874
transform 1 0 3952 0 1 1770
box -8 -3 16 105
use FILL  FILL_7381
timestamp 1680363874
transform 1 0 3960 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_80
timestamp 1680363874
transform -1 0 3992 0 1 1770
box -8 -3 32 105
use M3_M2  M3_M2_5655
timestamp 1680363874
transform 1 0 4020 0 1 1775
box -3 -3 3 3
use BUFX2  BUFX2_70
timestamp 1680363874
transform 1 0 3992 0 1 1770
box -5 -3 28 105
use NOR2X1  NOR2X1_81
timestamp 1680363874
transform -1 0 4040 0 1 1770
box -8 -3 32 105
use FILL  FILL_7382
timestamp 1680363874
transform 1 0 4040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7383
timestamp 1680363874
transform 1 0 4048 0 1 1770
box -8 -3 16 105
use FILL  FILL_7393
timestamp 1680363874
transform 1 0 4056 0 1 1770
box -8 -3 16 105
use FILL  FILL_7395
timestamp 1680363874
transform 1 0 4064 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_72
timestamp 1680363874
transform 1 0 4072 0 1 1770
box -5 -3 28 105
use INVX2  INVX2_444
timestamp 1680363874
transform 1 0 4096 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5656
timestamp 1680363874
transform 1 0 4164 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1680363874
transform 1 0 4212 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_387
timestamp 1680363874
transform -1 0 4208 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_388
timestamp 1680363874
transform 1 0 4208 0 1 1770
box -8 -3 104 105
use FILL  FILL_7397
timestamp 1680363874
transform 1 0 4304 0 1 1770
box -8 -3 16 105
use FILL  FILL_7398
timestamp 1680363874
transform 1 0 4312 0 1 1770
box -8 -3 16 105
use FILL  FILL_7413
timestamp 1680363874
transform 1 0 4320 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_389
timestamp 1680363874
transform 1 0 4328 0 1 1770
box -8 -3 104 105
use FILL  FILL_7415
timestamp 1680363874
transform 1 0 4424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7422
timestamp 1680363874
transform 1 0 4432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7424
timestamp 1680363874
transform 1 0 4440 0 1 1770
box -8 -3 16 105
use FILL  FILL_7426
timestamp 1680363874
transform 1 0 4448 0 1 1770
box -8 -3 16 105
use FILL  FILL_7428
timestamp 1680363874
transform 1 0 4456 0 1 1770
box -8 -3 16 105
use FILL  FILL_7430
timestamp 1680363874
transform 1 0 4464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7432
timestamp 1680363874
transform 1 0 4472 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_390
timestamp 1680363874
transform 1 0 4480 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_447
timestamp 1680363874
transform 1 0 4576 0 1 1770
box -9 -3 26 105
use FILL  FILL_7433
timestamp 1680363874
transform 1 0 4592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7443
timestamp 1680363874
transform 1 0 4600 0 1 1770
box -8 -3 16 105
use FILL  FILL_7445
timestamp 1680363874
transform 1 0 4608 0 1 1770
box -8 -3 16 105
use FILL  FILL_7447
timestamp 1680363874
transform 1 0 4616 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5658
timestamp 1680363874
transform 1 0 4636 0 1 1775
box -3 -3 3 3
use FILL  FILL_7449
timestamp 1680363874
transform 1 0 4624 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_241
timestamp 1680363874
transform 1 0 4632 0 1 1770
box -8 -3 46 105
use FILL  FILL_7451
timestamp 1680363874
transform 1 0 4672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7453
timestamp 1680363874
transform 1 0 4680 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_449
timestamp 1680363874
transform 1 0 4688 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5659
timestamp 1680363874
transform 1 0 4764 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_391
timestamp 1680363874
transform 1 0 4704 0 1 1770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_59
timestamp 1680363874
transform 1 0 4827 0 1 1770
box -10 -3 10 3
use M2_M1  M2_M1_6229
timestamp 1680363874
transform 1 0 100 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1680363874
transform 1 0 100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1680363874
transform 1 0 140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1680363874
transform 1 0 148 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1680363874
transform 1 0 164 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5704
timestamp 1680363874
transform 1 0 348 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6230
timestamp 1680363874
transform 1 0 284 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5759
timestamp 1680363874
transform 1 0 284 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1680363874
transform 1 0 380 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1680363874
transform 1 0 436 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6231
timestamp 1680363874
transform 1 0 380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1680363874
transform 1 0 332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1680363874
transform 1 0 364 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5760
timestamp 1680363874
transform 1 0 380 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6311
timestamp 1680363874
transform 1 0 404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1680363874
transform 1 0 476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5662
timestamp 1680363874
transform 1 0 492 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1680363874
transform 1 0 508 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6232
timestamp 1680363874
transform 1 0 492 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5761
timestamp 1680363874
transform 1 0 492 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6313
timestamp 1680363874
transform 1 0 516 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5762
timestamp 1680363874
transform 1 0 564 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6314
timestamp 1680363874
transform 1 0 580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1680363874
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5851
timestamp 1680363874
transform 1 0 596 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1680363874
transform 1 0 676 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1680363874
transform 1 0 700 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6228
timestamp 1680363874
transform 1 0 732 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1680363874
transform 1 0 628 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5763
timestamp 1680363874
transform 1 0 628 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6315
timestamp 1680363874
transform 1 0 636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1680363874
transform 1 0 644 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5764
timestamp 1680363874
transform 1 0 676 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1680363874
transform 1 0 644 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6317
timestamp 1680363874
transform 1 0 756 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5706
timestamp 1680363874
transform 1 0 772 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1680363874
transform 1 0 788 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1680363874
transform 1 0 812 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1680363874
transform 1 0 804 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1680363874
transform 1 0 884 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6235
timestamp 1680363874
transform 1 0 804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1680363874
transform 1 0 852 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1680363874
transform 1 0 924 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5665
timestamp 1680363874
transform 1 0 1020 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1680363874
transform 1 0 988 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6236
timestamp 1680363874
transform 1 0 964 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5765
timestamp 1680363874
transform 1 0 964 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1680363874
transform 1 0 996 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6320
timestamp 1680363874
transform 1 0 1012 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5788
timestamp 1680363874
transform 1 0 1012 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1680363874
transform 1 0 1052 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6321
timestamp 1680363874
transform 1 0 1052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1680363874
transform 1 0 1076 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5709
timestamp 1680363874
transform 1 0 1092 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6237
timestamp 1680363874
transform 1 0 1092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1680363874
transform 1 0 1116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1680363874
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1680363874
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5789
timestamp 1680363874
transform 1 0 1116 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1680363874
transform 1 0 1100 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6239
timestamp 1680363874
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5710
timestamp 1680363874
transform 1 0 1156 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6240
timestamp 1680363874
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5829
timestamp 1680363874
transform 1 0 1196 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6241
timestamp 1680363874
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1680363874
transform 1 0 1228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1680363874
transform 1 0 1220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1680363874
transform 1 0 1236 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5790
timestamp 1680363874
transform 1 0 1228 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1680363874
transform 1 0 1284 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6243
timestamp 1680363874
transform 1 0 1276 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5737
timestamp 1680363874
transform 1 0 1308 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6327
timestamp 1680363874
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5667
timestamp 1680363874
transform 1 0 1332 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1680363874
transform 1 0 1388 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1680363874
transform 1 0 1380 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1680363874
transform 1 0 1324 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6244
timestamp 1680363874
transform 1 0 1396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1680363874
transform 1 0 1348 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5767
timestamp 1680363874
transform 1 0 1364 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1680363874
transform 1 0 1396 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1680363874
transform 1 0 1348 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1680363874
transform 1 0 1508 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1680363874
transform 1 0 1444 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6245
timestamp 1680363874
transform 1 0 1428 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5739
timestamp 1680363874
transform 1 0 1476 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6329
timestamp 1680363874
transform 1 0 1476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5670
timestamp 1680363874
transform 1 0 1524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1680363874
transform 1 0 1532 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6246
timestamp 1680363874
transform 1 0 1524 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5769
timestamp 1680363874
transform 1 0 1516 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1680363874
transform 1 0 1556 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6247
timestamp 1680363874
transform 1 0 1564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1680363874
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1680363874
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1680363874
transform 1 0 1548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1680363874
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5770
timestamp 1680363874
transform 1 0 1564 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6332
timestamp 1680363874
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5792
timestamp 1680363874
transform 1 0 1548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1680363874
transform 1 0 1572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1680363874
transform 1 0 1588 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6333
timestamp 1680363874
transform 1 0 1628 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5831
timestamp 1680363874
transform 1 0 1628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1680363874
transform 1 0 1660 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1680363874
transform 1 0 1780 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1680363874
transform 1 0 1756 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1680363874
transform 1 0 1780 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6250
timestamp 1680363874
transform 1 0 1804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1680363874
transform 1 0 1716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1680363874
transform 1 0 1724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1680363874
transform 1 0 1756 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5795
timestamp 1680363874
transform 1 0 1756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1680363874
transform 1 0 1804 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1680363874
transform 1 0 1756 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1680363874
transform 1 0 1796 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1680363874
transform 1 0 1820 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1680363874
transform 1 0 1844 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1680363874
transform 1 0 1836 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1680363874
transform 1 0 1892 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1680363874
transform 1 0 1844 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6251
timestamp 1680363874
transform 1 0 1844 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5743
timestamp 1680363874
transform 1 0 1876 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1680363874
transform 1 0 1844 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6337
timestamp 1680363874
transform 1 0 1876 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5797
timestamp 1680363874
transform 1 0 1876 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1680363874
transform 1 0 1908 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1680363874
transform 1 0 1860 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1680363874
transform 1 0 1892 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1680363874
transform 1 0 1852 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5869
timestamp 1680363874
transform 1 0 1884 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6338
timestamp 1680363874
transform 1 0 1940 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5687
timestamp 1680363874
transform 1 0 2156 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1680363874
transform 1 0 1996 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1680363874
transform 1 0 2076 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1680363874
transform 1 0 2108 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6252
timestamp 1680363874
transform 1 0 1996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1680363874
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5870
timestamp 1680363874
transform 1 0 2004 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1680363874
transform 1 0 2044 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6253
timestamp 1680363874
transform 1 0 2108 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5744
timestamp 1680363874
transform 1 0 2172 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6340
timestamp 1680363874
transform 1 0 2092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1680363874
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5798
timestamp 1680363874
transform 1 0 2156 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1680363874
transform 1 0 2196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1680363874
transform 1 0 2220 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6342
timestamp 1680363874
transform 1 0 2220 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5800
timestamp 1680363874
transform 1 0 2220 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1680363874
transform 1 0 2260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1680363874
transform 1 0 2252 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1680363874
transform 1 0 2276 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1680363874
transform 1 0 2292 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1680363874
transform 1 0 2316 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6254
timestamp 1680363874
transform 1 0 2284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1680363874
transform 1 0 2300 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5746
timestamp 1680363874
transform 1 0 2308 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6343
timestamp 1680363874
transform 1 0 2276 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5773
timestamp 1680363874
transform 1 0 2284 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6344
timestamp 1680363874
transform 1 0 2292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1680363874
transform 1 0 2308 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5801
timestamp 1680363874
transform 1 0 2300 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6407
timestamp 1680363874
transform 1 0 2324 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5690
timestamp 1680363874
transform 1 0 2356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1680363874
transform 1 0 2348 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6346
timestamp 1680363874
transform 1 0 2388 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5774
timestamp 1680363874
transform 1 0 2396 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1680363874
transform 1 0 2388 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6408
timestamp 1680363874
transform 1 0 2404 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1680363874
transform 1 0 2396 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5691
timestamp 1680363874
transform 1 0 2428 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1680363874
transform 1 0 2444 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6256
timestamp 1680363874
transform 1 0 2452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1680363874
transform 1 0 2500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1680363874
transform 1 0 2532 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5804
timestamp 1680363874
transform 1 0 2500 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1680363874
transform 1 0 2484 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1680363874
transform 1 0 2532 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1680363874
transform 1 0 2556 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6349
timestamp 1680363874
transform 1 0 2548 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5747
timestamp 1680363874
transform 1 0 2564 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6350
timestamp 1680363874
transform 1 0 2572 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5805
timestamp 1680363874
transform 1 0 2588 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6257
timestamp 1680363874
transform 1 0 2604 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5719
timestamp 1680363874
transform 1 0 2620 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6351
timestamp 1680363874
transform 1 0 2620 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1680363874
transform 1 0 2612 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5806
timestamp 1680363874
transform 1 0 2620 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1680363874
transform 1 0 2652 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1680363874
transform 1 0 2716 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1680363874
transform 1 0 2652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1680363874
transform 1 0 2724 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6258
timestamp 1680363874
transform 1 0 2652 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5674
timestamp 1680363874
transform 1 0 2788 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6259
timestamp 1680363874
transform 1 0 2772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1680363874
transform 1 0 2676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1680363874
transform 1 0 2732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1680363874
transform 1 0 2748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1680363874
transform 1 0 2636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1680363874
transform 1 0 2628 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5855
timestamp 1680363874
transform 1 0 2628 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1680363874
transform 1 0 2684 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1680363874
transform 1 0 2732 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1680363874
transform 1 0 2836 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6260
timestamp 1680363874
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1680363874
transform 1 0 2836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1680363874
transform 1 0 2788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1680363874
transform 1 0 2740 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1680363874
transform 1 0 2764 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5836
timestamp 1680363874
transform 1 0 2724 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6417
timestamp 1680363874
transform 1 0 2740 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1680363874
transform 1 0 2756 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5837
timestamp 1680363874
transform 1 0 2764 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1680363874
transform 1 0 2676 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1680363874
transform 1 0 2740 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1680363874
transform 1 0 2652 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6262
timestamp 1680363874
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1680363874
transform 1 0 2820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1680363874
transform 1 0 2844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1680363874
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1680363874
transform 1 0 2868 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5838
timestamp 1680363874
transform 1 0 2868 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1680363874
transform 1 0 2860 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6264
timestamp 1680363874
transform 1 0 2908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1680363874
transform 1 0 2916 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5809
timestamp 1680363874
transform 1 0 2916 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1680363874
transform 1 0 2908 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1680363874
transform 1 0 2948 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6265
timestamp 1680363874
transform 1 0 2940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1680363874
transform 1 0 2948 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5858
timestamp 1680363874
transform 1 0 2948 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6266
timestamp 1680363874
transform 1 0 2980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1680363874
transform 1 0 3004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1680363874
transform 1 0 3012 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1680363874
transform 1 0 2988 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5810
timestamp 1680363874
transform 1 0 2988 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1680363874
transform 1 0 3020 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6362
timestamp 1680363874
transform 1 0 3028 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5811
timestamp 1680363874
transform 1 0 3028 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6269
timestamp 1680363874
transform 1 0 3052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1680363874
transform 1 0 3068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1680363874
transform 1 0 3060 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5859
timestamp 1680363874
transform 1 0 3060 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6271
timestamp 1680363874
transform 1 0 3092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1680363874
transform 1 0 3100 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5860
timestamp 1680363874
transform 1 0 3100 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1680363874
transform 1 0 3132 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6272
timestamp 1680363874
transform 1 0 3148 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5695
timestamp 1680363874
transform 1 0 3188 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1680363874
transform 1 0 3260 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6273
timestamp 1680363874
transform 1 0 3188 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5749
timestamp 1680363874
transform 1 0 3236 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1680363874
transform 1 0 3228 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6365
timestamp 1680363874
transform 1 0 3236 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5776
timestamp 1680363874
transform 1 0 3260 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6366
timestamp 1680363874
transform 1 0 3268 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1680363874
transform 1 0 3276 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5812
timestamp 1680363874
transform 1 0 3236 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1680363874
transform 1 0 3276 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1680363874
transform 1 0 3356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1680363874
transform 1 0 3348 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6274
timestamp 1680363874
transform 1 0 3340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1680363874
transform 1 0 3348 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5723
timestamp 1680363874
transform 1 0 3372 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6368
timestamp 1680363874
transform 1 0 3356 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5777
timestamp 1680363874
transform 1 0 3364 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6369
timestamp 1680363874
transform 1 0 3372 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5814
timestamp 1680363874
transform 1 0 3372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1680363874
transform 1 0 3396 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1680363874
transform 1 0 3388 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1680363874
transform 1 0 3420 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6276
timestamp 1680363874
transform 1 0 3428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1680363874
transform 1 0 3436 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5815
timestamp 1680363874
transform 1 0 3428 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1680363874
transform 1 0 3452 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1680363874
transform 1 0 3468 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1680363874
transform 1 0 3476 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6277
timestamp 1680363874
transform 1 0 3484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1680363874
transform 1 0 3500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1680363874
transform 1 0 3508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1680363874
transform 1 0 3476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1680363874
transform 1 0 3492 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5778
timestamp 1680363874
transform 1 0 3500 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6373
timestamp 1680363874
transform 1 0 3508 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5816
timestamp 1680363874
transform 1 0 3492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1680363874
transform 1 0 3476 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1680363874
transform 1 0 3500 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1680363874
transform 1 0 3604 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6374
timestamp 1680363874
transform 1 0 3612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1680363874
transform 1 0 3732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1680363874
transform 1 0 3684 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5874
timestamp 1680363874
transform 1 0 3676 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1680363874
transform 1 0 3732 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1680363874
transform 1 0 3788 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6281
timestamp 1680363874
transform 1 0 3804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1680363874
transform 1 0 3812 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5817
timestamp 1680363874
transform 1 0 3804 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1680363874
transform 1 0 3796 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6377
timestamp 1680363874
transform 1 0 3828 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5842
timestamp 1680363874
transform 1 0 3828 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1680363874
transform 1 0 3852 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1680363874
transform 1 0 3884 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6282
timestamp 1680363874
transform 1 0 3860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1680363874
transform 1 0 3884 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5843
timestamp 1680363874
transform 1 0 3844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1680363874
transform 1 0 3892 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6378
timestamp 1680363874
transform 1 0 3876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1680363874
transform 1 0 3892 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5818
timestamp 1680363874
transform 1 0 3876 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1680363874
transform 1 0 3892 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1680363874
transform 1 0 3884 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1680363874
transform 1 0 3916 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6284
timestamp 1680363874
transform 1 0 3908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1680363874
transform 1 0 3908 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5727
timestamp 1680363874
transform 1 0 3956 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6285
timestamp 1680363874
transform 1 0 3940 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5755
timestamp 1680363874
transform 1 0 3948 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6286
timestamp 1680363874
transform 1 0 3956 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5756
timestamp 1680363874
transform 1 0 3964 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6287
timestamp 1680363874
transform 1 0 3972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1680363874
transform 1 0 3948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1680363874
transform 1 0 3964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1680363874
transform 1 0 3980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5820
timestamp 1680363874
transform 1 0 3940 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1680363874
transform 1 0 3964 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1680363874
transform 1 0 3980 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1680363874
transform 1 0 3956 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6384
timestamp 1680363874
transform 1 0 3996 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5700
timestamp 1680363874
transform 1 0 4044 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6288
timestamp 1680363874
transform 1 0 4044 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5701
timestamp 1680363874
transform 1 0 4108 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1680363874
transform 1 0 4092 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6289
timestamp 1680363874
transform 1 0 4084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1680363874
transform 1 0 4092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1680363874
transform 1 0 4116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1680363874
transform 1 0 4084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1680363874
transform 1 0 4100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1680363874
transform 1 0 4116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1680363874
transform 1 0 4076 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5822
timestamp 1680363874
transform 1 0 4116 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1680363874
transform 1 0 4148 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1680363874
transform 1 0 4140 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6292
timestamp 1680363874
transform 1 0 4140 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5780
timestamp 1680363874
transform 1 0 4132 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1680363874
transform 1 0 4172 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6293
timestamp 1680363874
transform 1 0 4180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1680363874
transform 1 0 4156 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5781
timestamp 1680363874
transform 1 0 4164 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6389
timestamp 1680363874
transform 1 0 4172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1680363874
transform 1 0 4188 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5823
timestamp 1680363874
transform 1 0 4188 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1680363874
transform 1 0 4204 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1680363874
transform 1 0 4204 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1680363874
transform 1 0 4220 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1680363874
transform 1 0 4220 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1680363874
transform 1 0 4228 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6294
timestamp 1680363874
transform 1 0 4236 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5824
timestamp 1680363874
transform 1 0 4236 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1680363874
transform 1 0 4260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1680363874
transform 1 0 4268 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6295
timestamp 1680363874
transform 1 0 4260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1680363874
transform 1 0 4252 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5783
timestamp 1680363874
transform 1 0 4260 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1680363874
transform 1 0 4284 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6296
timestamp 1680363874
transform 1 0 4300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1680363874
transform 1 0 4276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1680363874
transform 1 0 4292 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5825
timestamp 1680363874
transform 1 0 4292 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6394
timestamp 1680363874
transform 1 0 4316 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5845
timestamp 1680363874
transform 1 0 4316 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6395
timestamp 1680363874
transform 1 0 4364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1680363874
transform 1 0 4388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1680363874
transform 1 0 4396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1680363874
transform 1 0 4420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1680363874
transform 1 0 4380 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5846
timestamp 1680363874
transform 1 0 4380 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1680363874
transform 1 0 4396 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6397
timestamp 1680363874
transform 1 0 4404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1680363874
transform 1 0 4420 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5847
timestamp 1680363874
transform 1 0 4420 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1680363874
transform 1 0 4444 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6300
timestamp 1680363874
transform 1 0 4444 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5785
timestamp 1680363874
transform 1 0 4444 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1680363874
transform 1 0 4468 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6301
timestamp 1680363874
transform 1 0 4468 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5734
timestamp 1680363874
transform 1 0 4484 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1680363874
transform 1 0 4492 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1680363874
transform 1 0 4580 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6302
timestamp 1680363874
transform 1 0 4564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1680363874
transform 1 0 4580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1680363874
transform 1 0 4556 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5876
timestamp 1680363874
transform 1 0 4548 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1680363874
transform 1 0 4564 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6400
timestamp 1680363874
transform 1 0 4572 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5736
timestamp 1680363874
transform 1 0 4604 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1680363874
transform 1 0 4596 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6401
timestamp 1680363874
transform 1 0 4620 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1680363874
transform 1 0 4644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1680363874
transform 1 0 4660 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1680363874
transform 1 0 4636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1680363874
transform 1 0 4652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1680363874
transform 1 0 4668 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5849
timestamp 1680363874
transform 1 0 4628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1680363874
transform 1 0 4652 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1680363874
transform 1 0 4668 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1680363874
transform 1 0 4692 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6306
timestamp 1680363874
transform 1 0 4716 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5827
timestamp 1680363874
transform 1 0 4716 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6405
timestamp 1680363874
transform 1 0 4740 0 1 1725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_60
timestamp 1680363874
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_6967
timestamp 1680363874
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6973
timestamp 1680363874
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_425
timestamp 1680363874
transform -1 0 104 0 -1 1770
box -9 -3 26 105
use FILL  FILL_6974
timestamp 1680363874
transform 1 0 104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6975
timestamp 1680363874
transform 1 0 112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6976
timestamp 1680363874
transform 1 0 120 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_50
timestamp 1680363874
transform 1 0 128 0 -1 1770
box -8 -3 40 105
use FILL  FILL_6977
timestamp 1680363874
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6979
timestamp 1680363874
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6981
timestamp 1680363874
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6983
timestamp 1680363874
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6986
timestamp 1680363874
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6987
timestamp 1680363874
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6988
timestamp 1680363874
transform 1 0 208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6989
timestamp 1680363874
transform 1 0 216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6991
timestamp 1680363874
transform 1 0 224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_6993
timestamp 1680363874
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7003
timestamp 1680363874
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7004
timestamp 1680363874
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7005
timestamp 1680363874
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7006
timestamp 1680363874
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_365
timestamp 1680363874
transform 1 0 272 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_366
timestamp 1680363874
transform 1 0 368 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7007
timestamp 1680363874
transform 1 0 464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7009
timestamp 1680363874
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_367
timestamp 1680363874
transform 1 0 480 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7023
timestamp 1680363874
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7025
timestamp 1680363874
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7027
timestamp 1680363874
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7029
timestamp 1680363874
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7037
timestamp 1680363874
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7038
timestamp 1680363874
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FAX1  FAX1_19
timestamp 1680363874
transform 1 0 624 0 -1 1770
box -5 -3 126 105
use FILL  FILL_7039
timestamp 1680363874
transform 1 0 744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7040
timestamp 1680363874
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7041
timestamp 1680363874
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7042
timestamp 1680363874
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7043
timestamp 1680363874
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7044
timestamp 1680363874
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_369
timestamp 1680363874
transform 1 0 792 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7058
timestamp 1680363874
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7065
timestamp 1680363874
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7066
timestamp 1680363874
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7067
timestamp 1680363874
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7068
timestamp 1680363874
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7069
timestamp 1680363874
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7070
timestamp 1680363874
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7071
timestamp 1680363874
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_371
timestamp 1680363874
transform 1 0 952 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7072
timestamp 1680363874
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7074
timestamp 1680363874
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7076
timestamp 1680363874
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7078
timestamp 1680363874
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7080
timestamp 1680363874
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7082
timestamp 1680363874
transform 1 0 1088 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_285
timestamp 1680363874
transform 1 0 1096 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7089
timestamp 1680363874
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7090
timestamp 1680363874
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7091
timestamp 1680363874
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7092
timestamp 1680363874
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7093
timestamp 1680363874
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7094
timestamp 1680363874
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7096
timestamp 1680363874
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7098
timestamp 1680363874
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7100
timestamp 1680363874
transform 1 0 1200 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_287
timestamp 1680363874
transform 1 0 1208 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7106
timestamp 1680363874
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7107
timestamp 1680363874
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7108
timestamp 1680363874
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7109
timestamp 1680363874
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7110
timestamp 1680363874
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7112
timestamp 1680363874
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7124
timestamp 1680363874
transform 1 0 1296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7125
timestamp 1680363874
transform 1 0 1304 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_372
timestamp 1680363874
transform -1 0 1408 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7126
timestamp 1680363874
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_373
timestamp 1680363874
transform 1 0 1416 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7136
timestamp 1680363874
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7138
timestamp 1680363874
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7139
timestamp 1680363874
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7140
timestamp 1680363874
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_288
timestamp 1680363874
transform 1 0 1544 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7141
timestamp 1680363874
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7142
timestamp 1680363874
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7143
timestamp 1680363874
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7144
timestamp 1680363874
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7145
timestamp 1680363874
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7147
timestamp 1680363874
transform 1 0 1624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7149
timestamp 1680363874
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7151
timestamp 1680363874
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_431
timestamp 1680363874
transform 1 0 1648 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7153
timestamp 1680363874
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7155
timestamp 1680363874
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7157
timestamp 1680363874
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7159
timestamp 1680363874
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7161
timestamp 1680363874
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7172
timestamp 1680363874
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7173
timestamp 1680363874
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_375
timestamp 1680363874
transform -1 0 1816 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7174
timestamp 1680363874
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7176
timestamp 1680363874
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5878
timestamp 1680363874
transform 1 0 1876 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1680363874
transform 1 0 1916 0 1 1675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_376
timestamp 1680363874
transform 1 0 1832 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7185
timestamp 1680363874
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7186
timestamp 1680363874
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7187
timestamp 1680363874
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7188
timestamp 1680363874
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7189
timestamp 1680363874
transform 1 0 1960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7190
timestamp 1680363874
transform 1 0 1968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7192
timestamp 1680363874
transform 1 0 1976 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_377
timestamp 1680363874
transform 1 0 1984 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_432
timestamp 1680363874
transform 1 0 2080 0 -1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_378
timestamp 1680363874
transform 1 0 2096 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7209
timestamp 1680363874
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7210
timestamp 1680363874
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_433
timestamp 1680363874
transform 1 0 2208 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7211
timestamp 1680363874
transform 1 0 2224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7213
timestamp 1680363874
transform 1 0 2232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7215
timestamp 1680363874
transform 1 0 2240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7217
timestamp 1680363874
transform 1 0 2248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7227
timestamp 1680363874
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7228
timestamp 1680363874
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5880
timestamp 1680363874
transform 1 0 2284 0 1 1675
box -3 -3 3 3
use AOI22X1  AOI22X1_229
timestamp 1680363874
transform -1 0 2312 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7229
timestamp 1680363874
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7230
timestamp 1680363874
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7231
timestamp 1680363874
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7232
timestamp 1680363874
transform 1 0 2336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7233
timestamp 1680363874
transform 1 0 2344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7234
timestamp 1680363874
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7235
timestamp 1680363874
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7236
timestamp 1680363874
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_52
timestamp 1680363874
transform 1 0 2376 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7237
timestamp 1680363874
transform 1 0 2408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7238
timestamp 1680363874
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7239
timestamp 1680363874
transform 1 0 2424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7240
timestamp 1680363874
transform 1 0 2432 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_380
timestamp 1680363874
transform 1 0 2440 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7241
timestamp 1680363874
transform 1 0 2536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7256
timestamp 1680363874
transform 1 0 2544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7257
timestamp 1680363874
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7258
timestamp 1680363874
transform 1 0 2560 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_52
timestamp 1680363874
transform 1 0 2568 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7259
timestamp 1680363874
transform 1 0 2592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7260
timestamp 1680363874
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_53
timestamp 1680363874
transform 1 0 2608 0 -1 1770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_382
timestamp 1680363874
transform 1 0 2640 0 -1 1770
box -8 -3 104 105
use NAND3X1  NAND3X1_54
timestamp 1680363874
transform 1 0 2736 0 -1 1770
box -8 -3 40 105
use BUFX2  BUFX2_53
timestamp 1680363874
transform -1 0 2792 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_54
timestamp 1680363874
transform 1 0 2792 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_55
timestamp 1680363874
transform 1 0 2816 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_56
timestamp 1680363874
transform 1 0 2840 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7261
timestamp 1680363874
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7262
timestamp 1680363874
transform 1 0 2872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7263
timestamp 1680363874
transform 1 0 2880 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_57
timestamp 1680363874
transform 1 0 2888 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7264
timestamp 1680363874
transform 1 0 2912 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_58
timestamp 1680363874
transform 1 0 2920 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7265
timestamp 1680363874
transform 1 0 2944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7266
timestamp 1680363874
transform 1 0 2952 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_60
timestamp 1680363874
transform 1 0 2960 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_61
timestamp 1680363874
transform 1 0 2984 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_62
timestamp 1680363874
transform -1 0 3032 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_63
timestamp 1680363874
transform 1 0 3032 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7277
timestamp 1680363874
transform 1 0 3056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7278
timestamp 1680363874
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5881
timestamp 1680363874
transform 1 0 3100 0 1 1675
box -3 -3 3 3
use BUFX2  BUFX2_64
timestamp 1680363874
transform 1 0 3072 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7279
timestamp 1680363874
transform 1 0 3096 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_66
timestamp 1680363874
transform 1 0 3104 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7283
timestamp 1680363874
transform 1 0 3128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7284
timestamp 1680363874
transform 1 0 3136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7285
timestamp 1680363874
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7287
timestamp 1680363874
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7297
timestamp 1680363874
transform 1 0 3160 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5882
timestamp 1680363874
transform 1 0 3180 0 1 1675
box -3 -3 3 3
use FILL  FILL_7298
timestamp 1680363874
transform 1 0 3168 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_383
timestamp 1680363874
transform 1 0 3176 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7299
timestamp 1680363874
transform 1 0 3272 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_439
timestamp 1680363874
transform -1 0 3296 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7300
timestamp 1680363874
transform 1 0 3296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7301
timestamp 1680363874
transform 1 0 3304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7302
timestamp 1680363874
transform 1 0 3312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7304
timestamp 1680363874
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7306
timestamp 1680363874
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7308
timestamp 1680363874
transform 1 0 3336 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_43
timestamp 1680363874
transform 1 0 3344 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7311
timestamp 1680363874
transform 1 0 3376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7313
timestamp 1680363874
transform 1 0 3384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7315
timestamp 1680363874
transform 1 0 3392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7319
timestamp 1680363874
transform 1 0 3400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7320
timestamp 1680363874
transform 1 0 3408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7321
timestamp 1680363874
transform 1 0 3416 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_440
timestamp 1680363874
transform 1 0 3424 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7322
timestamp 1680363874
transform 1 0 3440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7323
timestamp 1680363874
transform 1 0 3448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7324
timestamp 1680363874
transform 1 0 3456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7325
timestamp 1680363874
transform 1 0 3464 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_232
timestamp 1680363874
transform -1 0 3512 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7326
timestamp 1680363874
transform 1 0 3512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7328
timestamp 1680363874
transform 1 0 3520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7330
timestamp 1680363874
transform 1 0 3528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7332
timestamp 1680363874
transform 1 0 3536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7334
timestamp 1680363874
transform 1 0 3544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7336
timestamp 1680363874
transform 1 0 3552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7337
timestamp 1680363874
transform 1 0 3560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7338
timestamp 1680363874
transform 1 0 3568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7339
timestamp 1680363874
transform 1 0 3576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7340
timestamp 1680363874
transform 1 0 3584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7341
timestamp 1680363874
transform 1 0 3592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7343
timestamp 1680363874
transform 1 0 3600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7345
timestamp 1680363874
transform 1 0 3608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7347
timestamp 1680363874
transform 1 0 3616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7349
timestamp 1680363874
transform 1 0 3624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7351
timestamp 1680363874
transform 1 0 3632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7359
timestamp 1680363874
transform 1 0 3640 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_385
timestamp 1680363874
transform -1 0 3744 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7360
timestamp 1680363874
transform 1 0 3744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7361
timestamp 1680363874
transform 1 0 3752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7362
timestamp 1680363874
transform 1 0 3760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7363
timestamp 1680363874
transform 1 0 3768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7368
timestamp 1680363874
transform 1 0 3776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7369
timestamp 1680363874
transform 1 0 3784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7370
timestamp 1680363874
transform 1 0 3792 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_442
timestamp 1680363874
transform 1 0 3800 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7371
timestamp 1680363874
transform 1 0 3816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7372
timestamp 1680363874
transform 1 0 3824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7373
timestamp 1680363874
transform 1 0 3832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7374
timestamp 1680363874
transform 1 0 3840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7375
timestamp 1680363874
transform 1 0 3848 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_234
timestamp 1680363874
transform -1 0 3896 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7376
timestamp 1680363874
transform 1 0 3896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7384
timestamp 1680363874
transform 1 0 3904 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5883
timestamp 1680363874
transform 1 0 3924 0 1 1675
box -3 -3 3 3
use FILL  FILL_7385
timestamp 1680363874
transform 1 0 3912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7386
timestamp 1680363874
transform 1 0 3920 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_443
timestamp 1680363874
transform -1 0 3944 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_235
timestamp 1680363874
transform 1 0 3944 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7387
timestamp 1680363874
transform 1 0 3984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7388
timestamp 1680363874
transform 1 0 3992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7389
timestamp 1680363874
transform 1 0 4000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7390
timestamp 1680363874
transform 1 0 4008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7391
timestamp 1680363874
transform 1 0 4016 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_71
timestamp 1680363874
transform 1 0 4024 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7392
timestamp 1680363874
transform 1 0 4048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7394
timestamp 1680363874
transform 1 0 4056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7396
timestamp 1680363874
transform 1 0 4064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7399
timestamp 1680363874
transform 1 0 4072 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_236
timestamp 1680363874
transform 1 0 4080 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7400
timestamp 1680363874
transform 1 0 4120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7401
timestamp 1680363874
transform 1 0 4128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7402
timestamp 1680363874
transform 1 0 4136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7403
timestamp 1680363874
transform 1 0 4144 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_237
timestamp 1680363874
transform 1 0 4152 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7404
timestamp 1680363874
transform 1 0 4192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7405
timestamp 1680363874
transform 1 0 4200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7406
timestamp 1680363874
transform 1 0 4208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7407
timestamp 1680363874
transform 1 0 4216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7408
timestamp 1680363874
transform 1 0 4224 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_445
timestamp 1680363874
transform 1 0 4232 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7409
timestamp 1680363874
transform 1 0 4248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7410
timestamp 1680363874
transform 1 0 4256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7411
timestamp 1680363874
transform 1 0 4264 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_238
timestamp 1680363874
transform 1 0 4272 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7412
timestamp 1680363874
transform 1 0 4312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7414
timestamp 1680363874
transform 1 0 4320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7416
timestamp 1680363874
transform 1 0 4328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7417
timestamp 1680363874
transform 1 0 4336 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_446
timestamp 1680363874
transform -1 0 4360 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7418
timestamp 1680363874
transform 1 0 4360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7419
timestamp 1680363874
transform 1 0 4368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7420
timestamp 1680363874
transform 1 0 4376 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_239
timestamp 1680363874
transform 1 0 4384 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7421
timestamp 1680363874
transform 1 0 4424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7423
timestamp 1680363874
transform 1 0 4432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7425
timestamp 1680363874
transform 1 0 4440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7427
timestamp 1680363874
transform 1 0 4448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7429
timestamp 1680363874
transform 1 0 4456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7431
timestamp 1680363874
transform 1 0 4464 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_448
timestamp 1680363874
transform 1 0 4472 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7434
timestamp 1680363874
transform 1 0 4488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7435
timestamp 1680363874
transform 1 0 4496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7436
timestamp 1680363874
transform 1 0 4504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7437
timestamp 1680363874
transform 1 0 4512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7438
timestamp 1680363874
transform 1 0 4520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7439
timestamp 1680363874
transform 1 0 4528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7440
timestamp 1680363874
transform 1 0 4536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7441
timestamp 1680363874
transform 1 0 4544 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_240
timestamp 1680363874
transform -1 0 4592 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7442
timestamp 1680363874
transform 1 0 4592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7444
timestamp 1680363874
transform 1 0 4600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7446
timestamp 1680363874
transform 1 0 4608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7448
timestamp 1680363874
transform 1 0 4616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7450
timestamp 1680363874
transform 1 0 4624 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_242
timestamp 1680363874
transform 1 0 4632 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7452
timestamp 1680363874
transform 1 0 4672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7454
timestamp 1680363874
transform 1 0 4680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7455
timestamp 1680363874
transform 1 0 4688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7456
timestamp 1680363874
transform 1 0 4696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7457
timestamp 1680363874
transform 1 0 4704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7458
timestamp 1680363874
transform 1 0 4712 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_450
timestamp 1680363874
transform 1 0 4720 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7459
timestamp 1680363874
transform 1 0 4736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7460
timestamp 1680363874
transform 1 0 4744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7461
timestamp 1680363874
transform 1 0 4752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7462
timestamp 1680363874
transform 1 0 4760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7463
timestamp 1680363874
transform 1 0 4768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7464
timestamp 1680363874
transform 1 0 4776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7465
timestamp 1680363874
transform 1 0 4784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7466
timestamp 1680363874
transform 1 0 4792 0 -1 1770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_61
timestamp 1680363874
transform 1 0 4851 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_6433
timestamp 1680363874
transform 1 0 116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1680363874
transform 1 0 108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1680363874
transform 1 0 100 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5945
timestamp 1680363874
transform 1 0 140 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6423
timestamp 1680363874
transform 1 0 164 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1680363874
transform 1 0 196 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5946
timestamp 1680363874
transform 1 0 220 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6434
timestamp 1680363874
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1680363874
transform 1 0 228 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5913
timestamp 1680363874
transform 1 0 412 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1680363874
transform 1 0 340 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1680363874
transform 1 0 356 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6435
timestamp 1680363874
transform 1 0 316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1680363874
transform 1 0 356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1680363874
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1680363874
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5975
timestamp 1680363874
transform 1 0 388 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6538
timestamp 1680363874
transform 1 0 268 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1680363874
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6016
timestamp 1680363874
transform 1 0 284 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1680363874
transform 1 0 356 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6626
timestamp 1680363874
transform 1 0 460 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_6018
timestamp 1680363874
transform 1 0 468 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6627
timestamp 1680363874
transform 1 0 476 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5914
timestamp 1680363874
transform 1 0 524 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5915
timestamp 1680363874
transform 1 0 580 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5949
timestamp 1680363874
transform 1 0 596 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1680363874
transform 1 0 564 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1680363874
transform 1 0 580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6439
timestamp 1680363874
transform 1 0 596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1680363874
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5978
timestamp 1680363874
transform 1 0 612 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5988
timestamp 1680363874
transform 1 0 596 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6540
timestamp 1680363874
transform 1 0 612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1680363874
transform 1 0 508 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1680363874
transform 1 0 628 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5916
timestamp 1680363874
transform 1 0 660 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1680363874
transform 1 0 740 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1680363874
transform 1 0 652 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6542
timestamp 1680363874
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1680363874
transform 1 0 756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1680363874
transform 1 0 772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1680363874
transform 1 0 668 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1680363874
transform 1 0 788 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5951
timestamp 1680363874
transform 1 0 820 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6443
timestamp 1680363874
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1680363874
transform 1 0 860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1680363874
transform 1 0 884 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5989
timestamp 1680363874
transform 1 0 900 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6633
timestamp 1680363874
transform 1 0 900 0 1 1585
box -2 -2 2 2
use M3_M2  M3_M2_5952
timestamp 1680363874
transform 1 0 916 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6545
timestamp 1680363874
transform 1 0 916 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6019
timestamp 1680363874
transform 1 0 916 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1680363874
transform 1 0 988 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1680363874
transform 1 0 980 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6445
timestamp 1680363874
transform 1 0 980 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5918
timestamp 1680363874
transform 1 0 1020 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1680363874
transform 1 0 1036 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6446
timestamp 1680363874
transform 1 0 1036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1680363874
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5990
timestamp 1680363874
transform 1 0 1036 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1680363874
transform 1 0 1116 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6447
timestamp 1680363874
transform 1 0 1116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1680363874
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6043
timestamp 1680363874
transform 1 0 1140 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1680363874
transform 1 0 1164 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6448
timestamp 1680363874
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5991
timestamp 1680363874
transform 1 0 1164 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6419
timestamp 1680363874
transform 1 0 1196 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1680363874
transform 1 0 1172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1680363874
transform 1 0 1188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1680363874
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5992
timestamp 1680363874
transform 1 0 1212 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6550
timestamp 1680363874
transform 1 0 1284 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5979
timestamp 1680363874
transform 1 0 1308 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6551
timestamp 1680363874
transform 1 0 1308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1680363874
transform 1 0 1324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1680363874
transform 1 0 1332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1680363874
transform 1 0 1348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1680363874
transform 1 0 1364 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5980
timestamp 1680363874
transform 1 0 1372 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6453
timestamp 1680363874
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1680363874
transform 1 0 1340 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5993
timestamp 1680363874
transform 1 0 1348 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6554
timestamp 1680363874
transform 1 0 1356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1680363874
transform 1 0 1372 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6020
timestamp 1680363874
transform 1 0 1356 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1680363874
transform 1 0 1372 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6454
timestamp 1680363874
transform 1 0 1436 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5994
timestamp 1680363874
transform 1 0 1444 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6556
timestamp 1680363874
transform 1 0 1484 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6021
timestamp 1680363874
transform 1 0 1436 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6455
timestamp 1680363874
transform 1 0 1500 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5995
timestamp 1680363874
transform 1 0 1500 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6557
timestamp 1680363874
transform 1 0 1508 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6045
timestamp 1680363874
transform 1 0 1508 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6558
timestamp 1680363874
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5922
timestamp 1680363874
transform 1 0 1556 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6456
timestamp 1680363874
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1680363874
transform 1 0 1564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1680363874
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6022
timestamp 1680363874
transform 1 0 1580 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1680363874
transform 1 0 1588 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6560
timestamp 1680363874
transform 1 0 1604 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5901
timestamp 1680363874
transform 1 0 1652 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6458
timestamp 1680363874
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1680363874
transform 1 0 1668 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5981
timestamp 1680363874
transform 1 0 1676 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6460
timestamp 1680363874
transform 1 0 1684 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1680363874
transform 1 0 1644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1680363874
transform 1 0 1660 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5996
timestamp 1680363874
transform 1 0 1668 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6563
timestamp 1680363874
transform 1 0 1676 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5997
timestamp 1680363874
transform 1 0 1684 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1680363874
transform 1 0 1676 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1680363874
transform 1 0 1748 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6461
timestamp 1680363874
transform 1 0 1748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1680363874
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6024
timestamp 1680363874
transform 1 0 1756 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5902
timestamp 1680363874
transform 1 0 1780 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6462
timestamp 1680363874
transform 1 0 1796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1680363874
transform 1 0 1812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1680363874
transform 1 0 1788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1680363874
transform 1 0 1804 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5998
timestamp 1680363874
transform 1 0 1812 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6567
timestamp 1680363874
transform 1 0 1820 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6047
timestamp 1680363874
transform 1 0 1820 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5903
timestamp 1680363874
transform 1 0 1836 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6464
timestamp 1680363874
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1680363874
transform 1 0 1844 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6025
timestamp 1680363874
transform 1 0 1836 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6569
timestamp 1680363874
transform 1 0 1860 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5924
timestamp 1680363874
transform 1 0 1900 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6465
timestamp 1680363874
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1680363874
transform 1 0 1916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1680363874
transform 1 0 1892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1680363874
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5999
timestamp 1680363874
transform 1 0 1916 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1680363874
transform 1 0 1924 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1680363874
transform 1 0 1948 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6467
timestamp 1680363874
transform 1 0 1948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1680363874
transform 1 0 1940 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5904
timestamp 1680363874
transform 1 0 1972 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6468
timestamp 1680363874
transform 1 0 1972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1680363874
transform 1 0 1980 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1680363874
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5905
timestamp 1680363874
transform 1 0 2052 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6470
timestamp 1680363874
transform 1 0 2052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1680363874
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1680363874
transform 1 0 2028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1680363874
transform 1 0 2044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1680363874
transform 1 0 2052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1680363874
transform 1 0 2068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1680363874
transform 1 0 2124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1680363874
transform 1 0 2116 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6000
timestamp 1680363874
transform 1 0 2124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5906
timestamp 1680363874
transform 1 0 2140 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6472
timestamp 1680363874
transform 1 0 2140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1680363874
transform 1 0 2132 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6048
timestamp 1680363874
transform 1 0 2132 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6473
timestamp 1680363874
transform 1 0 2164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1680363874
transform 1 0 2156 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5926
timestamp 1680363874
transform 1 0 2180 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6474
timestamp 1680363874
transform 1 0 2204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1680363874
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6027
timestamp 1680363874
transform 1 0 2172 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1680363874
transform 1 0 2188 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6583
timestamp 1680363874
transform 1 0 2196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1680363874
transform 1 0 2212 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6049
timestamp 1680363874
transform 1 0 2180 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1680363874
transform 1 0 2228 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1680363874
transform 1 0 2220 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6050
timestamp 1680363874
transform 1 0 2212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1680363874
transform 1 0 2268 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1680363874
transform 1 0 2292 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1680363874
transform 1 0 2244 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6475
timestamp 1680363874
transform 1 0 2276 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1680363874
transform 1 0 2332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1680363874
transform 1 0 2252 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6029
timestamp 1680363874
transform 1 0 2252 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1680363874
transform 1 0 2276 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1680363874
transform 1 0 2356 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6477
timestamp 1680363874
transform 1 0 2380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1680363874
transform 1 0 2356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6003
timestamp 1680363874
transform 1 0 2428 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1680363874
transform 1 0 2420 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1680363874
transform 1 0 2452 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6478
timestamp 1680363874
transform 1 0 2444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1680363874
transform 1 0 2452 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6031
timestamp 1680363874
transform 1 0 2444 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1680363874
transform 1 0 2468 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6479
timestamp 1680363874
transform 1 0 2492 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6005
timestamp 1680363874
transform 1 0 2484 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6588
timestamp 1680363874
transform 1 0 2492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1680363874
transform 1 0 2484 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_6032
timestamp 1680363874
transform 1 0 2492 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1680363874
transform 1 0 2492 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6480
timestamp 1680363874
transform 1 0 2516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1680363874
transform 1 0 2532 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6006
timestamp 1680363874
transform 1 0 2516 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1680363874
transform 1 0 2532 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6424
timestamp 1680363874
transform 1 0 2564 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_6007
timestamp 1680363874
transform 1 0 2556 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6425
timestamp 1680363874
transform 1 0 2588 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1680363874
transform 1 0 2588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1680363874
transform 1 0 2628 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1680363874
transform 1 0 2612 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1680363874
transform 1 0 2620 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6008
timestamp 1680363874
transform 1 0 2628 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1680363874
transform 1 0 2676 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6421
timestamp 1680363874
transform 1 0 2684 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1680363874
transform 1 0 2676 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1680363874
transform 1 0 2692 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5954
timestamp 1680363874
transform 1 0 2700 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6484
timestamp 1680363874
transform 1 0 2692 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5884
timestamp 1680363874
transform 1 0 2732 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5928
timestamp 1680363874
transform 1 0 2748 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6422
timestamp 1680363874
transform 1 0 2756 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5955
timestamp 1680363874
transform 1 0 2740 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6429
timestamp 1680363874
transform 1 0 2748 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1680363874
transform 1 0 2756 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5956
timestamp 1680363874
transform 1 0 2764 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6485
timestamp 1680363874
transform 1 0 2764 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5929
timestamp 1680363874
transform 1 0 2788 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6486
timestamp 1680363874
transform 1 0 2788 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5885
timestamp 1680363874
transform 1 0 2812 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1680363874
transform 1 0 2812 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6431
timestamp 1680363874
transform 1 0 2812 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5957
timestamp 1680363874
transform 1 0 2820 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6487
timestamp 1680363874
transform 1 0 2820 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5886
timestamp 1680363874
transform 1 0 2844 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1680363874
transform 1 0 2860 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1680363874
transform 1 0 2852 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6488
timestamp 1680363874
transform 1 0 2852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1680363874
transform 1 0 2844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1680363874
transform 1 0 2876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1680363874
transform 1 0 2884 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5895
timestamp 1680363874
transform 1 0 2916 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1680363874
transform 1 0 2948 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1680363874
transform 1 0 2980 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6490
timestamp 1680363874
transform 1 0 2948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1680363874
transform 1 0 2972 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6033
timestamp 1680363874
transform 1 0 2972 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6491
timestamp 1680363874
transform 1 0 2988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1680363874
transform 1 0 3044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1680363874
transform 1 0 3076 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6034
timestamp 1680363874
transform 1 0 3076 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6634
timestamp 1680363874
transform 1 0 3092 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1680363874
transform 1 0 3108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1680363874
transform 1 0 3100 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5959
timestamp 1680363874
transform 1 0 3132 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6494
timestamp 1680363874
transform 1 0 3124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1680363874
transform 1 0 3132 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6009
timestamp 1680363874
transform 1 0 3124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1680363874
transform 1 0 3116 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1680363874
transform 1 0 3164 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6496
timestamp 1680363874
transform 1 0 3164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1680363874
transform 1 0 3156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1680363874
transform 1 0 3180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1680363874
transform 1 0 3252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1680363874
transform 1 0 3204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5887
timestamp 1680363874
transform 1 0 3316 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1680363874
transform 1 0 3316 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1680363874
transform 1 0 3340 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1680363874
transform 1 0 3380 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1680363874
transform 1 0 3348 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1680363874
transform 1 0 3372 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6498
timestamp 1680363874
transform 1 0 3332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1680363874
transform 1 0 3340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1680363874
transform 1 0 3356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1680363874
transform 1 0 3340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1680363874
transform 1 0 3348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1680363874
transform 1 0 3364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1680363874
transform 1 0 3372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1680363874
transform 1 0 3388 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5963
timestamp 1680363874
transform 1 0 3404 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6501
timestamp 1680363874
transform 1 0 3404 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6010
timestamp 1680363874
transform 1 0 3436 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6631
timestamp 1680363874
transform 1 0 3428 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5964
timestamp 1680363874
transform 1 0 3476 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6502
timestamp 1680363874
transform 1 0 3476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1680363874
transform 1 0 3532 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6054
timestamp 1680363874
transform 1 0 3548 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1680363874
transform 1 0 3612 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6503
timestamp 1680363874
transform 1 0 3572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1680363874
transform 1 0 3580 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1680363874
transform 1 0 3596 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5982
timestamp 1680363874
transform 1 0 3604 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6506
timestamp 1680363874
transform 1 0 3612 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6011
timestamp 1680363874
transform 1 0 3580 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6603
timestamp 1680363874
transform 1 0 3612 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6055
timestamp 1680363874
transform 1 0 3612 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1680363874
transform 1 0 3660 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1680363874
transform 1 0 3732 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1680363874
transform 1 0 3692 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6507
timestamp 1680363874
transform 1 0 3740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1680363874
transform 1 0 3692 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6036
timestamp 1680363874
transform 1 0 3716 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1680363874
transform 1 0 3708 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6508
timestamp 1680363874
transform 1 0 3780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1680363874
transform 1 0 3788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1680363874
transform 1 0 3796 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6057
timestamp 1680363874
transform 1 0 3788 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6510
timestamp 1680363874
transform 1 0 3828 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5983
timestamp 1680363874
transform 1 0 3836 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1680363874
transform 1 0 3868 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1680363874
transform 1 0 3852 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1680363874
transform 1 0 3868 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1680363874
transform 1 0 3852 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6511
timestamp 1680363874
transform 1 0 3844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1680363874
transform 1 0 3836 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6012
timestamp 1680363874
transform 1 0 3844 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6512
timestamp 1680363874
transform 1 0 3908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1680363874
transform 1 0 3868 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6037
timestamp 1680363874
transform 1 0 3868 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1680363874
transform 1 0 3956 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5938
timestamp 1680363874
transform 1 0 3980 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6513
timestamp 1680363874
transform 1 0 3972 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5898
timestamp 1680363874
transform 1 0 4012 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1680363874
transform 1 0 3996 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5899
timestamp 1680363874
transform 1 0 4036 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1680363874
transform 1 0 4124 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1680363874
transform 1 0 4020 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1680363874
transform 1 0 4084 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6514
timestamp 1680363874
transform 1 0 3996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1680363874
transform 1 0 4020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1680363874
transform 1 0 4084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1680363874
transform 1 0 4116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1680363874
transform 1 0 4124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1680363874
transform 1 0 4148 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5984
timestamp 1680363874
transform 1 0 4156 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6608
timestamp 1680363874
transform 1 0 4004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1680363874
transform 1 0 4020 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1680363874
transform 1 0 4036 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6013
timestamp 1680363874
transform 1 0 4116 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6611
timestamp 1680363874
transform 1 0 4124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1680363874
transform 1 0 4140 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6014
timestamp 1680363874
transform 1 0 4148 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6613
timestamp 1680363874
transform 1 0 4156 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6038
timestamp 1680363874
transform 1 0 4036 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6432
timestamp 1680363874
transform 1 0 4172 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5985
timestamp 1680363874
transform 1 0 4172 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6614
timestamp 1680363874
transform 1 0 4180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5900
timestamp 1680363874
transform 1 0 4196 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1680363874
transform 1 0 4204 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6520
timestamp 1680363874
transform 1 0 4204 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5912
timestamp 1680363874
transform 1 0 4316 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6521
timestamp 1680363874
transform 1 0 4268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1680363874
transform 1 0 4324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1680363874
transform 1 0 4244 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6039
timestamp 1680363874
transform 1 0 4292 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1680363874
transform 1 0 4244 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1680363874
transform 1 0 4428 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1680363874
transform 1 0 4396 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1680363874
transform 1 0 4436 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6523
timestamp 1680363874
transform 1 0 4396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1680363874
transform 1 0 4428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1680363874
transform 1 0 4436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1680363874
transform 1 0 4444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1680363874
transform 1 0 4348 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6059
timestamp 1680363874
transform 1 0 4348 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1680363874
transform 1 0 4500 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6527
timestamp 1680363874
transform 1 0 4492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1680363874
transform 1 0 4508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1680363874
transform 1 0 4492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1680363874
transform 1 0 4500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1680363874
transform 1 0 4516 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6040
timestamp 1680363874
transform 1 0 4516 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6620
timestamp 1680363874
transform 1 0 4532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1680363874
transform 1 0 4548 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5971
timestamp 1680363874
transform 1 0 4564 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6632
timestamp 1680363874
transform 1 0 4572 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_6060
timestamp 1680363874
transform 1 0 4572 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5972
timestamp 1680363874
transform 1 0 4612 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1680363874
transform 1 0 4636 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6530
timestamp 1680363874
transform 1 0 4612 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5986
timestamp 1680363874
transform 1 0 4620 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6531
timestamp 1680363874
transform 1 0 4628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1680363874
transform 1 0 4644 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5973
timestamp 1680363874
transform 1 0 4660 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6621
timestamp 1680363874
transform 1 0 4620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1680363874
transform 1 0 4636 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6015
timestamp 1680363874
transform 1 0 4652 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6623
timestamp 1680363874
transform 1 0 4660 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6061
timestamp 1680363874
transform 1 0 4636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1680363874
transform 1 0 4692 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6041
timestamp 1680363874
transform 1 0 4700 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1680363874
transform 1 0 4868 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1680363874
transform 1 0 4796 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6533
timestamp 1680363874
transform 1 0 4740 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5987
timestamp 1680363874
transform 1 0 4748 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6534
timestamp 1680363874
transform 1 0 4796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1680363874
transform 1 0 4716 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6042
timestamp 1680363874
transform 1 0 4716 0 1 1595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_62
timestamp 1680363874
transform 1 0 48 0 1 1570
box -10 -3 10 3
use FILL  FILL_7467
timestamp 1680363874
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_7469
timestamp 1680363874
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_7471
timestamp 1680363874
transform 1 0 88 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_82
timestamp 1680363874
transform 1 0 96 0 1 1570
box -8 -3 32 105
use FILL  FILL_7473
timestamp 1680363874
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_7475
timestamp 1680363874
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_7477
timestamp 1680363874
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7479
timestamp 1680363874
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_7481
timestamp 1680363874
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_7482
timestamp 1680363874
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_7483
timestamp 1680363874
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_7484
timestamp 1680363874
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7485
timestamp 1680363874
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7486
timestamp 1680363874
transform 1 0 192 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_145
timestamp 1680363874
transform -1 0 232 0 1 1570
box -8 -3 34 105
use FILL  FILL_7487
timestamp 1680363874
transform 1 0 232 0 1 1570
box -8 -3 16 105
use FILL  FILL_7488
timestamp 1680363874
transform 1 0 240 0 1 1570
box -8 -3 16 105
use FILL  FILL_7489
timestamp 1680363874
transform 1 0 248 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_393
timestamp 1680363874
transform 1 0 256 0 1 1570
box -8 -3 104 105
use FAX1  FAX1_20
timestamp 1680363874
transform 1 0 352 0 1 1570
box -5 -3 126 105
use FILL  FILL_7491
timestamp 1680363874
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_7492
timestamp 1680363874
transform 1 0 480 0 1 1570
box -8 -3 16 105
use FILL  FILL_7493
timestamp 1680363874
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FAX1  FAX1_21
timestamp 1680363874
transform -1 0 616 0 1 1570
box -5 -3 126 105
use FILL  FILL_7494
timestamp 1680363874
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7495
timestamp 1680363874
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7496
timestamp 1680363874
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_7497
timestamp 1680363874
transform 1 0 640 0 1 1570
box -8 -3 16 105
use FILL  FILL_7498
timestamp 1680363874
transform 1 0 648 0 1 1570
box -8 -3 16 105
use FAX1  FAX1_22
timestamp 1680363874
transform -1 0 776 0 1 1570
box -5 -3 126 105
use FILL  FILL_7499
timestamp 1680363874
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_7529
timestamp 1680363874
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7531
timestamp 1680363874
transform 1 0 792 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_394
timestamp 1680363874
transform -1 0 896 0 1 1570
box -8 -3 104 105
use FILL  FILL_7532
timestamp 1680363874
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_7533
timestamp 1680363874
transform 1 0 904 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_452
timestamp 1680363874
transform 1 0 912 0 1 1570
box -9 -3 26 105
use FILL  FILL_7534
timestamp 1680363874
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_7535
timestamp 1680363874
transform 1 0 936 0 1 1570
box -8 -3 16 105
use FILL  FILL_7536
timestamp 1680363874
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_7537
timestamp 1680363874
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7538
timestamp 1680363874
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7539
timestamp 1680363874
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_7540
timestamp 1680363874
transform 1 0 976 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_395
timestamp 1680363874
transform 1 0 984 0 1 1570
box -8 -3 104 105
use FILL  FILL_7541
timestamp 1680363874
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7560
timestamp 1680363874
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_454
timestamp 1680363874
transform 1 0 1096 0 1 1570
box -9 -3 26 105
use FILL  FILL_7562
timestamp 1680363874
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_7566
timestamp 1680363874
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_7568
timestamp 1680363874
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_7570
timestamp 1680363874
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7572
timestamp 1680363874
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_293
timestamp 1680363874
transform -1 0 1192 0 1 1570
box -8 -3 46 105
use FILL  FILL_7573
timestamp 1680363874
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_7581
timestamp 1680363874
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_7583
timestamp 1680363874
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_7585
timestamp 1680363874
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_7587
timestamp 1680363874
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use FILL  FILL_7589
timestamp 1680363874
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use FILL  FILL_7590
timestamp 1680363874
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_7591
timestamp 1680363874
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_7592
timestamp 1680363874
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_7593
timestamp 1680363874
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_7594
timestamp 1680363874
transform 1 0 1272 0 1 1570
box -8 -3 16 105
use FILL  FILL_7595
timestamp 1680363874
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_7596
timestamp 1680363874
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_7597
timestamp 1680363874
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_455
timestamp 1680363874
transform 1 0 1304 0 1 1570
box -9 -3 26 105
use FILL  FILL_7598
timestamp 1680363874
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_7599
timestamp 1680363874
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_294
timestamp 1680363874
transform 1 0 1336 0 1 1570
box -8 -3 46 105
use FILL  FILL_7601
timestamp 1680363874
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_7608
timestamp 1680363874
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_7609
timestamp 1680363874
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_398
timestamp 1680363874
transform -1 0 1496 0 1 1570
box -8 -3 104 105
use FILL  FILL_7610
timestamp 1680363874
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_7618
timestamp 1680363874
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_456
timestamp 1680363874
transform 1 0 1512 0 1 1570
box -9 -3 26 105
use FILL  FILL_7620
timestamp 1680363874
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_7624
timestamp 1680363874
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7626
timestamp 1680363874
transform 1 0 1544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7628
timestamp 1680363874
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7629
timestamp 1680363874
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7630
timestamp 1680363874
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_457
timestamp 1680363874
transform 1 0 1576 0 1 1570
box -9 -3 26 105
use FILL  FILL_7631
timestamp 1680363874
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_7633
timestamp 1680363874
transform 1 0 1600 0 1 1570
box -8 -3 16 105
use FILL  FILL_7635
timestamp 1680363874
transform 1 0 1608 0 1 1570
box -8 -3 16 105
use FILL  FILL_7637
timestamp 1680363874
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7639
timestamp 1680363874
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7641
timestamp 1680363874
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6062
timestamp 1680363874
transform 1 0 1676 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_297
timestamp 1680363874
transform 1 0 1640 0 1 1570
box -8 -3 46 105
use FILL  FILL_7643
timestamp 1680363874
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_7644
timestamp 1680363874
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_7645
timestamp 1680363874
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_7649
timestamp 1680363874
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_7651
timestamp 1680363874
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_7653
timestamp 1680363874
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_458
timestamp 1680363874
transform -1 0 1744 0 1 1570
box -9 -3 26 105
use FILL  FILL_7654
timestamp 1680363874
transform 1 0 1744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7655
timestamp 1680363874
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7658
timestamp 1680363874
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_7660
timestamp 1680363874
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_7662
timestamp 1680363874
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6063
timestamp 1680363874
transform 1 0 1820 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_298
timestamp 1680363874
transform 1 0 1784 0 1 1570
box -8 -3 46 105
use FILL  FILL_7663
timestamp 1680363874
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_7666
timestamp 1680363874
transform 1 0 1832 0 1 1570
box -8 -3 16 105
use FILL  FILL_7667
timestamp 1680363874
transform 1 0 1840 0 1 1570
box -8 -3 16 105
use FILL  FILL_7668
timestamp 1680363874
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_7669
timestamp 1680363874
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_7672
timestamp 1680363874
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6064
timestamp 1680363874
transform 1 0 1908 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_299
timestamp 1680363874
transform 1 0 1872 0 1 1570
box -8 -3 46 105
use FILL  FILL_7674
timestamp 1680363874
transform 1 0 1912 0 1 1570
box -8 -3 16 105
use FILL  FILL_7675
timestamp 1680363874
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_460
timestamp 1680363874
transform -1 0 1944 0 1 1570
box -9 -3 26 105
use FILL  FILL_7676
timestamp 1680363874
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_461
timestamp 1680363874
transform -1 0 1968 0 1 1570
box -9 -3 26 105
use FILL  FILL_7677
timestamp 1680363874
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_7678
timestamp 1680363874
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7679
timestamp 1680363874
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7683
timestamp 1680363874
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_7685
timestamp 1680363874
transform 1 0 2000 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6065
timestamp 1680363874
transform 1 0 2044 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_300
timestamp 1680363874
transform 1 0 2008 0 1 1570
box -8 -3 46 105
use FILL  FILL_7687
timestamp 1680363874
transform 1 0 2048 0 1 1570
box -8 -3 16 105
use FILL  FILL_7694
timestamp 1680363874
transform 1 0 2056 0 1 1570
box -8 -3 16 105
use FILL  FILL_7696
timestamp 1680363874
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_7697
timestamp 1680363874
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_7698
timestamp 1680363874
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7699
timestamp 1680363874
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6066
timestamp 1680363874
transform 1 0 2132 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_301
timestamp 1680363874
transform 1 0 2096 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_6067
timestamp 1680363874
transform 1 0 2148 0 1 1575
box -3 -3 3 3
use FILL  FILL_7700
timestamp 1680363874
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7701
timestamp 1680363874
transform 1 0 2144 0 1 1570
box -8 -3 16 105
use FILL  FILL_7702
timestamp 1680363874
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_7703
timestamp 1680363874
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_7705
timestamp 1680363874
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6068
timestamp 1680363874
transform 1 0 2196 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_302
timestamp 1680363874
transform 1 0 2176 0 1 1570
box -8 -3 46 105
use FILL  FILL_7707
timestamp 1680363874
transform 1 0 2216 0 1 1570
box -8 -3 16 105
use FILL  FILL_7712
timestamp 1680363874
transform 1 0 2224 0 1 1570
box -8 -3 16 105
use FILL  FILL_7714
timestamp 1680363874
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_401
timestamp 1680363874
transform 1 0 2240 0 1 1570
box -8 -3 104 105
use FILL  FILL_7715
timestamp 1680363874
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6069
timestamp 1680363874
transform 1 0 2380 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_402
timestamp 1680363874
transform 1 0 2344 0 1 1570
box -8 -3 104 105
use FILL  FILL_7716
timestamp 1680363874
transform 1 0 2440 0 1 1570
box -8 -3 16 105
use FILL  FILL_7717
timestamp 1680363874
transform 1 0 2448 0 1 1570
box -8 -3 16 105
use FILL  FILL_7718
timestamp 1680363874
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_84
timestamp 1680363874
transform -1 0 2488 0 1 1570
box -8 -3 32 105
use FILL  FILL_7719
timestamp 1680363874
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_7731
timestamp 1680363874
transform 1 0 2496 0 1 1570
box -8 -3 16 105
use AND2X2  AND2X2_45
timestamp 1680363874
transform 1 0 2504 0 1 1570
box -8 -3 40 105
use FILL  FILL_7733
timestamp 1680363874
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7737
timestamp 1680363874
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7739
timestamp 1680363874
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7740
timestamp 1680363874
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6070
timestamp 1680363874
transform 1 0 2612 0 1 1575
box -3 -3 3 3
use NAND3X1  NAND3X1_55
timestamp 1680363874
transform -1 0 2600 0 1 1570
box -8 -3 40 105
use FILL  FILL_7741
timestamp 1680363874
transform 1 0 2600 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_56
timestamp 1680363874
transform 1 0 2608 0 1 1570
box -8 -3 40 105
use FILL  FILL_7742
timestamp 1680363874
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_7749
timestamp 1680363874
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use FILL  FILL_7750
timestamp 1680363874
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_7751
timestamp 1680363874
transform 1 0 2664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7752
timestamp 1680363874
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_58
timestamp 1680363874
transform 1 0 2680 0 1 1570
box -8 -3 40 105
use FILL  FILL_7753
timestamp 1680363874
transform 1 0 2712 0 1 1570
box -8 -3 16 105
use FILL  FILL_7759
timestamp 1680363874
transform 1 0 2720 0 1 1570
box -8 -3 16 105
use FILL  FILL_7761
timestamp 1680363874
transform 1 0 2728 0 1 1570
box -8 -3 16 105
use FILL  FILL_7763
timestamp 1680363874
transform 1 0 2736 0 1 1570
box -8 -3 16 105
use FILL  FILL_7764
timestamp 1680363874
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_59
timestamp 1680363874
transform 1 0 2752 0 1 1570
box -8 -3 40 105
use FILL  FILL_7765
timestamp 1680363874
transform 1 0 2784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7769
timestamp 1680363874
transform 1 0 2792 0 1 1570
box -8 -3 16 105
use FILL  FILL_7771
timestamp 1680363874
transform 1 0 2800 0 1 1570
box -8 -3 16 105
use FILL  FILL_7772
timestamp 1680363874
transform 1 0 2808 0 1 1570
box -8 -3 16 105
use FILL  FILL_7773
timestamp 1680363874
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_77
timestamp 1680363874
transform 1 0 2824 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_78
timestamp 1680363874
transform 1 0 2848 0 1 1570
box -5 -3 28 105
use FILL  FILL_7774
timestamp 1680363874
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_7775
timestamp 1680363874
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_403
timestamp 1680363874
transform -1 0 2984 0 1 1570
box -8 -3 104 105
use FILL  FILL_7776
timestamp 1680363874
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_404
timestamp 1680363874
transform -1 0 3088 0 1 1570
box -8 -3 104 105
use FILL  FILL_7777
timestamp 1680363874
transform 1 0 3088 0 1 1570
box -8 -3 16 105
use FILL  FILL_7778
timestamp 1680363874
transform 1 0 3096 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_467
timestamp 1680363874
transform 1 0 3104 0 1 1570
box -9 -3 26 105
use FILL  FILL_7779
timestamp 1680363874
transform 1 0 3120 0 1 1570
box -8 -3 16 105
use FILL  FILL_7804
timestamp 1680363874
transform 1 0 3128 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_79
timestamp 1680363874
transform 1 0 3136 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_80
timestamp 1680363874
transform 1 0 3160 0 1 1570
box -5 -3 28 105
use FILL  FILL_7806
timestamp 1680363874
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_405
timestamp 1680363874
transform 1 0 3192 0 1 1570
box -8 -3 104 105
use FILL  FILL_7807
timestamp 1680363874
transform 1 0 3288 0 1 1570
box -8 -3 16 105
use FILL  FILL_7816
timestamp 1680363874
transform 1 0 3296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7818
timestamp 1680363874
transform 1 0 3304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7819
timestamp 1680363874
transform 1 0 3312 0 1 1570
box -8 -3 16 105
use FILL  FILL_7820
timestamp 1680363874
transform 1 0 3320 0 1 1570
box -8 -3 16 105
use FILL  FILL_7821
timestamp 1680363874
transform 1 0 3328 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_249
timestamp 1680363874
transform 1 0 3336 0 1 1570
box -8 -3 46 105
use FILL  FILL_7824
timestamp 1680363874
transform 1 0 3376 0 1 1570
box -8 -3 16 105
use FILL  FILL_7831
timestamp 1680363874
transform 1 0 3384 0 1 1570
box -8 -3 16 105
use FILL  FILL_7833
timestamp 1680363874
transform 1 0 3392 0 1 1570
box -8 -3 16 105
use FILL  FILL_7835
timestamp 1680363874
transform 1 0 3400 0 1 1570
box -8 -3 16 105
use FILL  FILL_7837
timestamp 1680363874
transform 1 0 3408 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6071
timestamp 1680363874
transform 1 0 3428 0 1 1575
box -3 -3 3 3
use FILL  FILL_7839
timestamp 1680363874
transform 1 0 3416 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_86
timestamp 1680363874
transform 1 0 3424 0 1 1570
box -8 -3 32 105
use FILL  FILL_7840
timestamp 1680363874
transform 1 0 3448 0 1 1570
box -8 -3 16 105
use FILL  FILL_7841
timestamp 1680363874
transform 1 0 3456 0 1 1570
box -8 -3 16 105
use FILL  FILL_7842
timestamp 1680363874
transform 1 0 3464 0 1 1570
box -8 -3 16 105
use FILL  FILL_7845
timestamp 1680363874
transform 1 0 3472 0 1 1570
box -8 -3 16 105
use FILL  FILL_7847
timestamp 1680363874
transform 1 0 3480 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6072
timestamp 1680363874
transform 1 0 3500 0 1 1575
box -3 -3 3 3
use FILL  FILL_7848
timestamp 1680363874
transform 1 0 3488 0 1 1570
box -8 -3 16 105
use FILL  FILL_7849
timestamp 1680363874
transform 1 0 3496 0 1 1570
box -8 -3 16 105
use FILL  FILL_7850
timestamp 1680363874
transform 1 0 3504 0 1 1570
box -8 -3 16 105
use FILL  FILL_7851
timestamp 1680363874
transform 1 0 3512 0 1 1570
box -8 -3 16 105
use FILL  FILL_7852
timestamp 1680363874
transform 1 0 3520 0 1 1570
box -8 -3 16 105
use FILL  FILL_7853
timestamp 1680363874
transform 1 0 3528 0 1 1570
box -8 -3 16 105
use FILL  FILL_7856
timestamp 1680363874
transform 1 0 3536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7858
timestamp 1680363874
transform 1 0 3544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7860
timestamp 1680363874
transform 1 0 3552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7862
timestamp 1680363874
transform 1 0 3560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7863
timestamp 1680363874
transform 1 0 3568 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_250
timestamp 1680363874
transform -1 0 3616 0 1 1570
box -8 -3 46 105
use FILL  FILL_7864
timestamp 1680363874
transform 1 0 3616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7865
timestamp 1680363874
transform 1 0 3624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7866
timestamp 1680363874
transform 1 0 3632 0 1 1570
box -8 -3 16 105
use FILL  FILL_7867
timestamp 1680363874
transform 1 0 3640 0 1 1570
box -8 -3 16 105
use FILL  FILL_7868
timestamp 1680363874
transform 1 0 3648 0 1 1570
box -8 -3 16 105
use FILL  FILL_7869
timestamp 1680363874
transform 1 0 3656 0 1 1570
box -8 -3 16 105
use FILL  FILL_7870
timestamp 1680363874
transform 1 0 3664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7871
timestamp 1680363874
transform 1 0 3672 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6073
timestamp 1680363874
transform 1 0 3788 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_407
timestamp 1680363874
transform 1 0 3680 0 1 1570
box -8 -3 104 105
use FILL  FILL_7872
timestamp 1680363874
transform 1 0 3776 0 1 1570
box -8 -3 16 105
use FILL  FILL_7873
timestamp 1680363874
transform 1 0 3784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7874
timestamp 1680363874
transform 1 0 3792 0 1 1570
box -8 -3 16 105
use FILL  FILL_7875
timestamp 1680363874
transform 1 0 3800 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6074
timestamp 1680363874
transform 1 0 3852 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_251
timestamp 1680363874
transform 1 0 3808 0 1 1570
box -8 -3 46 105
use FILL  FILL_7883
timestamp 1680363874
transform 1 0 3848 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_409
timestamp 1680363874
transform 1 0 3856 0 1 1570
box -8 -3 104 105
use FILL  FILL_7884
timestamp 1680363874
transform 1 0 3952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7885
timestamp 1680363874
transform 1 0 3960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7901
timestamp 1680363874
transform 1 0 3968 0 1 1570
box -8 -3 16 105
use FILL  FILL_7903
timestamp 1680363874
transform 1 0 3976 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_308
timestamp 1680363874
transform -1 0 4024 0 1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_410
timestamp 1680363874
transform 1 0 4024 0 1 1570
box -8 -3 104 105
use OAI22X1  OAI22X1_309
timestamp 1680363874
transform 1 0 4120 0 1 1570
box -8 -3 46 105
use FILL  FILL_7904
timestamp 1680363874
transform 1 0 4160 0 1 1570
box -8 -3 16 105
use FILL  FILL_7922
timestamp 1680363874
transform 1 0 4168 0 1 1570
box -8 -3 16 105
use FILL  FILL_7924
timestamp 1680363874
transform 1 0 4176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7926
timestamp 1680363874
transform 1 0 4184 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_474
timestamp 1680363874
transform 1 0 4192 0 1 1570
box -9 -3 26 105
use FILL  FILL_7928
timestamp 1680363874
transform 1 0 4208 0 1 1570
box -8 -3 16 105
use FILL  FILL_7932
timestamp 1680363874
transform 1 0 4216 0 1 1570
box -8 -3 16 105
use FILL  FILL_7934
timestamp 1680363874
transform 1 0 4224 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_411
timestamp 1680363874
transform 1 0 4232 0 1 1570
box -8 -3 104 105
use FILL  FILL_7936
timestamp 1680363874
transform 1 0 4328 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_412
timestamp 1680363874
transform 1 0 4336 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_475
timestamp 1680363874
transform -1 0 4448 0 1 1570
box -9 -3 26 105
use FILL  FILL_7937
timestamp 1680363874
transform 1 0 4448 0 1 1570
box -8 -3 16 105
use FILL  FILL_7958
timestamp 1680363874
transform 1 0 4456 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6075
timestamp 1680363874
transform 1 0 4476 0 1 1575
box -3 -3 3 3
use FILL  FILL_7959
timestamp 1680363874
transform 1 0 4464 0 1 1570
box -8 -3 16 105
use FILL  FILL_7960
timestamp 1680363874
transform 1 0 4472 0 1 1570
box -8 -3 16 105
use FILL  FILL_7961
timestamp 1680363874
transform 1 0 4480 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_253
timestamp 1680363874
transform -1 0 4528 0 1 1570
box -8 -3 46 105
use FILL  FILL_7962
timestamp 1680363874
transform 1 0 4528 0 1 1570
box -8 -3 16 105
use FILL  FILL_7963
timestamp 1680363874
transform 1 0 4536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7964
timestamp 1680363874
transform 1 0 4544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7965
timestamp 1680363874
transform 1 0 4552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7971
timestamp 1680363874
transform 1 0 4560 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_91
timestamp 1680363874
transform 1 0 4568 0 1 1570
box -8 -3 32 105
use FILL  FILL_7973
timestamp 1680363874
transform 1 0 4592 0 1 1570
box -8 -3 16 105
use FILL  FILL_7974
timestamp 1680363874
transform 1 0 4600 0 1 1570
box -8 -3 16 105
use FILL  FILL_7975
timestamp 1680363874
transform 1 0 4608 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6076
timestamp 1680363874
transform 1 0 4636 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_312
timestamp 1680363874
transform -1 0 4656 0 1 1570
box -8 -3 46 105
use FILL  FILL_7976
timestamp 1680363874
transform 1 0 4656 0 1 1570
box -8 -3 16 105
use FILL  FILL_7977
timestamp 1680363874
transform 1 0 4664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7978
timestamp 1680363874
transform 1 0 4672 0 1 1570
box -8 -3 16 105
use FILL  FILL_7979
timestamp 1680363874
transform 1 0 4680 0 1 1570
box -8 -3 16 105
use FILL  FILL_7980
timestamp 1680363874
transform 1 0 4688 0 1 1570
box -8 -3 16 105
use FILL  FILL_7981
timestamp 1680363874
transform 1 0 4696 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_413
timestamp 1680363874
transform 1 0 4704 0 1 1570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_63
timestamp 1680363874
transform 1 0 4827 0 1 1570
box -10 -3 10 3
use M2_M1  M2_M1_6635
timestamp 1680363874
transform 1 0 92 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_6168
timestamp 1680363874
transform 1 0 92 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6643
timestamp 1680363874
transform 1 0 124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6738
timestamp 1680363874
transform 1 0 116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1680363874
transform 1 0 164 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6169
timestamp 1680363874
transform 1 0 164 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6739
timestamp 1680363874
transform 1 0 188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6740
timestamp 1680363874
transform 1 0 244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1680363874
transform 1 0 276 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_6170
timestamp 1680363874
transform 1 0 268 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6741
timestamp 1680363874
transform 1 0 316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1680363874
transform 1 0 356 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6140
timestamp 1680363874
transform 1 0 364 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6742
timestamp 1680363874
transform 1 0 364 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1680363874
transform 1 0 372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1680363874
transform 1 0 388 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_6141
timestamp 1680363874
transform 1 0 460 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6647
timestamp 1680363874
transform 1 0 492 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6171
timestamp 1680363874
transform 1 0 388 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6743
timestamp 1680363874
transform 1 0 476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6744
timestamp 1680363874
transform 1 0 484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6210
timestamp 1680363874
transform 1 0 460 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6745
timestamp 1680363874
transform 1 0 500 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6118
timestamp 1680363874
transform 1 0 524 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6648
timestamp 1680363874
transform 1 0 524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1680363874
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1680363874
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6172
timestamp 1680363874
transform 1 0 548 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6077
timestamp 1680363874
transform 1 0 588 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6747
timestamp 1680363874
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6078
timestamp 1680363874
transform 1 0 612 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1680363874
transform 1 0 620 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1680363874
transform 1 0 644 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6650
timestamp 1680363874
transform 1 0 596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1680363874
transform 1 0 644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6748
timestamp 1680363874
transform 1 0 612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1680363874
transform 1 0 660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1680363874
transform 1 0 692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6750
timestamp 1680363874
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6090
timestamp 1680363874
transform 1 0 740 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6653
timestamp 1680363874
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6187
timestamp 1680363874
transform 1 0 764 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1680363874
transform 1 0 772 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6654
timestamp 1680363874
transform 1 0 772 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6173
timestamp 1680363874
transform 1 0 772 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6224
timestamp 1680363874
transform 1 0 788 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6751
timestamp 1680363874
transform 1 0 804 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6119
timestamp 1680363874
transform 1 0 852 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6655
timestamp 1680363874
transform 1 0 836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1680363874
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6092
timestamp 1680363874
transform 1 0 868 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6142
timestamp 1680363874
transform 1 0 868 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6752
timestamp 1680363874
transform 1 0 844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6753
timestamp 1680363874
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6754
timestamp 1680363874
transform 1 0 868 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6188
timestamp 1680363874
transform 1 0 844 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6120
timestamp 1680363874
transform 1 0 988 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6657
timestamp 1680363874
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1680363874
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6755
timestamp 1680363874
transform 1 0 900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6756
timestamp 1680363874
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6231
timestamp 1680363874
transform 1 0 1148 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6189
timestamp 1680363874
transform 1 0 1228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6121
timestamp 1680363874
transform 1 0 1244 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6659
timestamp 1680363874
transform 1 0 1244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6757
timestamp 1680363874
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6758
timestamp 1680363874
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6190
timestamp 1680363874
transform 1 0 1268 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6211
timestamp 1680363874
transform 1 0 1308 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6232
timestamp 1680363874
transform 1 0 1260 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6191
timestamp 1680363874
transform 1 0 1332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6212
timestamp 1680363874
transform 1 0 1332 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6660
timestamp 1680363874
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1680363874
transform 1 0 1396 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6192
timestamp 1680363874
transform 1 0 1396 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1680363874
transform 1 0 1420 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6759
timestamp 1680363874
transform 1 0 1412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6760
timestamp 1680363874
transform 1 0 1444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6123
timestamp 1680363874
transform 1 0 1484 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6662
timestamp 1680363874
transform 1 0 1460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1680363874
transform 1 0 1476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1680363874
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6213
timestamp 1680363874
transform 1 0 1460 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6214
timestamp 1680363874
transform 1 0 1492 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1680363874
transform 1 0 1508 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6664
timestamp 1680363874
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6762
timestamp 1680363874
transform 1 0 1508 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6124
timestamp 1680363874
transform 1 0 1556 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6094
timestamp 1680363874
transform 1 0 1588 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6665
timestamp 1680363874
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1680363874
transform 1 0 1572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1680363874
transform 1 0 1588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6763
timestamp 1680363874
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6764
timestamp 1680363874
transform 1 0 1580 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6193
timestamp 1680363874
transform 1 0 1580 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1680363874
transform 1 0 1604 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6765
timestamp 1680363874
transform 1 0 1612 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6215
timestamp 1680363874
transform 1 0 1620 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6079
timestamp 1680363874
transform 1 0 1644 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6095
timestamp 1680363874
transform 1 0 1652 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1680363874
transform 1 0 1692 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6668
timestamp 1680363874
transform 1 0 1668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1680363874
transform 1 0 1684 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6766
timestamp 1680363874
transform 1 0 1676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6767
timestamp 1680363874
transform 1 0 1692 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6194
timestamp 1680363874
transform 1 0 1684 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6216
timestamp 1680363874
transform 1 0 1668 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6217
timestamp 1680363874
transform 1 0 1700 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6768
timestamp 1680363874
transform 1 0 1732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1680363874
transform 1 0 1748 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6097
timestamp 1680363874
transform 1 0 1764 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6671
timestamp 1680363874
transform 1 0 1764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1680363874
transform 1 0 1756 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6098
timestamp 1680363874
transform 1 0 1804 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6672
timestamp 1680363874
transform 1 0 1788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1680363874
transform 1 0 1796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1680363874
transform 1 0 1812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1680363874
transform 1 0 1788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6771
timestamp 1680363874
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6772
timestamp 1680363874
transform 1 0 1836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1680363874
transform 1 0 1844 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6099
timestamp 1680363874
transform 1 0 1892 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1680363874
transform 1 0 1924 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6675
timestamp 1680363874
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6774
timestamp 1680363874
transform 1 0 1876 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6195
timestamp 1680363874
transform 1 0 1884 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6676
timestamp 1680363874
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6775
timestamp 1680363874
transform 1 0 1924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6776
timestamp 1680363874
transform 1 0 1980 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6126
timestamp 1680363874
transform 1 0 2060 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6101
timestamp 1680363874
transform 1 0 2140 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6677
timestamp 1680363874
transform 1 0 2076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6777
timestamp 1680363874
transform 1 0 2116 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6127
timestamp 1680363874
transform 1 0 2204 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6778
timestamp 1680363874
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6779
timestamp 1680363874
transform 1 0 2196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1680363874
transform 1 0 2204 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6218
timestamp 1680363874
transform 1 0 2228 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6679
timestamp 1680363874
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6780
timestamp 1680363874
transform 1 0 2260 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6219
timestamp 1680363874
transform 1 0 2260 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6781
timestamp 1680363874
transform 1 0 2276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1680363874
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6102
timestamp 1680363874
transform 1 0 2324 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6681
timestamp 1680363874
transform 1 0 2316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6782
timestamp 1680363874
transform 1 0 2316 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6220
timestamp 1680363874
transform 1 0 2316 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6682
timestamp 1680363874
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1680363874
transform 1 0 2364 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6143
timestamp 1680363874
transform 1 0 2380 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6783
timestamp 1680363874
transform 1 0 2388 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6103
timestamp 1680363874
transform 1 0 2412 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6638
timestamp 1680363874
transform 1 0 2420 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_6144
timestamp 1680363874
transform 1 0 2420 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1680363874
transform 1 0 2452 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6684
timestamp 1680363874
transform 1 0 2428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1680363874
transform 1 0 2444 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6145
timestamp 1680363874
transform 1 0 2452 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6146
timestamp 1680363874
transform 1 0 2476 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6686
timestamp 1680363874
transform 1 0 2484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6784
timestamp 1680363874
transform 1 0 2452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6785
timestamp 1680363874
transform 1 0 2468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6786
timestamp 1680363874
transform 1 0 2476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6787
timestamp 1680363874
transform 1 0 2484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6221
timestamp 1680363874
transform 1 0 2484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6225
timestamp 1680363874
transform 1 0 2500 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6128
timestamp 1680363874
transform 1 0 2532 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6687
timestamp 1680363874
transform 1 0 2532 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6129
timestamp 1680363874
transform 1 0 2564 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6688
timestamp 1680363874
transform 1 0 2556 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6147
timestamp 1680363874
transform 1 0 2588 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6788
timestamp 1680363874
transform 1 0 2588 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6080
timestamp 1680363874
transform 1 0 2604 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6148
timestamp 1680363874
transform 1 0 2620 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6789
timestamp 1680363874
transform 1 0 2620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6838
timestamp 1680363874
transform 1 0 2604 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6839
timestamp 1680363874
transform 1 0 2628 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6845
timestamp 1680363874
transform 1 0 2612 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6226
timestamp 1680363874
transform 1 0 2628 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6840
timestamp 1680363874
transform 1 0 2644 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1680363874
transform 1 0 2660 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6174
timestamp 1680363874
transform 1 0 2660 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6690
timestamp 1680363874
transform 1 0 2692 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6149
timestamp 1680363874
transform 1 0 2700 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1680363874
transform 1 0 2700 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6846
timestamp 1680363874
transform 1 0 2708 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6227
timestamp 1680363874
transform 1 0 2708 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6790
timestamp 1680363874
transform 1 0 2732 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6150
timestamp 1680363874
transform 1 0 2748 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6791
timestamp 1680363874
transform 1 0 2748 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6841
timestamp 1680363874
transform 1 0 2740 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1680363874
transform 1 0 2756 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6842
timestamp 1680363874
transform 1 0 2796 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1680363874
transform 1 0 2812 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6151
timestamp 1680363874
transform 1 0 2820 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6692
timestamp 1680363874
transform 1 0 2828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1680363874
transform 1 0 2820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6793
timestamp 1680363874
transform 1 0 2860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1680363874
transform 1 0 2868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1680363874
transform 1 0 2876 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6176
timestamp 1680363874
transform 1 0 2876 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6695
timestamp 1680363874
transform 1 0 2892 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6177
timestamp 1680363874
transform 1 0 2900 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6196
timestamp 1680363874
transform 1 0 2908 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6152
timestamp 1680363874
transform 1 0 2940 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6130
timestamp 1680363874
transform 1 0 2964 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6696
timestamp 1680363874
transform 1 0 2964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1680363874
transform 1 0 2980 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6153
timestamp 1680363874
transform 1 0 2988 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6794
timestamp 1680363874
transform 1 0 2948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6795
timestamp 1680363874
transform 1 0 2956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6796
timestamp 1680363874
transform 1 0 2972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6797
timestamp 1680363874
transform 1 0 2988 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6131
timestamp 1680363874
transform 1 0 3004 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6698
timestamp 1680363874
transform 1 0 3004 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6178
timestamp 1680363874
transform 1 0 3076 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6699
timestamp 1680363874
transform 1 0 3092 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6154
timestamp 1680363874
transform 1 0 3116 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6798
timestamp 1680363874
transform 1 0 3084 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1680363874
transform 1 0 3100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1680363874
transform 1 0 3116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1680363874
transform 1 0 3124 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6105
timestamp 1680363874
transform 1 0 3148 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6132
timestamp 1680363874
transform 1 0 3252 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6155
timestamp 1680363874
transform 1 0 3220 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6700
timestamp 1680363874
transform 1 0 3252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6802
timestamp 1680363874
transform 1 0 3204 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6179
timestamp 1680363874
transform 1 0 3252 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1680363874
transform 1 0 3276 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6701
timestamp 1680363874
transform 1 0 3268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6803
timestamp 1680363874
transform 1 0 3276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1680363874
transform 1 0 3300 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6180
timestamp 1680363874
transform 1 0 3300 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1680363874
transform 1 0 3316 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6703
timestamp 1680363874
transform 1 0 3332 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6107
timestamp 1680363874
transform 1 0 3364 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6704
timestamp 1680363874
transform 1 0 3356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6804
timestamp 1680363874
transform 1 0 3348 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6081
timestamp 1680363874
transform 1 0 3396 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6134
timestamp 1680363874
transform 1 0 3412 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6705
timestamp 1680363874
transform 1 0 3444 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6156
timestamp 1680363874
transform 1 0 3452 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6181
timestamp 1680363874
transform 1 0 3428 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6805
timestamp 1680363874
transform 1 0 3436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1680363874
transform 1 0 3452 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6197
timestamp 1680363874
transform 1 0 3468 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1680363874
transform 1 0 3492 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6135
timestamp 1680363874
transform 1 0 3508 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6706
timestamp 1680363874
transform 1 0 3484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1680363874
transform 1 0 3492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1680363874
transform 1 0 3508 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6157
timestamp 1680363874
transform 1 0 3516 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6182
timestamp 1680363874
transform 1 0 3492 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6807
timestamp 1680363874
transform 1 0 3500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1680363874
transform 1 0 3516 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6198
timestamp 1680363874
transform 1 0 3500 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6233
timestamp 1680363874
transform 1 0 3492 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6709
timestamp 1680363874
transform 1 0 3532 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6183
timestamp 1680363874
transform 1 0 3532 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6809
timestamp 1680363874
transform 1 0 3556 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6222
timestamp 1680363874
transform 1 0 3564 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6710
timestamp 1680363874
transform 1 0 3580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1680363874
transform 1 0 3580 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6082
timestamp 1680363874
transform 1 0 3700 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1680363874
transform 1 0 3692 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6639
timestamp 1680363874
transform 1 0 3692 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1680363874
transform 1 0 3676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6811
timestamp 1680363874
transform 1 0 3588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6812
timestamp 1680363874
transform 1 0 3596 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6184
timestamp 1680363874
transform 1 0 3604 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6813
timestamp 1680363874
transform 1 0 3628 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6199
timestamp 1680363874
transform 1 0 3588 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6200
timestamp 1680363874
transform 1 0 3628 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6223
timestamp 1680363874
transform 1 0 3588 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6712
timestamp 1680363874
transform 1 0 3700 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6158
timestamp 1680363874
transform 1 0 3740 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1680363874
transform 1 0 3764 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1680363874
transform 1 0 3780 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6110
timestamp 1680363874
transform 1 0 3780 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6713
timestamp 1680363874
transform 1 0 3764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1680363874
transform 1 0 3780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1680363874
transform 1 0 3796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6814
timestamp 1680363874
transform 1 0 3756 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6201
timestamp 1680363874
transform 1 0 3756 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6815
timestamp 1680363874
transform 1 0 3772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6816
timestamp 1680363874
transform 1 0 3788 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6234
timestamp 1680363874
transform 1 0 3764 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6159
timestamp 1680363874
transform 1 0 3804 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6817
timestamp 1680363874
transform 1 0 3804 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6202
timestamp 1680363874
transform 1 0 3812 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6085
timestamp 1680363874
transform 1 0 3836 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6716
timestamp 1680363874
transform 1 0 3828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1680363874
transform 1 0 3900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6818
timestamp 1680363874
transform 1 0 3932 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6235
timestamp 1680363874
transform 1 0 3980 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6640
timestamp 1680363874
transform 1 0 4004 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6819
timestamp 1680363874
transform 1 0 4060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1680363874
transform 1 0 4084 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1680363874
transform 1 0 4116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1680363874
transform 1 0 4124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1680363874
transform 1 0 4140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6821
timestamp 1680363874
transform 1 0 4132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6203
timestamp 1680363874
transform 1 0 4116 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6204
timestamp 1680363874
transform 1 0 4132 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6822
timestamp 1680363874
transform 1 0 4156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6823
timestamp 1680363874
transform 1 0 4172 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6228
timestamp 1680363874
transform 1 0 4196 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6843
timestamp 1680363874
transform 1 0 4212 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6844
timestamp 1680363874
transform 1 0 4260 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6160
timestamp 1680363874
transform 1 0 4284 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6721
timestamp 1680363874
transform 1 0 4292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1680363874
transform 1 0 4300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1680363874
transform 1 0 4324 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6111
timestamp 1680363874
transform 1 0 4340 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6724
timestamp 1680363874
transform 1 0 4348 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6161
timestamp 1680363874
transform 1 0 4356 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6824
timestamp 1680363874
transform 1 0 4332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6825
timestamp 1680363874
transform 1 0 4356 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6205
timestamp 1680363874
transform 1 0 4332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1680363874
transform 1 0 4372 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6641
timestamp 1680363874
transform 1 0 4372 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1680363874
transform 1 0 4388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1680363874
transform 1 0 4412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6826
timestamp 1680363874
transform 1 0 4404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6827
timestamp 1680363874
transform 1 0 4412 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6206
timestamp 1680363874
transform 1 0 4412 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6727
timestamp 1680363874
transform 1 0 4428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1680363874
transform 1 0 4476 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6162
timestamp 1680363874
transform 1 0 4484 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6729
timestamp 1680363874
transform 1 0 4492 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6185
timestamp 1680363874
transform 1 0 4468 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6828
timestamp 1680363874
transform 1 0 4484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6229
timestamp 1680363874
transform 1 0 4484 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6236
timestamp 1680363874
transform 1 0 4484 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6163
timestamp 1680363874
transform 1 0 4500 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6237
timestamp 1680363874
transform 1 0 4500 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6136
timestamp 1680363874
transform 1 0 4516 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1680363874
transform 1 0 4532 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6642
timestamp 1680363874
transform 1 0 4532 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1680363874
transform 1 0 4524 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6238
timestamp 1680363874
transform 1 0 4540 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6164
timestamp 1680363874
transform 1 0 4564 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6829
timestamp 1680363874
transform 1 0 4564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6731
timestamp 1680363874
transform 1 0 4572 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6086
timestamp 1680363874
transform 1 0 4604 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6114
timestamp 1680363874
transform 1 0 4596 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6137
timestamp 1680363874
transform 1 0 4588 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6165
timestamp 1680363874
transform 1 0 4588 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6732
timestamp 1680363874
transform 1 0 4596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6830
timestamp 1680363874
transform 1 0 4588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6831
timestamp 1680363874
transform 1 0 4604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6207
timestamp 1680363874
transform 1 0 4604 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6230
timestamp 1680363874
transform 1 0 4588 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6166
timestamp 1680363874
transform 1 0 4628 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1680363874
transform 1 0 4644 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6115
timestamp 1680363874
transform 1 0 4644 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1680363874
transform 1 0 4668 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1680363874
transform 1 0 4660 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6139
timestamp 1680363874
transform 1 0 4676 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6733
timestamp 1680363874
transform 1 0 4644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6734
timestamp 1680363874
transform 1 0 4652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1680363874
transform 1 0 4668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6736
timestamp 1680363874
transform 1 0 4676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6832
timestamp 1680363874
transform 1 0 4636 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6239
timestamp 1680363874
transform 1 0 4628 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6186
timestamp 1680363874
transform 1 0 4652 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6833
timestamp 1680363874
transform 1 0 4660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1680363874
transform 1 0 4676 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6167
timestamp 1680363874
transform 1 0 4692 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6117
timestamp 1680363874
transform 1 0 4788 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6737
timestamp 1680363874
transform 1 0 4708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6835
timestamp 1680363874
transform 1 0 4692 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6836
timestamp 1680363874
transform 1 0 4732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6837
timestamp 1680363874
transform 1 0 4788 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6208
timestamp 1680363874
transform 1 0 4692 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6209
timestamp 1680363874
transform 1 0 4732 0 1 1515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_64
timestamp 1680363874
transform 1 0 24 0 1 1470
box -10 -3 10 3
use FILL  FILL_7468
timestamp 1680363874
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7470
timestamp 1680363874
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7472
timestamp 1680363874
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_83
timestamp 1680363874
transform 1 0 96 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7474
timestamp 1680363874
transform 1 0 120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7476
timestamp 1680363874
transform 1 0 128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7478
timestamp 1680363874
transform 1 0 136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7480
timestamp 1680363874
transform 1 0 144 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_392
timestamp 1680363874
transform 1 0 152 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7490
timestamp 1680363874
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7500
timestamp 1680363874
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7501
timestamp 1680363874
transform 1 0 264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7502
timestamp 1680363874
transform 1 0 272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7503
timestamp 1680363874
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7504
timestamp 1680363874
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7505
timestamp 1680363874
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7506
timestamp 1680363874
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_14
timestamp 1680363874
transform -1 0 344 0 -1 1570
box -7 -3 39 105
use FILL  FILL_7507
timestamp 1680363874
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7508
timestamp 1680363874
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7509
timestamp 1680363874
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7510
timestamp 1680363874
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FAX1  FAX1_23
timestamp 1680363874
transform -1 0 496 0 -1 1570
box -5 -3 126 105
use FILL  FILL_7511
timestamp 1680363874
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7512
timestamp 1680363874
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7513
timestamp 1680363874
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_243
timestamp 1680363874
transform 1 0 520 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7514
timestamp 1680363874
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7515
timestamp 1680363874
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7516
timestamp 1680363874
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7517
timestamp 1680363874
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_3
timestamp 1680363874
transform -1 0 648 0 -1 1570
box -8 -3 64 105
use FILL  FILL_7518
timestamp 1680363874
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7519
timestamp 1680363874
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7520
timestamp 1680363874
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7521
timestamp 1680363874
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_15
timestamp 1680363874
transform 1 0 680 0 -1 1570
box -7 -3 39 105
use FILL  FILL_7522
timestamp 1680363874
transform 1 0 712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7523
timestamp 1680363874
transform 1 0 720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7524
timestamp 1680363874
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7525
timestamp 1680363874
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_451
timestamp 1680363874
transform -1 0 760 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7526
timestamp 1680363874
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7527
timestamp 1680363874
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7528
timestamp 1680363874
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7530
timestamp 1680363874
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7542
timestamp 1680363874
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7543
timestamp 1680363874
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7544
timestamp 1680363874
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7545
timestamp 1680363874
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_244
timestamp 1680363874
transform -1 0 864 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7546
timestamp 1680363874
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7547
timestamp 1680363874
transform 1 0 872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7548
timestamp 1680363874
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_453
timestamp 1680363874
transform -1 0 904 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_396
timestamp 1680363874
transform -1 0 1000 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7549
timestamp 1680363874
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7550
timestamp 1680363874
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7551
timestamp 1680363874
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7552
timestamp 1680363874
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7553
timestamp 1680363874
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7554
timestamp 1680363874
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7555
timestamp 1680363874
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7556
timestamp 1680363874
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7557
timestamp 1680363874
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7558
timestamp 1680363874
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7559
timestamp 1680363874
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7561
timestamp 1680363874
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7563
timestamp 1680363874
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7564
timestamp 1680363874
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7565
timestamp 1680363874
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7567
timestamp 1680363874
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7569
timestamp 1680363874
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7571
timestamp 1680363874
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7574
timestamp 1680363874
transform 1 0 1144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7575
timestamp 1680363874
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7576
timestamp 1680363874
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7577
timestamp 1680363874
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7578
timestamp 1680363874
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7579
timestamp 1680363874
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7580
timestamp 1680363874
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7582
timestamp 1680363874
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7584
timestamp 1680363874
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7586
timestamp 1680363874
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7588
timestamp 1680363874
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_397
timestamp 1680363874
transform 1 0 1232 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7600
timestamp 1680363874
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7602
timestamp 1680363874
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7603
timestamp 1680363874
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7604
timestamp 1680363874
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7605
timestamp 1680363874
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7606
timestamp 1680363874
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7607
timestamp 1680363874
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7611
timestamp 1680363874
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_73
timestamp 1680363874
transform -1 0 1416 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7612
timestamp 1680363874
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7613
timestamp 1680363874
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7614
timestamp 1680363874
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7615
timestamp 1680363874
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7616
timestamp 1680363874
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_295
timestamp 1680363874
transform 1 0 1456 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7617
timestamp 1680363874
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7619
timestamp 1680363874
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7621
timestamp 1680363874
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7622
timestamp 1680363874
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7623
timestamp 1680363874
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7625
timestamp 1680363874
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7627
timestamp 1680363874
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_296
timestamp 1680363874
transform 1 0 1552 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7632
timestamp 1680363874
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7634
timestamp 1680363874
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7636
timestamp 1680363874
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7638
timestamp 1680363874
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7640
timestamp 1680363874
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7642
timestamp 1680363874
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7646
timestamp 1680363874
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7647
timestamp 1680363874
transform 1 0 1648 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_245
timestamp 1680363874
transform 1 0 1656 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7648
timestamp 1680363874
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7650
timestamp 1680363874
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7652
timestamp 1680363874
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7656
timestamp 1680363874
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_74
timestamp 1680363874
transform 1 0 1728 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7657
timestamp 1680363874
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7659
timestamp 1680363874
transform 1 0 1760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7661
timestamp 1680363874
transform 1 0 1768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7664
timestamp 1680363874
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_246
timestamp 1680363874
transform -1 0 1824 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7665
timestamp 1680363874
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7670
timestamp 1680363874
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_459
timestamp 1680363874
transform -1 0 1856 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7671
timestamp 1680363874
transform 1 0 1856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7673
timestamp 1680363874
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7680
timestamp 1680363874
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7681
timestamp 1680363874
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_399
timestamp 1680363874
transform 1 0 1888 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7682
timestamp 1680363874
transform 1 0 1984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7684
timestamp 1680363874
transform 1 0 1992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7686
timestamp 1680363874
transform 1 0 2000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7688
timestamp 1680363874
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7689
timestamp 1680363874
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7690
timestamp 1680363874
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7691
timestamp 1680363874
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7692
timestamp 1680363874
transform 1 0 2040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7693
timestamp 1680363874
transform 1 0 2048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7695
timestamp 1680363874
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_400
timestamp 1680363874
transform 1 0 2064 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7704
timestamp 1680363874
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7706
timestamp 1680363874
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_462
timestamp 1680363874
transform 1 0 2176 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7708
timestamp 1680363874
transform 1 0 2192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7709
timestamp 1680363874
transform 1 0 2200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7710
timestamp 1680363874
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7711
timestamp 1680363874
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7713
timestamp 1680363874
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_303
timestamp 1680363874
transform 1 0 2232 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7720
timestamp 1680363874
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7721
timestamp 1680363874
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7722
timestamp 1680363874
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7723
timestamp 1680363874
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_463
timestamp 1680363874
transform -1 0 2320 0 -1 1570
box -9 -3 26 105
use BUFX2  BUFX2_75
timestamp 1680363874
transform 1 0 2320 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7724
timestamp 1680363874
transform 1 0 2344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7725
timestamp 1680363874
transform 1 0 2352 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_76
timestamp 1680363874
transform -1 0 2384 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7726
timestamp 1680363874
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7727
timestamp 1680363874
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7728
timestamp 1680363874
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7729
timestamp 1680363874
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_85
timestamp 1680363874
transform 1 0 2416 0 -1 1570
box -8 -3 32 105
use AND2X2  AND2X2_44
timestamp 1680363874
transform 1 0 2440 0 -1 1570
box -8 -3 40 105
use INVX2  INVX2_464
timestamp 1680363874
transform -1 0 2488 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7730
timestamp 1680363874
transform 1 0 2488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7732
timestamp 1680363874
transform 1 0 2496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7734
timestamp 1680363874
transform 1 0 2504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7735
timestamp 1680363874
transform 1 0 2512 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_465
timestamp 1680363874
transform -1 0 2536 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7736
timestamp 1680363874
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7738
timestamp 1680363874
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_466
timestamp 1680363874
transform 1 0 2552 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7743
timestamp 1680363874
transform 1 0 2568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7744
timestamp 1680363874
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7745
timestamp 1680363874
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7746
timestamp 1680363874
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_57
timestamp 1680363874
transform -1 0 2632 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7747
timestamp 1680363874
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7748
timestamp 1680363874
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7754
timestamp 1680363874
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_146
timestamp 1680363874
transform -1 0 2688 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7755
timestamp 1680363874
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7756
timestamp 1680363874
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7757
timestamp 1680363874
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7758
timestamp 1680363874
transform 1 0 2712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7760
timestamp 1680363874
transform 1 0 2720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7762
timestamp 1680363874
transform 1 0 2728 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_60
timestamp 1680363874
transform 1 0 2736 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7766
timestamp 1680363874
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7767
timestamp 1680363874
transform 1 0 2776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7768
timestamp 1680363874
transform 1 0 2784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7770
timestamp 1680363874
transform 1 0 2792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7780
timestamp 1680363874
transform 1 0 2800 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_304
timestamp 1680363874
transform -1 0 2848 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7781
timestamp 1680363874
transform 1 0 2848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7782
timestamp 1680363874
transform 1 0 2856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7783
timestamp 1680363874
transform 1 0 2864 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_468
timestamp 1680363874
transform 1 0 2872 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7784
timestamp 1680363874
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7785
timestamp 1680363874
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7786
timestamp 1680363874
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7787
timestamp 1680363874
transform 1 0 2912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7788
timestamp 1680363874
transform 1 0 2920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7789
timestamp 1680363874
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7790
timestamp 1680363874
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7791
timestamp 1680363874
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_247
timestamp 1680363874
transform 1 0 2952 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7792
timestamp 1680363874
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7793
timestamp 1680363874
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7794
timestamp 1680363874
transform 1 0 3008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7795
timestamp 1680363874
transform 1 0 3016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7796
timestamp 1680363874
transform 1 0 3024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7797
timestamp 1680363874
transform 1 0 3032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7798
timestamp 1680363874
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7799
timestamp 1680363874
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7800
timestamp 1680363874
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7801
timestamp 1680363874
transform 1 0 3064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7802
timestamp 1680363874
transform 1 0 3072 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_248
timestamp 1680363874
transform 1 0 3080 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7803
timestamp 1680363874
transform 1 0 3120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7805
timestamp 1680363874
transform 1 0 3128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7808
timestamp 1680363874
transform 1 0 3136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7809
timestamp 1680363874
transform 1 0 3144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7810
timestamp 1680363874
transform 1 0 3152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7811
timestamp 1680363874
transform 1 0 3160 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_406
timestamp 1680363874
transform -1 0 3264 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7812
timestamp 1680363874
transform 1 0 3264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7813
timestamp 1680363874
transform 1 0 3272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7814
timestamp 1680363874
transform 1 0 3280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7815
timestamp 1680363874
transform 1 0 3288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7817
timestamp 1680363874
transform 1 0 3296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7822
timestamp 1680363874
transform 1 0 3304 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_469
timestamp 1680363874
transform -1 0 3328 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7823
timestamp 1680363874
transform 1 0 3328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7825
timestamp 1680363874
transform 1 0 3336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7826
timestamp 1680363874
transform 1 0 3344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7827
timestamp 1680363874
transform 1 0 3352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7828
timestamp 1680363874
transform 1 0 3360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7829
timestamp 1680363874
transform 1 0 3368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7830
timestamp 1680363874
transform 1 0 3376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7832
timestamp 1680363874
transform 1 0 3384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7834
timestamp 1680363874
transform 1 0 3392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7836
timestamp 1680363874
transform 1 0 3400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7838
timestamp 1680363874
transform 1 0 3408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7843
timestamp 1680363874
transform 1 0 3416 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_305
timestamp 1680363874
transform -1 0 3464 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7844
timestamp 1680363874
transform 1 0 3464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7846
timestamp 1680363874
transform 1 0 3472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7854
timestamp 1680363874
transform 1 0 3480 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_306
timestamp 1680363874
transform -1 0 3528 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7855
timestamp 1680363874
transform 1 0 3528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7857
timestamp 1680363874
transform 1 0 3536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7859
timestamp 1680363874
transform 1 0 3544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7861
timestamp 1680363874
transform 1 0 3552 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_470
timestamp 1680363874
transform 1 0 3560 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_471
timestamp 1680363874
transform 1 0 3576 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_408
timestamp 1680363874
transform -1 0 3688 0 -1 1570
box -8 -3 104 105
use NOR2X1  NOR2X1_87
timestamp 1680363874
transform 1 0 3688 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7876
timestamp 1680363874
transform 1 0 3712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7877
timestamp 1680363874
transform 1 0 3720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7878
timestamp 1680363874
transform 1 0 3728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7879
timestamp 1680363874
transform 1 0 3736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7880
timestamp 1680363874
transform 1 0 3744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7881
timestamp 1680363874
transform 1 0 3752 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_307
timestamp 1680363874
transform -1 0 3800 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7882
timestamp 1680363874
transform 1 0 3800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7886
timestamp 1680363874
transform 1 0 3808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7887
timestamp 1680363874
transform 1 0 3816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7888
timestamp 1680363874
transform 1 0 3824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7889
timestamp 1680363874
transform 1 0 3832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7890
timestamp 1680363874
transform 1 0 3840 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_472
timestamp 1680363874
transform 1 0 3848 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7891
timestamp 1680363874
transform 1 0 3864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7892
timestamp 1680363874
transform 1 0 3872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7893
timestamp 1680363874
transform 1 0 3880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7894
timestamp 1680363874
transform 1 0 3888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7895
timestamp 1680363874
transform 1 0 3896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7896
timestamp 1680363874
transform 1 0 3904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7897
timestamp 1680363874
transform 1 0 3912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7898
timestamp 1680363874
transform 1 0 3920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7899
timestamp 1680363874
transform 1 0 3928 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_88
timestamp 1680363874
transform -1 0 3960 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7900
timestamp 1680363874
transform 1 0 3960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7902
timestamp 1680363874
transform 1 0 3968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7905
timestamp 1680363874
transform 1 0 3976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7906
timestamp 1680363874
transform 1 0 3984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7907
timestamp 1680363874
transform 1 0 3992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7908
timestamp 1680363874
transform 1 0 4000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7909
timestamp 1680363874
transform 1 0 4008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7910
timestamp 1680363874
transform 1 0 4016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7911
timestamp 1680363874
transform 1 0 4024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7912
timestamp 1680363874
transform 1 0 4032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7913
timestamp 1680363874
transform 1 0 4040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7914
timestamp 1680363874
transform 1 0 4048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7915
timestamp 1680363874
transform 1 0 4056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7916
timestamp 1680363874
transform 1 0 4064 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_473
timestamp 1680363874
transform -1 0 4088 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7917
timestamp 1680363874
transform 1 0 4088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7918
timestamp 1680363874
transform 1 0 4096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7919
timestamp 1680363874
transform 1 0 4104 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_252
timestamp 1680363874
transform -1 0 4152 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7920
timestamp 1680363874
transform 1 0 4152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7921
timestamp 1680363874
transform 1 0 4160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7923
timestamp 1680363874
transform 1 0 4168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7925
timestamp 1680363874
transform 1 0 4176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7927
timestamp 1680363874
transform 1 0 4184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7929
timestamp 1680363874
transform 1 0 4192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7930
timestamp 1680363874
transform 1 0 4200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7931
timestamp 1680363874
transform 1 0 4208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7933
timestamp 1680363874
transform 1 0 4216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7935
timestamp 1680363874
transform 1 0 4224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7938
timestamp 1680363874
transform 1 0 4232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7939
timestamp 1680363874
transform 1 0 4240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7940
timestamp 1680363874
transform 1 0 4248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7941
timestamp 1680363874
transform 1 0 4256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7942
timestamp 1680363874
transform 1 0 4264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7943
timestamp 1680363874
transform 1 0 4272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7944
timestamp 1680363874
transform 1 0 4280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7945
timestamp 1680363874
transform 1 0 4288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7946
timestamp 1680363874
transform 1 0 4296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7947
timestamp 1680363874
transform 1 0 4304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7948
timestamp 1680363874
transform 1 0 4312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7949
timestamp 1680363874
transform 1 0 4320 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_310
timestamp 1680363874
transform 1 0 4328 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7950
timestamp 1680363874
transform 1 0 4368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7951
timestamp 1680363874
transform 1 0 4376 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_89
timestamp 1680363874
transform 1 0 4384 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7952
timestamp 1680363874
transform 1 0 4408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7953
timestamp 1680363874
transform 1 0 4416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7954
timestamp 1680363874
transform 1 0 4424 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6240
timestamp 1680363874
transform 1 0 4444 0 1 1475
box -3 -3 3 3
use FILL  FILL_7955
timestamp 1680363874
transform 1 0 4432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7956
timestamp 1680363874
transform 1 0 4440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7957
timestamp 1680363874
transform 1 0 4448 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_311
timestamp 1680363874
transform 1 0 4456 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7966
timestamp 1680363874
transform 1 0 4496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7967
timestamp 1680363874
transform 1 0 4504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7968
timestamp 1680363874
transform 1 0 4512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7969
timestamp 1680363874
transform 1 0 4520 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_90
timestamp 1680363874
transform 1 0 4528 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7970
timestamp 1680363874
transform 1 0 4552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7972
timestamp 1680363874
transform 1 0 4560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7982
timestamp 1680363874
transform 1 0 4568 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_313
timestamp 1680363874
transform -1 0 4616 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7983
timestamp 1680363874
transform 1 0 4616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7984
timestamp 1680363874
transform 1 0 4624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7985
timestamp 1680363874
transform 1 0 4632 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6241
timestamp 1680363874
transform 1 0 4676 0 1 1475
box -3 -3 3 3
use AOI22X1  AOI22X1_254
timestamp 1680363874
transform 1 0 4640 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_476
timestamp 1680363874
transform 1 0 4680 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_414
timestamp 1680363874
transform 1 0 4696 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7986
timestamp 1680363874
transform 1 0 4792 0 -1 1570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_65
timestamp 1680363874
transform 1 0 4851 0 1 1470
box -10 -3 10 3
use M2_M1  M2_M1_6857
timestamp 1680363874
transform 1 0 124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6858
timestamp 1680363874
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6967
timestamp 1680363874
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6292
timestamp 1680363874
transform 1 0 196 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6859
timestamp 1680363874
transform 1 0 188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6968
timestamp 1680363874
transform 1 0 180 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6325
timestamp 1680363874
transform 1 0 196 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6265
timestamp 1680363874
transform 1 0 220 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6860
timestamp 1680363874
transform 1 0 228 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6326
timestamp 1680363874
transform 1 0 236 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6293
timestamp 1680363874
transform 1 0 252 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6861
timestamp 1680363874
transform 1 0 244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6969
timestamp 1680363874
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6970
timestamp 1680363874
transform 1 0 236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6971
timestamp 1680363874
transform 1 0 244 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6398
timestamp 1680363874
transform 1 0 236 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6399
timestamp 1680363874
transform 1 0 260 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6862
timestamp 1680363874
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6327
timestamp 1680363874
transform 1 0 324 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6972
timestamp 1680363874
transform 1 0 324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6863
timestamp 1680363874
transform 1 0 340 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6266
timestamp 1680363874
transform 1 0 380 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6864
timestamp 1680363874
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6973
timestamp 1680363874
transform 1 0 380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6974
timestamp 1680363874
transform 1 0 388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6865
timestamp 1680363874
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6866
timestamp 1680363874
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6867
timestamp 1680363874
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6975
timestamp 1680363874
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6364
timestamp 1680363874
transform 1 0 452 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6868
timestamp 1680363874
transform 1 0 484 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6344
timestamp 1680363874
transform 1 0 492 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7062
timestamp 1680363874
transform 1 0 492 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6267
timestamp 1680363874
transform 1 0 524 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6869
timestamp 1680363874
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6870
timestamp 1680363874
transform 1 0 524 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6345
timestamp 1680363874
transform 1 0 524 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6976
timestamp 1680363874
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6977
timestamp 1680363874
transform 1 0 540 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6365
timestamp 1680363874
transform 1 0 532 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6328
timestamp 1680363874
transform 1 0 548 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6978
timestamp 1680363874
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6366
timestamp 1680363874
transform 1 0 572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6268
timestamp 1680363874
transform 1 0 604 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6871
timestamp 1680363874
transform 1 0 612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6872
timestamp 1680363874
transform 1 0 644 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6979
timestamp 1680363874
transform 1 0 620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6980
timestamp 1680363874
transform 1 0 636 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6367
timestamp 1680363874
transform 1 0 628 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6368
timestamp 1680363874
transform 1 0 652 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6873
timestamp 1680363874
transform 1 0 668 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6346
timestamp 1680363874
transform 1 0 684 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6981
timestamp 1680363874
transform 1 0 692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7063
timestamp 1680363874
transform 1 0 684 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6982
timestamp 1680363874
transform 1 0 724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7064
timestamp 1680363874
transform 1 0 716 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6874
timestamp 1680363874
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6347
timestamp 1680363874
transform 1 0 732 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6294
timestamp 1680363874
transform 1 0 780 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6983
timestamp 1680363874
transform 1 0 780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6984
timestamp 1680363874
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6369
timestamp 1680363874
transform 1 0 788 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6248
timestamp 1680363874
transform 1 0 804 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6269
timestamp 1680363874
transform 1 0 812 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6875
timestamp 1680363874
transform 1 0 804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6876
timestamp 1680363874
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6329
timestamp 1680363874
transform 1 0 836 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6249
timestamp 1680363874
transform 1 0 860 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6985
timestamp 1680363874
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6295
timestamp 1680363874
transform 1 0 876 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6877
timestamp 1680363874
transform 1 0 876 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6330
timestamp 1680363874
transform 1 0 884 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6986
timestamp 1680363874
transform 1 0 884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6987
timestamp 1680363874
transform 1 0 900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6878
timestamp 1680363874
transform 1 0 916 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6348
timestamp 1680363874
transform 1 0 956 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6270
timestamp 1680363874
transform 1 0 988 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6988
timestamp 1680363874
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6271
timestamp 1680363874
transform 1 0 1044 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6296
timestamp 1680363874
transform 1 0 1036 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6331
timestamp 1680363874
transform 1 0 1028 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6879
timestamp 1680363874
transform 1 0 1036 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6880
timestamp 1680363874
transform 1 0 1044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6881
timestamp 1680363874
transform 1 0 1060 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6370
timestamp 1680363874
transform 1 0 1052 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6400
timestamp 1680363874
transform 1 0 1044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6371
timestamp 1680363874
transform 1 0 1100 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6401
timestamp 1680363874
transform 1 0 1092 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6882
timestamp 1680363874
transform 1 0 1116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6851
timestamp 1680363874
transform 1 0 1132 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6297
timestamp 1680363874
transform 1 0 1148 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6883
timestamp 1680363874
transform 1 0 1148 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6332
timestamp 1680363874
transform 1 0 1172 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6989
timestamp 1680363874
transform 1 0 1140 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6990
timestamp 1680363874
transform 1 0 1156 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6349
timestamp 1680363874
transform 1 0 1164 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6991
timestamp 1680363874
transform 1 0 1172 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6372
timestamp 1680363874
transform 1 0 1140 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6884
timestamp 1680363874
transform 1 0 1212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6885
timestamp 1680363874
transform 1 0 1236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6886
timestamp 1680363874
transform 1 0 1252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6992
timestamp 1680363874
transform 1 0 1212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6993
timestamp 1680363874
transform 1 0 1228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6994
timestamp 1680363874
transform 1 0 1244 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6402
timestamp 1680363874
transform 1 0 1212 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6373
timestamp 1680363874
transform 1 0 1244 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6403
timestamp 1680363874
transform 1 0 1252 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6887
timestamp 1680363874
transform 1 0 1308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6995
timestamp 1680363874
transform 1 0 1324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6996
timestamp 1680363874
transform 1 0 1332 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6374
timestamp 1680363874
transform 1 0 1324 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6272
timestamp 1680363874
transform 1 0 1364 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6273
timestamp 1680363874
transform 1 0 1412 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6888
timestamp 1680363874
transform 1 0 1364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6889
timestamp 1680363874
transform 1 0 1372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6890
timestamp 1680363874
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6891
timestamp 1680363874
transform 1 0 1404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6997
timestamp 1680363874
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6998
timestamp 1680363874
transform 1 0 1396 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6333
timestamp 1680363874
transform 1 0 1420 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6892
timestamp 1680363874
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6893
timestamp 1680363874
transform 1 0 1500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6999
timestamp 1680363874
transform 1 0 1420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6375
timestamp 1680363874
transform 1 0 1452 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6298
timestamp 1680363874
transform 1 0 1596 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6334
timestamp 1680363874
transform 1 0 1548 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6894
timestamp 1680363874
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7000
timestamp 1680363874
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6299
timestamp 1680363874
transform 1 0 1692 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6895
timestamp 1680363874
transform 1 0 1684 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7001
timestamp 1680363874
transform 1 0 1692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7002
timestamp 1680363874
transform 1 0 1708 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6274
timestamp 1680363874
transform 1 0 1740 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6896
timestamp 1680363874
transform 1 0 1732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6897
timestamp 1680363874
transform 1 0 1740 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6376
timestamp 1680363874
transform 1 0 1732 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7003
timestamp 1680363874
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6377
timestamp 1680363874
transform 1 0 1756 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7004
timestamp 1680363874
transform 1 0 1772 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6350
timestamp 1680363874
transform 1 0 1804 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6898
timestamp 1680363874
transform 1 0 1876 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6899
timestamp 1680363874
transform 1 0 1908 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6351
timestamp 1680363874
transform 1 0 1908 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7005
timestamp 1680363874
transform 1 0 1956 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6378
timestamp 1680363874
transform 1 0 1956 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6850
timestamp 1680363874
transform 1 0 1996 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_6852
timestamp 1680363874
transform 1 0 1980 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6853
timestamp 1680363874
transform 1 0 2004 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6900
timestamp 1680363874
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6335
timestamp 1680363874
transform 1 0 1996 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6300
timestamp 1680363874
transform 1 0 2100 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6901
timestamp 1680363874
transform 1 0 2100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7006
timestamp 1680363874
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6379
timestamp 1680363874
transform 1 0 2052 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6380
timestamp 1680363874
transform 1 0 2076 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6381
timestamp 1680363874
transform 1 0 2100 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6404
timestamp 1680363874
transform 1 0 2044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6255
timestamp 1680363874
transform 1 0 2140 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_7007
timestamp 1680363874
transform 1 0 2140 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6256
timestamp 1680363874
transform 1 0 2204 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6902
timestamp 1680363874
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6903
timestamp 1680363874
transform 1 0 2172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6904
timestamp 1680363874
transform 1 0 2196 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6405
timestamp 1680363874
transform 1 0 2156 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6352
timestamp 1680363874
transform 1 0 2180 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7008
timestamp 1680363874
transform 1 0 2188 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6353
timestamp 1680363874
transform 1 0 2196 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7009
timestamp 1680363874
transform 1 0 2204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7010
timestamp 1680363874
transform 1 0 2212 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6382
timestamp 1680363874
transform 1 0 2188 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6905
timestamp 1680363874
transform 1 0 2236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7011
timestamp 1680363874
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6301
timestamp 1680363874
transform 1 0 2252 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6302
timestamp 1680363874
transform 1 0 2276 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6906
timestamp 1680363874
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6907
timestamp 1680363874
transform 1 0 2276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7012
timestamp 1680363874
transform 1 0 2268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7013
timestamp 1680363874
transform 1 0 2284 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6275
timestamp 1680363874
transform 1 0 2308 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6908
timestamp 1680363874
transform 1 0 2308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6909
timestamp 1680363874
transform 1 0 2316 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6276
timestamp 1680363874
transform 1 0 2356 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6910
timestamp 1680363874
transform 1 0 2356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6911
timestamp 1680363874
transform 1 0 2380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7014
timestamp 1680363874
transform 1 0 2372 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6383
timestamp 1680363874
transform 1 0 2372 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6336
timestamp 1680363874
transform 1 0 2388 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7015
timestamp 1680363874
transform 1 0 2388 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6303
timestamp 1680363874
transform 1 0 2436 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6912
timestamp 1680363874
transform 1 0 2420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6913
timestamp 1680363874
transform 1 0 2436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7065
timestamp 1680363874
transform 1 0 2412 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6406
timestamp 1680363874
transform 1 0 2412 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6337
timestamp 1680363874
transform 1 0 2444 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6277
timestamp 1680363874
transform 1 0 2468 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6304
timestamp 1680363874
transform 1 0 2468 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6914
timestamp 1680363874
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6915
timestamp 1680363874
transform 1 0 2484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7016
timestamp 1680363874
transform 1 0 2444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7017
timestamp 1680363874
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7018
timestamp 1680363874
transform 1 0 2460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6384
timestamp 1680363874
transform 1 0 2452 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6354
timestamp 1680363874
transform 1 0 2468 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6305
timestamp 1680363874
transform 1 0 2508 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6916
timestamp 1680363874
transform 1 0 2500 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6338
timestamp 1680363874
transform 1 0 2540 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6917
timestamp 1680363874
transform 1 0 2556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7019
timestamp 1680363874
transform 1 0 2580 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6385
timestamp 1680363874
transform 1 0 2580 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6250
timestamp 1680363874
transform 1 0 2620 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6257
timestamp 1680363874
transform 1 0 2604 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6258
timestamp 1680363874
transform 1 0 2660 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6306
timestamp 1680363874
transform 1 0 2636 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6918
timestamp 1680363874
transform 1 0 2636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6919
timestamp 1680363874
transform 1 0 2692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6920
timestamp 1680363874
transform 1 0 2700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7020
timestamp 1680363874
transform 1 0 2612 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6355
timestamp 1680363874
transform 1 0 2652 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6386
timestamp 1680363874
transform 1 0 2612 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7021
timestamp 1680363874
transform 1 0 2708 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6339
timestamp 1680363874
transform 1 0 2740 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7022
timestamp 1680363874
transform 1 0 2740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7023
timestamp 1680363874
transform 1 0 2756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6356
timestamp 1680363874
transform 1 0 2788 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7066
timestamp 1680363874
transform 1 0 2788 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6278
timestamp 1680363874
transform 1 0 2804 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6921
timestamp 1680363874
transform 1 0 2804 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6357
timestamp 1680363874
transform 1 0 2828 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6358
timestamp 1680363874
transform 1 0 2844 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6307
timestamp 1680363874
transform 1 0 2868 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6308
timestamp 1680363874
transform 1 0 2908 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6922
timestamp 1680363874
transform 1 0 2884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6923
timestamp 1680363874
transform 1 0 2900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7024
timestamp 1680363874
transform 1 0 2876 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6359
timestamp 1680363874
transform 1 0 2884 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7025
timestamp 1680363874
transform 1 0 2892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7026
timestamp 1680363874
transform 1 0 2908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7027
timestamp 1680363874
transform 1 0 2916 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6924
timestamp 1680363874
transform 1 0 2972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6854
timestamp 1680363874
transform 1 0 2988 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6925
timestamp 1680363874
transform 1 0 3044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7028
timestamp 1680363874
transform 1 0 3068 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6309
timestamp 1680363874
transform 1 0 3100 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6340
timestamp 1680363874
transform 1 0 3092 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6926
timestamp 1680363874
transform 1 0 3100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6927
timestamp 1680363874
transform 1 0 3116 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6310
timestamp 1680363874
transform 1 0 3132 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_7029
timestamp 1680363874
transform 1 0 3108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7030
timestamp 1680363874
transform 1 0 3124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7031
timestamp 1680363874
transform 1 0 3132 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6407
timestamp 1680363874
transform 1 0 3108 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6259
timestamp 1680363874
transform 1 0 3172 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6341
timestamp 1680363874
transform 1 0 3188 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7032
timestamp 1680363874
transform 1 0 3188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6928
timestamp 1680363874
transform 1 0 3204 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6279
timestamp 1680363874
transform 1 0 3220 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6929
timestamp 1680363874
transform 1 0 3236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6930
timestamp 1680363874
transform 1 0 3252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7033
timestamp 1680363874
transform 1 0 3260 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6280
timestamp 1680363874
transform 1 0 3276 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6931
timestamp 1680363874
transform 1 0 3276 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6311
timestamp 1680363874
transform 1 0 3284 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_7034
timestamp 1680363874
transform 1 0 3292 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6360
timestamp 1680363874
transform 1 0 3300 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6281
timestamp 1680363874
transform 1 0 3332 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6312
timestamp 1680363874
transform 1 0 3372 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6932
timestamp 1680363874
transform 1 0 3332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6933
timestamp 1680363874
transform 1 0 3348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6934
timestamp 1680363874
transform 1 0 3364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7035
timestamp 1680363874
transform 1 0 3340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7036
timestamp 1680363874
transform 1 0 3356 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6361
timestamp 1680363874
transform 1 0 3364 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7037
timestamp 1680363874
transform 1 0 3372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6855
timestamp 1680363874
transform 1 0 3404 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6260
timestamp 1680363874
transform 1 0 3452 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6856
timestamp 1680363874
transform 1 0 3444 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6935
timestamp 1680363874
transform 1 0 3452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7038
timestamp 1680363874
transform 1 0 3444 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6242
timestamp 1680363874
transform 1 0 3476 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6251
timestamp 1680363874
transform 1 0 3476 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6243
timestamp 1680363874
transform 1 0 3492 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6387
timestamp 1680363874
transform 1 0 3484 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6282
timestamp 1680363874
transform 1 0 3516 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6936
timestamp 1680363874
transform 1 0 3508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6937
timestamp 1680363874
transform 1 0 3516 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6252
timestamp 1680363874
transform 1 0 3540 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6261
timestamp 1680363874
transform 1 0 3564 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6938
timestamp 1680363874
transform 1 0 3548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6939
timestamp 1680363874
transform 1 0 3564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7039
timestamp 1680363874
transform 1 0 3540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7040
timestamp 1680363874
transform 1 0 3556 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6388
timestamp 1680363874
transform 1 0 3556 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6408
timestamp 1680363874
transform 1 0 3540 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6313
timestamp 1680363874
transform 1 0 3580 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6283
timestamp 1680363874
transform 1 0 3652 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6314
timestamp 1680363874
transform 1 0 3636 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6940
timestamp 1680363874
transform 1 0 3636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7041
timestamp 1680363874
transform 1 0 3684 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6389
timestamp 1680363874
transform 1 0 3684 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6409
timestamp 1680363874
transform 1 0 3612 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6941
timestamp 1680363874
transform 1 0 3708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7042
timestamp 1680363874
transform 1 0 3700 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6410
timestamp 1680363874
transform 1 0 3700 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6362
timestamp 1680363874
transform 1 0 3716 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6244
timestamp 1680363874
transform 1 0 3764 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6253
timestamp 1680363874
transform 1 0 3772 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6262
timestamp 1680363874
transform 1 0 3764 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6284
timestamp 1680363874
transform 1 0 3756 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6942
timestamp 1680363874
transform 1 0 3748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6943
timestamp 1680363874
transform 1 0 3764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7043
timestamp 1680363874
transform 1 0 3756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7044
timestamp 1680363874
transform 1 0 3764 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6263
timestamp 1680363874
transform 1 0 3788 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6285
timestamp 1680363874
transform 1 0 3796 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6264
timestamp 1680363874
transform 1 0 3820 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6286
timestamp 1680363874
transform 1 0 3828 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6315
timestamp 1680363874
transform 1 0 3820 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6254
timestamp 1680363874
transform 1 0 3916 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6316
timestamp 1680363874
transform 1 0 3860 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6944
timestamp 1680363874
transform 1 0 3820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6945
timestamp 1680363874
transform 1 0 3828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6946
timestamp 1680363874
transform 1 0 3860 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6363
timestamp 1680363874
transform 1 0 3820 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7045
timestamp 1680363874
transform 1 0 3908 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6390
timestamp 1680363874
transform 1 0 3908 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6947
timestamp 1680363874
transform 1 0 3948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7046
timestamp 1680363874
transform 1 0 3940 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6411
timestamp 1680363874
transform 1 0 3940 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6245
timestamp 1680363874
transform 1 0 3988 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6287
timestamp 1680363874
transform 1 0 3980 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6948
timestamp 1680363874
transform 1 0 3972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6949
timestamp 1680363874
transform 1 0 3988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7047
timestamp 1680363874
transform 1 0 3980 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6246
timestamp 1680363874
transform 1 0 4084 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6288
timestamp 1680363874
transform 1 0 4020 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6950
timestamp 1680363874
transform 1 0 4060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7048
timestamp 1680363874
transform 1 0 4028 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6391
timestamp 1680363874
transform 1 0 4028 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6392
timestamp 1680363874
transform 1 0 4060 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6951
timestamp 1680363874
transform 1 0 4124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7067
timestamp 1680363874
transform 1 0 4148 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6412
timestamp 1680363874
transform 1 0 4140 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6247
timestamp 1680363874
transform 1 0 4180 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6289
timestamp 1680363874
transform 1 0 4180 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6952
timestamp 1680363874
transform 1 0 4172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6953
timestamp 1680363874
transform 1 0 4180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7049
timestamp 1680363874
transform 1 0 4164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7050
timestamp 1680363874
transform 1 0 4180 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6413
timestamp 1680363874
transform 1 0 4180 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6317
timestamp 1680363874
transform 1 0 4228 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_7051
timestamp 1680363874
transform 1 0 4228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6393
timestamp 1680363874
transform 1 0 4244 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6290
timestamp 1680363874
transform 1 0 4292 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6318
timestamp 1680363874
transform 1 0 4276 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6954
timestamp 1680363874
transform 1 0 4252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6955
timestamp 1680363874
transform 1 0 4260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6956
timestamp 1680363874
transform 1 0 4276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6957
timestamp 1680363874
transform 1 0 4292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7052
timestamp 1680363874
transform 1 0 4252 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6394
timestamp 1680363874
transform 1 0 4260 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6414
timestamp 1680363874
transform 1 0 4252 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_7053
timestamp 1680363874
transform 1 0 4300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7054
timestamp 1680363874
transform 1 0 4316 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6319
timestamp 1680363874
transform 1 0 4340 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6320
timestamp 1680363874
transform 1 0 4380 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6395
timestamp 1680363874
transform 1 0 4380 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6291
timestamp 1680363874
transform 1 0 4444 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_7068
timestamp 1680363874
transform 1 0 4460 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6342
timestamp 1680363874
transform 1 0 4476 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7055
timestamp 1680363874
transform 1 0 4492 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6321
timestamp 1680363874
transform 1 0 4508 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6958
timestamp 1680363874
transform 1 0 4500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6959
timestamp 1680363874
transform 1 0 4508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6960
timestamp 1680363874
transform 1 0 4524 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6343
timestamp 1680363874
transform 1 0 4532 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6322
timestamp 1680363874
transform 1 0 4548 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6961
timestamp 1680363874
transform 1 0 4540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6962
timestamp 1680363874
transform 1 0 4548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7056
timestamp 1680363874
transform 1 0 4508 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7057
timestamp 1680363874
transform 1 0 4540 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6396
timestamp 1680363874
transform 1 0 4532 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6415
timestamp 1680363874
transform 1 0 4540 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6963
timestamp 1680363874
transform 1 0 4596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7058
timestamp 1680363874
transform 1 0 4572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7059
timestamp 1680363874
transform 1 0 4580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7060
timestamp 1680363874
transform 1 0 4604 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6397
timestamp 1680363874
transform 1 0 4596 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6416
timestamp 1680363874
transform 1 0 4588 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6417
timestamp 1680363874
transform 1 0 4604 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6848
timestamp 1680363874
transform 1 0 4620 0 1 1455
box -2 -2 2 2
use M2_M1  M2_M1_6964
timestamp 1680363874
transform 1 0 4636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1680363874
transform 1 0 4676 0 1 1455
box -2 -2 2 2
use M3_M2  M3_M2_6323
timestamp 1680363874
transform 1 0 4676 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6324
timestamp 1680363874
transform 1 0 4796 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6965
timestamp 1680363874
transform 1 0 4740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6966
timestamp 1680363874
transform 1 0 4796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7061
timestamp 1680363874
transform 1 0 4716 0 1 1405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_66
timestamp 1680363874
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_7987
timestamp 1680363874
transform 1 0 72 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_415
timestamp 1680363874
transform 1 0 80 0 1 1370
box -8 -3 104 105
use FILL  FILL_7989
timestamp 1680363874
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_7990
timestamp 1680363874
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_7991
timestamp 1680363874
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_7992
timestamp 1680363874
transform 1 0 200 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6418
timestamp 1680363874
transform 1 0 228 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_255
timestamp 1680363874
transform 1 0 208 0 1 1370
box -8 -3 46 105
use FILL  FILL_7993
timestamp 1680363874
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_7994
timestamp 1680363874
transform 1 0 256 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_477
timestamp 1680363874
transform 1 0 264 0 1 1370
box -9 -3 26 105
use FILL  FILL_7995
timestamp 1680363874
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_7996
timestamp 1680363874
transform 1 0 288 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6419
timestamp 1680363874
transform 1 0 308 0 1 1375
box -3 -3 3 3
use FILL  FILL_7997
timestamp 1680363874
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_7998
timestamp 1680363874
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_7999
timestamp 1680363874
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8000
timestamp 1680363874
transform 1 0 320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8001
timestamp 1680363874
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8012
timestamp 1680363874
transform 1 0 336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8014
timestamp 1680363874
transform 1 0 344 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_256
timestamp 1680363874
transform -1 0 392 0 1 1370
box -8 -3 46 105
use FILL  FILL_8015
timestamp 1680363874
transform 1 0 392 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_479
timestamp 1680363874
transform 1 0 400 0 1 1370
box -9 -3 26 105
use FILL  FILL_8019
timestamp 1680363874
transform 1 0 416 0 1 1370
box -8 -3 16 105
use FILL  FILL_8020
timestamp 1680363874
transform 1 0 424 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_16
timestamp 1680363874
transform -1 0 464 0 1 1370
box -7 -3 39 105
use FILL  FILL_8021
timestamp 1680363874
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_8022
timestamp 1680363874
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_8023
timestamp 1680363874
transform 1 0 480 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_17
timestamp 1680363874
transform -1 0 520 0 1 1370
box -7 -3 39 105
use FILL  FILL_8024
timestamp 1680363874
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_8025
timestamp 1680363874
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_8026
timestamp 1680363874
transform 1 0 536 0 1 1370
box -8 -3 16 105
use FILL  FILL_8027
timestamp 1680363874
transform 1 0 544 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_480
timestamp 1680363874
transform 1 0 552 0 1 1370
box -9 -3 26 105
use FILL  FILL_8028
timestamp 1680363874
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_8033
timestamp 1680363874
transform 1 0 576 0 1 1370
box -8 -3 16 105
use FILL  FILL_8035
timestamp 1680363874
transform 1 0 584 0 1 1370
box -8 -3 16 105
use FILL  FILL_8037
timestamp 1680363874
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_8039
timestamp 1680363874
transform 1 0 600 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_18
timestamp 1680363874
transform 1 0 608 0 1 1370
box -7 -3 39 105
use FILL  FILL_8040
timestamp 1680363874
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_8043
timestamp 1680363874
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_8045
timestamp 1680363874
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_8047
timestamp 1680363874
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_8049
timestamp 1680363874
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_8051
timestamp 1680363874
transform 1 0 680 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_19
timestamp 1680363874
transform 1 0 688 0 1 1370
box -7 -3 39 105
use FILL  FILL_8052
timestamp 1680363874
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_8055
timestamp 1680363874
transform 1 0 728 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_481
timestamp 1680363874
transform -1 0 752 0 1 1370
box -9 -3 26 105
use FILL  FILL_8056
timestamp 1680363874
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_8057
timestamp 1680363874
transform 1 0 760 0 1 1370
box -8 -3 16 105
use FILL  FILL_8058
timestamp 1680363874
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8063
timestamp 1680363874
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8065
timestamp 1680363874
transform 1 0 784 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_483
timestamp 1680363874
transform 1 0 792 0 1 1370
box -9 -3 26 105
use FILL  FILL_8067
timestamp 1680363874
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_8071
timestamp 1680363874
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_8073
timestamp 1680363874
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_8075
timestamp 1680363874
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_8077
timestamp 1680363874
transform 1 0 840 0 1 1370
box -8 -3 16 105
use FILL  FILL_8078
timestamp 1680363874
transform 1 0 848 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_257
timestamp 1680363874
transform 1 0 856 0 1 1370
box -8 -3 46 105
use FILL  FILL_8079
timestamp 1680363874
transform 1 0 896 0 1 1370
box -8 -3 16 105
use FILL  FILL_8083
timestamp 1680363874
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_8085
timestamp 1680363874
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_8087
timestamp 1680363874
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8089
timestamp 1680363874
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_8091
timestamp 1680363874
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_8093
timestamp 1680363874
transform 1 0 944 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_484
timestamp 1680363874
transform 1 0 952 0 1 1370
box -9 -3 26 105
use FILL  FILL_8095
timestamp 1680363874
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8099
timestamp 1680363874
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8101
timestamp 1680363874
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_8103
timestamp 1680363874
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_8104
timestamp 1680363874
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FILL  FILL_8105
timestamp 1680363874
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8107
timestamp 1680363874
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_8109
timestamp 1680363874
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8111
timestamp 1680363874
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_259
timestamp 1680363874
transform 1 0 1040 0 1 1370
box -8 -3 46 105
use FILL  FILL_8113
timestamp 1680363874
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_8114
timestamp 1680363874
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_8117
timestamp 1680363874
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_8119
timestamp 1680363874
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_8121
timestamp 1680363874
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8123
timestamp 1680363874
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_8125
timestamp 1680363874
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_315
timestamp 1680363874
transform -1 0 1176 0 1 1370
box -8 -3 46 105
use FILL  FILL_8126
timestamp 1680363874
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_8129
timestamp 1680363874
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_8131
timestamp 1680363874
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8133
timestamp 1680363874
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_316
timestamp 1680363874
transform 1 0 1208 0 1 1370
box -8 -3 46 105
use FILL  FILL_8135
timestamp 1680363874
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_486
timestamp 1680363874
transform -1 0 1272 0 1 1370
box -9 -3 26 105
use FILL  FILL_8136
timestamp 1680363874
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_8137
timestamp 1680363874
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_8138
timestamp 1680363874
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_8139
timestamp 1680363874
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_8140
timestamp 1680363874
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8141
timestamp 1680363874
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8149
timestamp 1680363874
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_81
timestamp 1680363874
transform -1 0 1352 0 1 1370
box -5 -3 28 105
use FILL  FILL_8150
timestamp 1680363874
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8151
timestamp 1680363874
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_262
timestamp 1680363874
transform 1 0 1368 0 1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_416
timestamp 1680363874
transform 1 0 1408 0 1 1370
box -8 -3 104 105
use FILL  FILL_8152
timestamp 1680363874
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_8153
timestamp 1680363874
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_8154
timestamp 1680363874
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_8165
timestamp 1680363874
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_418
timestamp 1680363874
transform 1 0 1536 0 1 1370
box -8 -3 104 105
use FILL  FILL_8167
timestamp 1680363874
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_8168
timestamp 1680363874
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_8169
timestamp 1680363874
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_490
timestamp 1680363874
transform 1 0 1656 0 1 1370
box -9 -3 26 105
use FILL  FILL_8170
timestamp 1680363874
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_8171
timestamp 1680363874
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8172
timestamp 1680363874
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_8173
timestamp 1680363874
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_8174
timestamp 1680363874
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_82
timestamp 1680363874
transform -1 0 1736 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_83
timestamp 1680363874
transform 1 0 1736 0 1 1370
box -5 -3 28 105
use FILL  FILL_8175
timestamp 1680363874
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_8188
timestamp 1680363874
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8190
timestamp 1680363874
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8192
timestamp 1680363874
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_8193
timestamp 1680363874
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_8194
timestamp 1680363874
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use FILL  FILL_8195
timestamp 1680363874
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_8196
timestamp 1680363874
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_8197
timestamp 1680363874
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_8199
timestamp 1680363874
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_8201
timestamp 1680363874
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_8203
timestamp 1680363874
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_8205
timestamp 1680363874
transform 1 0 1856 0 1 1370
box -8 -3 16 105
use FILL  FILL_8206
timestamp 1680363874
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_420
timestamp 1680363874
transform -1 0 1968 0 1 1370
box -8 -3 104 105
use FILL  FILL_8207
timestamp 1680363874
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_61
timestamp 1680363874
transform 1 0 1976 0 1 1370
box -8 -3 40 105
use FILL  FILL_8208
timestamp 1680363874
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8209
timestamp 1680363874
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_8222
timestamp 1680363874
transform 1 0 2024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8224
timestamp 1680363874
transform 1 0 2032 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_421
timestamp 1680363874
transform 1 0 2040 0 1 1370
box -8 -3 104 105
use FILL  FILL_8226
timestamp 1680363874
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_8227
timestamp 1680363874
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_8228
timestamp 1680363874
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_8229
timestamp 1680363874
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_318
timestamp 1680363874
transform 1 0 2168 0 1 1370
box -8 -3 46 105
use FILL  FILL_8230
timestamp 1680363874
transform 1 0 2208 0 1 1370
box -8 -3 16 105
use FILL  FILL_8241
timestamp 1680363874
transform 1 0 2216 0 1 1370
box -8 -3 16 105
use FILL  FILL_8242
timestamp 1680363874
transform 1 0 2224 0 1 1370
box -8 -3 16 105
use FILL  FILL_8243
timestamp 1680363874
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_266
timestamp 1680363874
transform 1 0 2240 0 1 1370
box -8 -3 46 105
use FILL  FILL_8245
timestamp 1680363874
transform 1 0 2280 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_84
timestamp 1680363874
transform -1 0 2312 0 1 1370
box -5 -3 28 105
use FILL  FILL_8246
timestamp 1680363874
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8253
timestamp 1680363874
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8254
timestamp 1680363874
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_50
timestamp 1680363874
transform -1 0 2368 0 1 1370
box -8 -3 40 105
use FILL  FILL_8255
timestamp 1680363874
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_94
timestamp 1680363874
transform -1 0 2400 0 1 1370
box -8 -3 32 105
use FILL  FILL_8256
timestamp 1680363874
transform 1 0 2400 0 1 1370
box -8 -3 16 105
use FILL  FILL_8257
timestamp 1680363874
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_51
timestamp 1680363874
transform -1 0 2448 0 1 1370
box -8 -3 40 105
use FILL  FILL_8258
timestamp 1680363874
transform 1 0 2448 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_52
timestamp 1680363874
transform 1 0 2456 0 1 1370
box -8 -3 40 105
use FILL  FILL_8259
timestamp 1680363874
transform 1 0 2488 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_422
timestamp 1680363874
transform -1 0 2592 0 1 1370
box -8 -3 104 105
use FILL  FILL_8260
timestamp 1680363874
transform 1 0 2592 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_423
timestamp 1680363874
transform 1 0 2600 0 1 1370
box -8 -3 104 105
use FILL  FILL_8279
timestamp 1680363874
transform 1 0 2696 0 1 1370
box -8 -3 16 105
use FILL  FILL_8280
timestamp 1680363874
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_8288
timestamp 1680363874
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_97
timestamp 1680363874
transform -1 0 2744 0 1 1370
box -8 -3 32 105
use FILL  FILL_8289
timestamp 1680363874
transform 1 0 2744 0 1 1370
box -8 -3 16 105
use FILL  FILL_8290
timestamp 1680363874
transform 1 0 2752 0 1 1370
box -8 -3 16 105
use FILL  FILL_8291
timestamp 1680363874
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FILL  FILL_8292
timestamp 1680363874
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8293
timestamp 1680363874
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8294
timestamp 1680363874
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_53
timestamp 1680363874
transform 1 0 2792 0 1 1370
box -8 -3 40 105
use FILL  FILL_8295
timestamp 1680363874
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_8299
timestamp 1680363874
transform 1 0 2832 0 1 1370
box -8 -3 16 105
use FILL  FILL_8301
timestamp 1680363874
transform 1 0 2840 0 1 1370
box -8 -3 16 105
use FILL  FILL_8302
timestamp 1680363874
transform 1 0 2848 0 1 1370
box -8 -3 16 105
use FILL  FILL_8303
timestamp 1680363874
transform 1 0 2856 0 1 1370
box -8 -3 16 105
use FILL  FILL_8305
timestamp 1680363874
transform 1 0 2864 0 1 1370
box -8 -3 16 105
use FILL  FILL_8307
timestamp 1680363874
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_269
timestamp 1680363874
transform 1 0 2880 0 1 1370
box -8 -3 46 105
use FILL  FILL_8309
timestamp 1680363874
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8314
timestamp 1680363874
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_8315
timestamp 1680363874
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_8316
timestamp 1680363874
transform 1 0 2944 0 1 1370
box -8 -3 16 105
use FILL  FILL_8317
timestamp 1680363874
transform 1 0 2952 0 1 1370
box -8 -3 16 105
use FILL  FILL_8318
timestamp 1680363874
transform 1 0 2960 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6420
timestamp 1680363874
transform 1 0 2980 0 1 1375
box -3 -3 3 3
use FILL  FILL_8319
timestamp 1680363874
transform 1 0 2968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8320
timestamp 1680363874
transform 1 0 2976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8321
timestamp 1680363874
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_8322
timestamp 1680363874
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_8323
timestamp 1680363874
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_8324
timestamp 1680363874
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8326
timestamp 1680363874
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_499
timestamp 1680363874
transform 1 0 3024 0 1 1370
box -9 -3 26 105
use FILL  FILL_8328
timestamp 1680363874
transform 1 0 3040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8332
timestamp 1680363874
transform 1 0 3048 0 1 1370
box -8 -3 16 105
use FILL  FILL_8333
timestamp 1680363874
transform 1 0 3056 0 1 1370
box -8 -3 16 105
use FILL  FILL_8334
timestamp 1680363874
transform 1 0 3064 0 1 1370
box -8 -3 16 105
use FILL  FILL_8335
timestamp 1680363874
transform 1 0 3072 0 1 1370
box -8 -3 16 105
use FILL  FILL_8336
timestamp 1680363874
transform 1 0 3080 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6421
timestamp 1680363874
transform 1 0 3116 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_321
timestamp 1680363874
transform -1 0 3128 0 1 1370
box -8 -3 46 105
use FILL  FILL_8337
timestamp 1680363874
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8338
timestamp 1680363874
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_8339
timestamp 1680363874
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_8340
timestamp 1680363874
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use FILL  FILL_8341
timestamp 1680363874
transform 1 0 3160 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_501
timestamp 1680363874
transform 1 0 3168 0 1 1370
box -9 -3 26 105
use FILL  FILL_8343
timestamp 1680363874
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_8344
timestamp 1680363874
transform 1 0 3192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8345
timestamp 1680363874
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6422
timestamp 1680363874
transform 1 0 3220 0 1 1375
box -3 -3 3 3
use FILL  FILL_8346
timestamp 1680363874
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_8347
timestamp 1680363874
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use FILL  FILL_8348
timestamp 1680363874
transform 1 0 3224 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_271
timestamp 1680363874
transform 1 0 3232 0 1 1370
box -8 -3 46 105
use FILL  FILL_8349
timestamp 1680363874
transform 1 0 3272 0 1 1370
box -8 -3 16 105
use FILL  FILL_8350
timestamp 1680363874
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use FILL  FILL_8351
timestamp 1680363874
transform 1 0 3288 0 1 1370
box -8 -3 16 105
use FILL  FILL_8352
timestamp 1680363874
transform 1 0 3296 0 1 1370
box -8 -3 16 105
use FILL  FILL_8353
timestamp 1680363874
transform 1 0 3304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8354
timestamp 1680363874
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8355
timestamp 1680363874
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_272
timestamp 1680363874
transform 1 0 3328 0 1 1370
box -8 -3 46 105
use FILL  FILL_8356
timestamp 1680363874
transform 1 0 3368 0 1 1370
box -8 -3 16 105
use FILL  FILL_8357
timestamp 1680363874
transform 1 0 3376 0 1 1370
box -8 -3 16 105
use FILL  FILL_8366
timestamp 1680363874
transform 1 0 3384 0 1 1370
box -8 -3 16 105
use FILL  FILL_8368
timestamp 1680363874
transform 1 0 3392 0 1 1370
box -8 -3 16 105
use FILL  FILL_8370
timestamp 1680363874
transform 1 0 3400 0 1 1370
box -8 -3 16 105
use FILL  FILL_8371
timestamp 1680363874
transform 1 0 3408 0 1 1370
box -8 -3 16 105
use FILL  FILL_8372
timestamp 1680363874
transform 1 0 3416 0 1 1370
box -8 -3 16 105
use FILL  FILL_8373
timestamp 1680363874
transform 1 0 3424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8375
timestamp 1680363874
transform 1 0 3432 0 1 1370
box -8 -3 16 105
use AND2X2  AND2X2_54
timestamp 1680363874
transform 1 0 3440 0 1 1370
box -8 -3 40 105
use FILL  FILL_8377
timestamp 1680363874
transform 1 0 3472 0 1 1370
box -8 -3 16 105
use FILL  FILL_8383
timestamp 1680363874
transform 1 0 3480 0 1 1370
box -8 -3 16 105
use FILL  FILL_8385
timestamp 1680363874
transform 1 0 3488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8386
timestamp 1680363874
transform 1 0 3496 0 1 1370
box -8 -3 16 105
use FILL  FILL_8387
timestamp 1680363874
transform 1 0 3504 0 1 1370
box -8 -3 16 105
use FILL  FILL_8388
timestamp 1680363874
transform 1 0 3512 0 1 1370
box -8 -3 16 105
use FILL  FILL_8389
timestamp 1680363874
transform 1 0 3520 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_273
timestamp 1680363874
transform 1 0 3528 0 1 1370
box -8 -3 46 105
use FILL  FILL_8391
timestamp 1680363874
transform 1 0 3568 0 1 1370
box -8 -3 16 105
use FILL  FILL_8392
timestamp 1680363874
transform 1 0 3576 0 1 1370
box -8 -3 16 105
use FILL  FILL_8393
timestamp 1680363874
transform 1 0 3584 0 1 1370
box -8 -3 16 105
use FILL  FILL_8398
timestamp 1680363874
transform 1 0 3592 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_427
timestamp 1680363874
transform -1 0 3696 0 1 1370
box -8 -3 104 105
use FILL  FILL_8399
timestamp 1680363874
transform 1 0 3696 0 1 1370
box -8 -3 16 105
use FILL  FILL_8400
timestamp 1680363874
transform 1 0 3704 0 1 1370
box -8 -3 16 105
use FILL  FILL_8401
timestamp 1680363874
transform 1 0 3712 0 1 1370
box -8 -3 16 105
use FILL  FILL_8402
timestamp 1680363874
transform 1 0 3720 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_274
timestamp 1680363874
transform 1 0 3728 0 1 1370
box -8 -3 46 105
use FILL  FILL_8403
timestamp 1680363874
transform 1 0 3768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8412
timestamp 1680363874
transform 1 0 3776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8414
timestamp 1680363874
transform 1 0 3784 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_503
timestamp 1680363874
transform 1 0 3792 0 1 1370
box -9 -3 26 105
use FILL  FILL_8415
timestamp 1680363874
transform 1 0 3808 0 1 1370
box -8 -3 16 105
use FILL  FILL_8416
timestamp 1680363874
transform 1 0 3816 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_429
timestamp 1680363874
transform -1 0 3920 0 1 1370
box -8 -3 104 105
use FILL  FILL_8417
timestamp 1680363874
transform 1 0 3920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8422
timestamp 1680363874
transform 1 0 3928 0 1 1370
box -8 -3 16 105
use FILL  FILL_8424
timestamp 1680363874
transform 1 0 3936 0 1 1370
box -8 -3 16 105
use FILL  FILL_8426
timestamp 1680363874
transform 1 0 3944 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_275
timestamp 1680363874
transform 1 0 3952 0 1 1370
box -8 -3 46 105
use FILL  FILL_8427
timestamp 1680363874
transform 1 0 3992 0 1 1370
box -8 -3 16 105
use FILL  FILL_8428
timestamp 1680363874
transform 1 0 4000 0 1 1370
box -8 -3 16 105
use FILL  FILL_8429
timestamp 1680363874
transform 1 0 4008 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_431
timestamp 1680363874
transform 1 0 4016 0 1 1370
box -8 -3 104 105
use FILL  FILL_8430
timestamp 1680363874
transform 1 0 4112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8431
timestamp 1680363874
transform 1 0 4120 0 1 1370
box -8 -3 16 105
use FILL  FILL_8432
timestamp 1680363874
transform 1 0 4128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8433
timestamp 1680363874
transform 1 0 4136 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_99
timestamp 1680363874
transform 1 0 4144 0 1 1370
box -8 -3 32 105
use FILL  FILL_8434
timestamp 1680363874
transform 1 0 4168 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_505
timestamp 1680363874
transform 1 0 4176 0 1 1370
box -9 -3 26 105
use FILL  FILL_8435
timestamp 1680363874
transform 1 0 4192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8436
timestamp 1680363874
transform 1 0 4200 0 1 1370
box -8 -3 16 105
use FILL  FILL_8437
timestamp 1680363874
transform 1 0 4208 0 1 1370
box -8 -3 16 105
use FILL  FILL_8438
timestamp 1680363874
transform 1 0 4216 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_506
timestamp 1680363874
transform 1 0 4224 0 1 1370
box -9 -3 26 105
use FILL  FILL_8439
timestamp 1680363874
transform 1 0 4240 0 1 1370
box -8 -3 16 105
use FILL  FILL_8440
timestamp 1680363874
transform 1 0 4248 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_276
timestamp 1680363874
transform 1 0 4256 0 1 1370
box -8 -3 46 105
use FILL  FILL_8441
timestamp 1680363874
transform 1 0 4296 0 1 1370
box -8 -3 16 105
use FILL  FILL_8442
timestamp 1680363874
transform 1 0 4304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8443
timestamp 1680363874
transform 1 0 4312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8444
timestamp 1680363874
transform 1 0 4320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8453
timestamp 1680363874
transform 1 0 4328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8455
timestamp 1680363874
transform 1 0 4336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8456
timestamp 1680363874
transform 1 0 4344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8457
timestamp 1680363874
transform 1 0 4352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8458
timestamp 1680363874
transform 1 0 4360 0 1 1370
box -8 -3 16 105
use FILL  FILL_8459
timestamp 1680363874
transform 1 0 4368 0 1 1370
box -8 -3 16 105
use FILL  FILL_8460
timestamp 1680363874
transform 1 0 4376 0 1 1370
box -8 -3 16 105
use FILL  FILL_8461
timestamp 1680363874
transform 1 0 4384 0 1 1370
box -8 -3 16 105
use FILL  FILL_8464
timestamp 1680363874
transform 1 0 4392 0 1 1370
box -8 -3 16 105
use FILL  FILL_8466
timestamp 1680363874
transform 1 0 4400 0 1 1370
box -8 -3 16 105
use FILL  FILL_8468
timestamp 1680363874
transform 1 0 4408 0 1 1370
box -8 -3 16 105
use FILL  FILL_8470
timestamp 1680363874
transform 1 0 4416 0 1 1370
box -8 -3 16 105
use FILL  FILL_8471
timestamp 1680363874
transform 1 0 4424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8472
timestamp 1680363874
transform 1 0 4432 0 1 1370
box -8 -3 16 105
use FILL  FILL_8473
timestamp 1680363874
transform 1 0 4440 0 1 1370
box -8 -3 16 105
use FILL  FILL_8474
timestamp 1680363874
transform 1 0 4448 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_100
timestamp 1680363874
transform 1 0 4456 0 1 1370
box -8 -3 32 105
use FILL  FILL_8475
timestamp 1680363874
transform 1 0 4480 0 1 1370
box -8 -3 16 105
use FILL  FILL_8476
timestamp 1680363874
transform 1 0 4488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8477
timestamp 1680363874
transform 1 0 4496 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_278
timestamp 1680363874
transform -1 0 4544 0 1 1370
box -8 -3 46 105
use FILL  FILL_8478
timestamp 1680363874
transform 1 0 4544 0 1 1370
box -8 -3 16 105
use FILL  FILL_8479
timestamp 1680363874
transform 1 0 4552 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6423
timestamp 1680363874
transform 1 0 4572 0 1 1375
box -3 -3 3 3
use FILL  FILL_8482
timestamp 1680363874
transform 1 0 4560 0 1 1370
box -8 -3 16 105
use FILL  FILL_8484
timestamp 1680363874
transform 1 0 4568 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_279
timestamp 1680363874
transform -1 0 4616 0 1 1370
box -8 -3 46 105
use FILL  FILL_8485
timestamp 1680363874
transform 1 0 4616 0 1 1370
box -8 -3 16 105
use FILL  FILL_8493
timestamp 1680363874
transform 1 0 4624 0 1 1370
box -8 -3 16 105
use FILL  FILL_8495
timestamp 1680363874
transform 1 0 4632 0 1 1370
box -8 -3 16 105
use FILL  FILL_8497
timestamp 1680363874
transform 1 0 4640 0 1 1370
box -8 -3 16 105
use FILL  FILL_8499
timestamp 1680363874
transform 1 0 4648 0 1 1370
box -8 -3 16 105
use FILL  FILL_8500
timestamp 1680363874
transform 1 0 4656 0 1 1370
box -8 -3 16 105
use FILL  FILL_8501
timestamp 1680363874
transform 1 0 4664 0 1 1370
box -8 -3 16 105
use FILL  FILL_8502
timestamp 1680363874
transform 1 0 4672 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6424
timestamp 1680363874
transform 1 0 4692 0 1 1375
box -3 -3 3 3
use FILL  FILL_8503
timestamp 1680363874
transform 1 0 4680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8504
timestamp 1680363874
transform 1 0 4688 0 1 1370
box -8 -3 16 105
use FILL  FILL_8506
timestamp 1680363874
transform 1 0 4696 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_436
timestamp 1680363874
transform 1 0 4704 0 1 1370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_67
timestamp 1680363874
transform 1 0 4827 0 1 1370
box -10 -3 10 3
use M3_M2  M3_M2_6425
timestamp 1680363874
transform 1 0 108 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7069
timestamp 1680363874
transform 1 0 100 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7075
timestamp 1680363874
transform 1 0 108 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6560
timestamp 1680363874
transform 1 0 100 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6496
timestamp 1680363874
transform 1 0 132 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6462
timestamp 1680363874
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6463
timestamp 1680363874
transform 1 0 180 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7076
timestamp 1680363874
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6464
timestamp 1680363874
transform 1 0 212 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7077
timestamp 1680363874
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7078
timestamp 1680363874
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7162
timestamp 1680363874
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7163
timestamp 1680363874
transform 1 0 196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7164
timestamp 1680363874
transform 1 0 204 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6523
timestamp 1680363874
transform 1 0 188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6561
timestamp 1680363874
transform 1 0 180 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6465
timestamp 1680363874
transform 1 0 244 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7079
timestamp 1680363874
transform 1 0 244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7165
timestamp 1680363874
transform 1 0 236 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6497
timestamp 1680363874
transform 1 0 260 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7080
timestamp 1680363874
transform 1 0 276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7166
timestamp 1680363874
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7167
timestamp 1680363874
transform 1 0 300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7275
timestamp 1680363874
transform 1 0 268 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6524
timestamp 1680363874
transform 1 0 300 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6426
timestamp 1680363874
transform 1 0 356 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6466
timestamp 1680363874
transform 1 0 388 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7081
timestamp 1680363874
transform 1 0 388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7082
timestamp 1680363874
transform 1 0 396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7168
timestamp 1680363874
transform 1 0 380 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6525
timestamp 1680363874
transform 1 0 396 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6427
timestamp 1680363874
transform 1 0 452 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6441
timestamp 1680363874
transform 1 0 412 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6442
timestamp 1680363874
transform 1 0 436 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6562
timestamp 1680363874
transform 1 0 404 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6467
timestamp 1680363874
transform 1 0 460 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7083
timestamp 1680363874
transform 1 0 460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7169
timestamp 1680363874
transform 1 0 436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7170
timestamp 1680363874
transform 1 0 444 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6526
timestamp 1680363874
transform 1 0 444 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6563
timestamp 1680363874
transform 1 0 436 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6594
timestamp 1680363874
transform 1 0 436 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6595
timestamp 1680363874
transform 1 0 460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6468
timestamp 1680363874
transform 1 0 476 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6469
timestamp 1680363874
transform 1 0 500 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7084
timestamp 1680363874
transform 1 0 500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7085
timestamp 1680363874
transform 1 0 508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7171
timestamp 1680363874
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6527
timestamp 1680363874
transform 1 0 508 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7172
timestamp 1680363874
transform 1 0 540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7173
timestamp 1680363874
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6528
timestamp 1680363874
transform 1 0 548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6564
timestamp 1680363874
transform 1 0 516 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6565
timestamp 1680363874
transform 1 0 540 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6470
timestamp 1680363874
transform 1 0 580 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7086
timestamp 1680363874
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7174
timestamp 1680363874
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7087
timestamp 1680363874
transform 1 0 684 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6508
timestamp 1680363874
transform 1 0 684 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7088
timestamp 1680363874
transform 1 0 724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7175
timestamp 1680363874
transform 1 0 692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7176
timestamp 1680363874
transform 1 0 708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7177
timestamp 1680363874
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7276
timestamp 1680363874
transform 1 0 684 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6566
timestamp 1680363874
transform 1 0 700 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6567
timestamp 1680363874
transform 1 0 716 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6509
timestamp 1680363874
transform 1 0 820 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6471
timestamp 1680363874
transform 1 0 844 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6472
timestamp 1680363874
transform 1 0 860 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7089
timestamp 1680363874
transform 1 0 844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7090
timestamp 1680363874
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7178
timestamp 1680363874
transform 1 0 844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7179
timestamp 1680363874
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7091
timestamp 1680363874
transform 1 0 884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7180
timestamp 1680363874
transform 1 0 924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7092
timestamp 1680363874
transform 1 0 996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7181
timestamp 1680363874
transform 1 0 1012 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6529
timestamp 1680363874
transform 1 0 1012 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6443
timestamp 1680363874
transform 1 0 1036 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7093
timestamp 1680363874
transform 1 0 1036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7094
timestamp 1680363874
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7095
timestamp 1680363874
transform 1 0 1084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7096
timestamp 1680363874
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7182
timestamp 1680363874
transform 1 0 1060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7183
timestamp 1680363874
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6530
timestamp 1680363874
transform 1 0 1076 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6568
timestamp 1680363874
transform 1 0 1060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6569
timestamp 1680363874
transform 1 0 1076 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6596
timestamp 1680363874
transform 1 0 1084 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6498
timestamp 1680363874
transform 1 0 1100 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7184
timestamp 1680363874
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6597
timestamp 1680363874
transform 1 0 1100 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7185
timestamp 1680363874
transform 1 0 1124 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6473
timestamp 1680363874
transform 1 0 1148 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7097
timestamp 1680363874
transform 1 0 1156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7186
timestamp 1680363874
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6444
timestamp 1680363874
transform 1 0 1188 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6474
timestamp 1680363874
transform 1 0 1196 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7098
timestamp 1680363874
transform 1 0 1212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7187
timestamp 1680363874
transform 1 0 1204 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6531
timestamp 1680363874
transform 1 0 1204 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6499
timestamp 1680363874
transform 1 0 1276 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7099
timestamp 1680363874
transform 1 0 1308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7188
timestamp 1680363874
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7189
timestamp 1680363874
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7190
timestamp 1680363874
transform 1 0 1292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7191
timestamp 1680363874
transform 1 0 1308 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6532
timestamp 1680363874
transform 1 0 1308 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7192
timestamp 1680363874
transform 1 0 1356 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6533
timestamp 1680363874
transform 1 0 1348 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6500
timestamp 1680363874
transform 1 0 1372 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6445
timestamp 1680363874
transform 1 0 1468 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7100
timestamp 1680363874
transform 1 0 1468 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6510
timestamp 1680363874
transform 1 0 1396 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7193
timestamp 1680363874
transform 1 0 1420 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6511
timestamp 1680363874
transform 1 0 1468 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6534
timestamp 1680363874
transform 1 0 1420 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6570
timestamp 1680363874
transform 1 0 1404 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6475
timestamp 1680363874
transform 1 0 1484 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7194
timestamp 1680363874
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7101
timestamp 1680363874
transform 1 0 1500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7102
timestamp 1680363874
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7195
timestamp 1680363874
transform 1 0 1556 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6476
timestamp 1680363874
transform 1 0 1588 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7103
timestamp 1680363874
transform 1 0 1588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7196
timestamp 1680363874
transform 1 0 1580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7197
timestamp 1680363874
transform 1 0 1596 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6535
timestamp 1680363874
transform 1 0 1580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6571
timestamp 1680363874
transform 1 0 1596 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7104
timestamp 1680363874
transform 1 0 1716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7198
timestamp 1680363874
transform 1 0 1636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7199
timestamp 1680363874
transform 1 0 1684 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6536
timestamp 1680363874
transform 1 0 1692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6572
timestamp 1680363874
transform 1 0 1724 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7105
timestamp 1680363874
transform 1 0 1764 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6573
timestamp 1680363874
transform 1 0 1764 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7200
timestamp 1680363874
transform 1 0 1780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7106
timestamp 1680363874
transform 1 0 1804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7107
timestamp 1680363874
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7201
timestamp 1680363874
transform 1 0 1812 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6537
timestamp 1680363874
transform 1 0 1812 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7108
timestamp 1680363874
transform 1 0 1844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7202
timestamp 1680363874
transform 1 0 1844 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6538
timestamp 1680363874
transform 1 0 1844 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7280
timestamp 1680363874
transform 1 0 1844 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_7109
timestamp 1680363874
transform 1 0 1876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7203
timestamp 1680363874
transform 1 0 1876 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6446
timestamp 1680363874
transform 1 0 1892 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6447
timestamp 1680363874
transform 1 0 1956 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6477
timestamp 1680363874
transform 1 0 2020 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7110
timestamp 1680363874
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7111
timestamp 1680363874
transform 1 0 2012 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7204
timestamp 1680363874
transform 1 0 1972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7205
timestamp 1680363874
transform 1 0 1980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7206
timestamp 1680363874
transform 1 0 1996 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6574
timestamp 1680363874
transform 1 0 1980 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6448
timestamp 1680363874
transform 1 0 2060 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6501
timestamp 1680363874
transform 1 0 2052 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6478
timestamp 1680363874
transform 1 0 2092 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7112
timestamp 1680363874
transform 1 0 2060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7113
timestamp 1680363874
transform 1 0 2076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7114
timestamp 1680363874
transform 1 0 2092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7115
timestamp 1680363874
transform 1 0 2100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7207
timestamp 1680363874
transform 1 0 2052 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7208
timestamp 1680363874
transform 1 0 2060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7209
timestamp 1680363874
transform 1 0 2084 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6575
timestamp 1680363874
transform 1 0 2052 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6428
timestamp 1680363874
transform 1 0 2108 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6539
timestamp 1680363874
transform 1 0 2100 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7210
timestamp 1680363874
transform 1 0 2116 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6576
timestamp 1680363874
transform 1 0 2116 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6449
timestamp 1680363874
transform 1 0 2140 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7116
timestamp 1680363874
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6502
timestamp 1680363874
transform 1 0 2156 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7117
timestamp 1680363874
transform 1 0 2172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7118
timestamp 1680363874
transform 1 0 2180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7211
timestamp 1680363874
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7212
timestamp 1680363874
transform 1 0 2156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7213
timestamp 1680363874
transform 1 0 2164 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6540
timestamp 1680363874
transform 1 0 2164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6577
timestamp 1680363874
transform 1 0 2140 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6603
timestamp 1680363874
transform 1 0 2164 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7214
timestamp 1680363874
transform 1 0 2228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7277
timestamp 1680363874
transform 1 0 2252 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6503
timestamp 1680363874
transform 1 0 2284 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7215
timestamp 1680363874
transform 1 0 2284 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6512
timestamp 1680363874
transform 1 0 2292 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7119
timestamp 1680363874
transform 1 0 2308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7278
timestamp 1680363874
transform 1 0 2300 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6578
timestamp 1680363874
transform 1 0 2284 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7281
timestamp 1680363874
transform 1 0 2292 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_7070
timestamp 1680363874
transform 1 0 2324 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6504
timestamp 1680363874
transform 1 0 2324 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6604
timestamp 1680363874
transform 1 0 2316 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6429
timestamp 1680363874
transform 1 0 2340 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7120
timestamp 1680363874
transform 1 0 2348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7216
timestamp 1680363874
transform 1 0 2340 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6513
timestamp 1680363874
transform 1 0 2348 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6430
timestamp 1680363874
transform 1 0 2380 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7217
timestamp 1680363874
transform 1 0 2388 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6431
timestamp 1680363874
transform 1 0 2412 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6479
timestamp 1680363874
transform 1 0 2420 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7121
timestamp 1680363874
transform 1 0 2412 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6450
timestamp 1680363874
transform 1 0 2444 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7071
timestamp 1680363874
transform 1 0 2444 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7218
timestamp 1680363874
transform 1 0 2468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7219
timestamp 1680363874
transform 1 0 2476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7279
timestamp 1680363874
transform 1 0 2452 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6514
timestamp 1680363874
transform 1 0 2484 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6579
timestamp 1680363874
transform 1 0 2476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6480
timestamp 1680363874
transform 1 0 2540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7122
timestamp 1680363874
transform 1 0 2500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7123
timestamp 1680363874
transform 1 0 2524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7124
timestamp 1680363874
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7220
timestamp 1680363874
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6515
timestamp 1680363874
transform 1 0 2524 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7221
timestamp 1680363874
transform 1 0 2532 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6605
timestamp 1680363874
transform 1 0 2532 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7222
timestamp 1680363874
transform 1 0 2556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7125
timestamp 1680363874
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6541
timestamp 1680363874
transform 1 0 2604 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7126
timestamp 1680363874
transform 1 0 2628 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6516
timestamp 1680363874
transform 1 0 2628 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7223
timestamp 1680363874
transform 1 0 2636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7127
timestamp 1680363874
transform 1 0 2692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7224
timestamp 1680363874
transform 1 0 2668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7225
timestamp 1680363874
transform 1 0 2684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7226
timestamp 1680363874
transform 1 0 2700 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6542
timestamp 1680363874
transform 1 0 2684 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6598
timestamp 1680363874
transform 1 0 2668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6580
timestamp 1680363874
transform 1 0 2700 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6481
timestamp 1680363874
transform 1 0 2780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7128
timestamp 1680363874
transform 1 0 2732 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6517
timestamp 1680363874
transform 1 0 2732 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7227
timestamp 1680363874
transform 1 0 2780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7228
timestamp 1680363874
transform 1 0 2812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7229
timestamp 1680363874
transform 1 0 2820 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6543
timestamp 1680363874
transform 1 0 2780 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6544
timestamp 1680363874
transform 1 0 2820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6599
timestamp 1680363874
transform 1 0 2820 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7129
timestamp 1680363874
transform 1 0 2844 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6482
timestamp 1680363874
transform 1 0 2900 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7130
timestamp 1680363874
transform 1 0 2892 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6545
timestamp 1680363874
transform 1 0 2892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6600
timestamp 1680363874
transform 1 0 2884 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6483
timestamp 1680363874
transform 1 0 2924 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7131
timestamp 1680363874
transform 1 0 2916 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6432
timestamp 1680363874
transform 1 0 2996 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6451
timestamp 1680363874
transform 1 0 2988 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6484
timestamp 1680363874
transform 1 0 2964 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6485
timestamp 1680363874
transform 1 0 3004 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7132
timestamp 1680363874
transform 1 0 2964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7133
timestamp 1680363874
transform 1 0 2972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7134
timestamp 1680363874
transform 1 0 2988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7135
timestamp 1680363874
transform 1 0 3004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7230
timestamp 1680363874
transform 1 0 2924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7231
timestamp 1680363874
transform 1 0 2932 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6581
timestamp 1680363874
transform 1 0 2924 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6518
timestamp 1680363874
transform 1 0 2940 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7232
timestamp 1680363874
transform 1 0 2948 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7233
timestamp 1680363874
transform 1 0 2972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7234
timestamp 1680363874
transform 1 0 2980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7235
timestamp 1680363874
transform 1 0 2996 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6546
timestamp 1680363874
transform 1 0 2948 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6582
timestamp 1680363874
transform 1 0 2964 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7136
timestamp 1680363874
transform 1 0 3020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7137
timestamp 1680363874
transform 1 0 3052 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6433
timestamp 1680363874
transform 1 0 3100 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6434
timestamp 1680363874
transform 1 0 3124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6435
timestamp 1680363874
transform 1 0 3140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6436
timestamp 1680363874
transform 1 0 3164 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6452
timestamp 1680363874
transform 1 0 3156 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7138
timestamp 1680363874
transform 1 0 3148 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6519
timestamp 1680363874
transform 1 0 3052 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7236
timestamp 1680363874
transform 1 0 3060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7237
timestamp 1680363874
transform 1 0 3068 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6520
timestamp 1680363874
transform 1 0 3076 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7238
timestamp 1680363874
transform 1 0 3100 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6583
timestamp 1680363874
transform 1 0 3060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6584
timestamp 1680363874
transform 1 0 3100 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6585
timestamp 1680363874
transform 1 0 3124 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6601
timestamp 1680363874
transform 1 0 3100 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6606
timestamp 1680363874
transform 1 0 3092 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6453
timestamp 1680363874
transform 1 0 3188 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6602
timestamp 1680363874
transform 1 0 3180 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7139
timestamp 1680363874
transform 1 0 3196 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6505
timestamp 1680363874
transform 1 0 3204 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7140
timestamp 1680363874
transform 1 0 3212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7239
timestamp 1680363874
transform 1 0 3204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7240
timestamp 1680363874
transform 1 0 3220 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6586
timestamp 1680363874
transform 1 0 3204 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7141
timestamp 1680363874
transform 1 0 3252 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6454
timestamp 1680363874
transform 1 0 3260 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7072
timestamp 1680363874
transform 1 0 3260 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6437
timestamp 1680363874
transform 1 0 3308 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6438
timestamp 1680363874
transform 1 0 3340 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6455
timestamp 1680363874
transform 1 0 3284 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6486
timestamp 1680363874
transform 1 0 3364 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7142
timestamp 1680363874
transform 1 0 3364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7241
timestamp 1680363874
transform 1 0 3276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7242
timestamp 1680363874
transform 1 0 3284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7243
timestamp 1680363874
transform 1 0 3324 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6521
timestamp 1680363874
transform 1 0 3332 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6522
timestamp 1680363874
transform 1 0 3364 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6587
timestamp 1680363874
transform 1 0 3276 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6588
timestamp 1680363874
transform 1 0 3324 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6487
timestamp 1680363874
transform 1 0 3396 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7073
timestamp 1680363874
transform 1 0 3404 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6488
timestamp 1680363874
transform 1 0 3444 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7074
timestamp 1680363874
transform 1 0 3452 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7244
timestamp 1680363874
transform 1 0 3436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7143
timestamp 1680363874
transform 1 0 3460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7245
timestamp 1680363874
transform 1 0 3500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6489
timestamp 1680363874
transform 1 0 3532 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7144
timestamp 1680363874
transform 1 0 3532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7246
timestamp 1680363874
transform 1 0 3532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7247
timestamp 1680363874
transform 1 0 3564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7248
timestamp 1680363874
transform 1 0 3580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7249
timestamp 1680363874
transform 1 0 3588 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6547
timestamp 1680363874
transform 1 0 3580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6490
timestamp 1680363874
transform 1 0 3708 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7145
timestamp 1680363874
transform 1 0 3708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7250
timestamp 1680363874
transform 1 0 3676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7251
timestamp 1680363874
transform 1 0 3724 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6607
timestamp 1680363874
transform 1 0 3700 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7146
timestamp 1680363874
transform 1 0 3740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7147
timestamp 1680363874
transform 1 0 3748 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6439
timestamp 1680363874
transform 1 0 3884 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6491
timestamp 1680363874
transform 1 0 3884 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7148
timestamp 1680363874
transform 1 0 3884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7252
timestamp 1680363874
transform 1 0 3796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7253
timestamp 1680363874
transform 1 0 3804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7254
timestamp 1680363874
transform 1 0 3836 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6548
timestamp 1680363874
transform 1 0 3796 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6549
timestamp 1680363874
transform 1 0 3836 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6550
timestamp 1680363874
transform 1 0 3884 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6440
timestamp 1680363874
transform 1 0 3916 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6551
timestamp 1680363874
transform 1 0 3932 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6492
timestamp 1680363874
transform 1 0 3940 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7149
timestamp 1680363874
transform 1 0 3940 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6493
timestamp 1680363874
transform 1 0 3972 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6456
timestamp 1680363874
transform 1 0 4036 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7150
timestamp 1680363874
transform 1 0 4060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7255
timestamp 1680363874
transform 1 0 3972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7256
timestamp 1680363874
transform 1 0 3980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7257
timestamp 1680363874
transform 1 0 4020 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6552
timestamp 1680363874
transform 1 0 3972 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6553
timestamp 1680363874
transform 1 0 4020 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6457
timestamp 1680363874
transform 1 0 4108 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7151
timestamp 1680363874
transform 1 0 4108 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6458
timestamp 1680363874
transform 1 0 4204 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7152
timestamp 1680363874
transform 1 0 4204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7258
timestamp 1680363874
transform 1 0 4132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7259
timestamp 1680363874
transform 1 0 4188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7260
timestamp 1680363874
transform 1 0 4252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7261
timestamp 1680363874
transform 1 0 4284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7262
timestamp 1680363874
transform 1 0 4292 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6554
timestamp 1680363874
transform 1 0 4252 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6555
timestamp 1680363874
transform 1 0 4292 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6589
timestamp 1680363874
transform 1 0 4284 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7153
timestamp 1680363874
transform 1 0 4348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7154
timestamp 1680363874
transform 1 0 4356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7263
timestamp 1680363874
transform 1 0 4340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7264
timestamp 1680363874
transform 1 0 4364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7265
timestamp 1680363874
transform 1 0 4380 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6590
timestamp 1680363874
transform 1 0 4356 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6494
timestamp 1680363874
transform 1 0 4396 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7155
timestamp 1680363874
transform 1 0 4396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7266
timestamp 1680363874
transform 1 0 4396 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6591
timestamp 1680363874
transform 1 0 4388 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6459
timestamp 1680363874
transform 1 0 4428 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7156
timestamp 1680363874
transform 1 0 4428 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6506
timestamp 1680363874
transform 1 0 4516 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6495
timestamp 1680363874
transform 1 0 4540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7157
timestamp 1680363874
transform 1 0 4524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7158
timestamp 1680363874
transform 1 0 4532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7267
timestamp 1680363874
transform 1 0 4468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7268
timestamp 1680363874
transform 1 0 4508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7269
timestamp 1680363874
transform 1 0 4516 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6556
timestamp 1680363874
transform 1 0 4468 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6557
timestamp 1680363874
transform 1 0 4516 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6592
timestamp 1680363874
transform 1 0 4492 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6593
timestamp 1680363874
transform 1 0 4508 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6507
timestamp 1680363874
transform 1 0 4540 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7159
timestamp 1680363874
transform 1 0 4604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7270
timestamp 1680363874
transform 1 0 4612 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6460
timestamp 1680363874
transform 1 0 4660 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7160
timestamp 1680363874
transform 1 0 4676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7271
timestamp 1680363874
transform 1 0 4652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7272
timestamp 1680363874
transform 1 0 4668 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6558
timestamp 1680363874
transform 1 0 4668 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7273
timestamp 1680363874
transform 1 0 4692 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6461
timestamp 1680363874
transform 1 0 4716 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7161
timestamp 1680363874
transform 1 0 4716 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6559
timestamp 1680363874
transform 1 0 4716 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7274
timestamp 1680363874
transform 1 0 4740 0 1 1325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_68
timestamp 1680363874
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_7988
timestamp 1680363874
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8002
timestamp 1680363874
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8003
timestamp 1680363874
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_92
timestamp 1680363874
transform 1 0 96 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8004
timestamp 1680363874
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8005
timestamp 1680363874
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8006
timestamp 1680363874
transform 1 0 136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8007
timestamp 1680363874
transform 1 0 144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8008
timestamp 1680363874
transform 1 0 152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8009
timestamp 1680363874
transform 1 0 160 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_46
timestamp 1680363874
transform 1 0 168 0 -1 1370
box -8 -3 40 105
use NOR2X1  NOR2X1_93
timestamp 1680363874
transform -1 0 224 0 -1 1370
box -8 -3 32 105
use INVX2  INVX2_478
timestamp 1680363874
transform 1 0 224 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8010
timestamp 1680363874
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1680363874
transform 1 0 248 0 -1 1370
box -8 -3 32 105
use XOR2X1  XOR2X1_4
timestamp 1680363874
transform 1 0 272 0 -1 1370
box -8 -3 64 105
use FILL  FILL_8011
timestamp 1680363874
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8013
timestamp 1680363874
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8016
timestamp 1680363874
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8017
timestamp 1680363874
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_47
timestamp 1680363874
transform -1 0 392 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8018
timestamp 1680363874
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8029
timestamp 1680363874
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_5
timestamp 1680363874
transform 1 0 408 0 -1 1370
box -8 -3 64 105
use FILL  FILL_8030
timestamp 1680363874
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_48
timestamp 1680363874
transform -1 0 504 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8031
timestamp 1680363874
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_6
timestamp 1680363874
transform 1 0 512 0 -1 1370
box -8 -3 64 105
use FILL  FILL_8032
timestamp 1680363874
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8034
timestamp 1680363874
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8036
timestamp 1680363874
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8038
timestamp 1680363874
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8041
timestamp 1680363874
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_49
timestamp 1680363874
transform -1 0 640 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8042
timestamp 1680363874
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8044
timestamp 1680363874
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8046
timestamp 1680363874
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8048
timestamp 1680363874
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8050
timestamp 1680363874
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8053
timestamp 1680363874
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_147
timestamp 1680363874
transform -1 0 720 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8054
timestamp 1680363874
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8059
timestamp 1680363874
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8060
timestamp 1680363874
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8061
timestamp 1680363874
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_482
timestamp 1680363874
transform -1 0 768 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8062
timestamp 1680363874
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8064
timestamp 1680363874
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8066
timestamp 1680363874
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8068
timestamp 1680363874
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8069
timestamp 1680363874
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8070
timestamp 1680363874
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8072
timestamp 1680363874
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8074
timestamp 1680363874
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8076
timestamp 1680363874
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_258
timestamp 1680363874
transform 1 0 840 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8080
timestamp 1680363874
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8081
timestamp 1680363874
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8082
timestamp 1680363874
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8084
timestamp 1680363874
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8086
timestamp 1680363874
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8088
timestamp 1680363874
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8090
timestamp 1680363874
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8092
timestamp 1680363874
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8094
timestamp 1680363874
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8096
timestamp 1680363874
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8097
timestamp 1680363874
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8098
timestamp 1680363874
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8100
timestamp 1680363874
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8102
timestamp 1680363874
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_485
timestamp 1680363874
transform 1 0 992 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8106
timestamp 1680363874
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8108
timestamp 1680363874
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8110
timestamp 1680363874
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8112
timestamp 1680363874
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8115
timestamp 1680363874
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_314
timestamp 1680363874
transform 1 0 1048 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8116
timestamp 1680363874
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8118
timestamp 1680363874
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8120
timestamp 1680363874
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8122
timestamp 1680363874
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8124
timestamp 1680363874
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_260
timestamp 1680363874
transform 1 0 1128 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8127
timestamp 1680363874
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8128
timestamp 1680363874
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8130
timestamp 1680363874
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8132
timestamp 1680363874
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8134
timestamp 1680363874
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_487
timestamp 1680363874
transform 1 0 1208 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8142
timestamp 1680363874
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8143
timestamp 1680363874
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8144
timestamp 1680363874
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8145
timestamp 1680363874
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8146
timestamp 1680363874
transform 1 0 1256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8147
timestamp 1680363874
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_261
timestamp 1680363874
transform 1 0 1272 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8148
timestamp 1680363874
transform 1 0 1312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8155
timestamp 1680363874
transform 1 0 1320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8156
timestamp 1680363874
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8157
timestamp 1680363874
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8158
timestamp 1680363874
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_488
timestamp 1680363874
transform -1 0 1368 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8159
timestamp 1680363874
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8160
timestamp 1680363874
transform 1 0 1376 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_417
timestamp 1680363874
transform -1 0 1480 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8161
timestamp 1680363874
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8162
timestamp 1680363874
transform 1 0 1488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8163
timestamp 1680363874
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_489
timestamp 1680363874
transform 1 0 1504 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8164
timestamp 1680363874
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8166
timestamp 1680363874
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8176
timestamp 1680363874
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8177
timestamp 1680363874
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8178
timestamp 1680363874
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_263
timestamp 1680363874
transform 1 0 1560 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8179
timestamp 1680363874
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8180
timestamp 1680363874
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8181
timestamp 1680363874
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8182
timestamp 1680363874
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_419
timestamp 1680363874
transform -1 0 1728 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8183
timestamp 1680363874
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8184
timestamp 1680363874
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8185
timestamp 1680363874
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8186
timestamp 1680363874
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8187
timestamp 1680363874
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8189
timestamp 1680363874
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8191
timestamp 1680363874
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6608
timestamp 1680363874
transform 1 0 1812 0 1 1275
box -3 -3 3 3
use OAI22X1  OAI22X1_317
timestamp 1680363874
transform 1 0 1784 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8198
timestamp 1680363874
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8200
timestamp 1680363874
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8202
timestamp 1680363874
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8204
timestamp 1680363874
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8210
timestamp 1680363874
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_491
timestamp 1680363874
transform -1 0 1880 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8211
timestamp 1680363874
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8212
timestamp 1680363874
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8213
timestamp 1680363874
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8214
timestamp 1680363874
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_492
timestamp 1680363874
transform 1 0 1912 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8215
timestamp 1680363874
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8216
timestamp 1680363874
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8217
timestamp 1680363874
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8218
timestamp 1680363874
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8219
timestamp 1680363874
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8220
timestamp 1680363874
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_264
timestamp 1680363874
transform -1 0 2016 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8221
timestamp 1680363874
transform 1 0 2016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8223
timestamp 1680363874
transform 1 0 2024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8225
timestamp 1680363874
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8231
timestamp 1680363874
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8232
timestamp 1680363874
transform 1 0 2048 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_319
timestamp 1680363874
transform 1 0 2056 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8233
timestamp 1680363874
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8234
timestamp 1680363874
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8235
timestamp 1680363874
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_265
timestamp 1680363874
transform -1 0 2160 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_493
timestamp 1680363874
transform -1 0 2176 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8236
timestamp 1680363874
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8237
timestamp 1680363874
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8238
timestamp 1680363874
transform 1 0 2192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8239
timestamp 1680363874
transform 1 0 2200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8240
timestamp 1680363874
transform 1 0 2208 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_494
timestamp 1680363874
transform 1 0 2216 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8244
timestamp 1680363874
transform 1 0 2232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8247
timestamp 1680363874
transform 1 0 2240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8248
timestamp 1680363874
transform 1 0 2248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8249
timestamp 1680363874
transform 1 0 2256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8250
timestamp 1680363874
transform 1 0 2264 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6609
timestamp 1680363874
transform 1 0 2308 0 1 1275
box -3 -3 3 3
use NAND3X1  NAND3X1_62
timestamp 1680363874
transform 1 0 2272 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8251
timestamp 1680363874
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8252
timestamp 1680363874
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_95
timestamp 1680363874
transform 1 0 2320 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8261
timestamp 1680363874
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8262
timestamp 1680363874
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8263
timestamp 1680363874
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8264
timestamp 1680363874
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8265
timestamp 1680363874
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_96
timestamp 1680363874
transform -1 0 2408 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8266
timestamp 1680363874
transform 1 0 2408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8267
timestamp 1680363874
transform 1 0 2416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8268
timestamp 1680363874
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8269
timestamp 1680363874
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8270
timestamp 1680363874
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_148
timestamp 1680363874
transform -1 0 2480 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8271
timestamp 1680363874
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8272
timestamp 1680363874
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_267
timestamp 1680363874
transform -1 0 2536 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8273
timestamp 1680363874
transform 1 0 2536 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_495
timestamp 1680363874
transform 1 0 2544 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8274
timestamp 1680363874
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8275
timestamp 1680363874
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8276
timestamp 1680363874
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8277
timestamp 1680363874
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8278
timestamp 1680363874
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_496
timestamp 1680363874
transform 1 0 2600 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8281
timestamp 1680363874
transform 1 0 2616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8282
timestamp 1680363874
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8283
timestamp 1680363874
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8284
timestamp 1680363874
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8285
timestamp 1680363874
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8286
timestamp 1680363874
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_268
timestamp 1680363874
transform 1 0 2664 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8287
timestamp 1680363874
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8296
timestamp 1680363874
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6610
timestamp 1680363874
transform 1 0 2804 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_424
timestamp 1680363874
transform 1 0 2720 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8297
timestamp 1680363874
transform 1 0 2816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8298
timestamp 1680363874
transform 1 0 2824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8300
timestamp 1680363874
transform 1 0 2832 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_497
timestamp 1680363874
transform 1 0 2840 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8304
timestamp 1680363874
transform 1 0 2856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8306
timestamp 1680363874
transform 1 0 2864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8308
timestamp 1680363874
transform 1 0 2872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8310
timestamp 1680363874
transform 1 0 2880 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6611
timestamp 1680363874
transform 1 0 2916 0 1 1275
box -3 -3 3 3
use INVX2  INVX2_498
timestamp 1680363874
transform 1 0 2888 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8311
timestamp 1680363874
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8312
timestamp 1680363874
transform 1 0 2912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8313
timestamp 1680363874
transform 1 0 2920 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_270
timestamp 1680363874
transform 1 0 2928 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_320
timestamp 1680363874
transform 1 0 2968 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8325
timestamp 1680363874
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8327
timestamp 1680363874
transform 1 0 3016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8329
timestamp 1680363874
transform 1 0 3024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8330
timestamp 1680363874
transform 1 0 3032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8331
timestamp 1680363874
transform 1 0 3040 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_500
timestamp 1680363874
transform 1 0 3048 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6612
timestamp 1680363874
transform 1 0 3084 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_425
timestamp 1680363874
transform -1 0 3160 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8342
timestamp 1680363874
transform 1 0 3160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8358
timestamp 1680363874
transform 1 0 3168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8359
timestamp 1680363874
transform 1 0 3176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8360
timestamp 1680363874
transform 1 0 3184 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_322
timestamp 1680363874
transform -1 0 3232 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8361
timestamp 1680363874
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8362
timestamp 1680363874
transform 1 0 3240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8363
timestamp 1680363874
transform 1 0 3248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8364
timestamp 1680363874
transform 1 0 3256 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_502
timestamp 1680363874
transform 1 0 3264 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_426
timestamp 1680363874
transform -1 0 3376 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8365
timestamp 1680363874
transform 1 0 3376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8367
timestamp 1680363874
transform 1 0 3384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8369
timestamp 1680363874
transform 1 0 3392 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_98
timestamp 1680363874
transform 1 0 3400 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8374
timestamp 1680363874
transform 1 0 3424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8376
timestamp 1680363874
transform 1 0 3432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8378
timestamp 1680363874
transform 1 0 3440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8379
timestamp 1680363874
transform 1 0 3448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8380
timestamp 1680363874
transform 1 0 3456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8381
timestamp 1680363874
transform 1 0 3464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8382
timestamp 1680363874
transform 1 0 3472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8384
timestamp 1680363874
transform 1 0 3480 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6613
timestamp 1680363874
transform 1 0 3508 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_6614
timestamp 1680363874
transform 1 0 3524 0 1 1275
box -3 -3 3 3
use AND2X2  AND2X2_55
timestamp 1680363874
transform 1 0 3488 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8390
timestamp 1680363874
transform 1 0 3520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8394
timestamp 1680363874
transform 1 0 3528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8395
timestamp 1680363874
transform 1 0 3536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8396
timestamp 1680363874
transform 1 0 3544 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_56
timestamp 1680363874
transform 1 0 3552 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8397
timestamp 1680363874
transform 1 0 3584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8404
timestamp 1680363874
transform 1 0 3592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8405
timestamp 1680363874
transform 1 0 3600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8406
timestamp 1680363874
transform 1 0 3608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8407
timestamp 1680363874
transform 1 0 3616 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_428
timestamp 1680363874
transform -1 0 3720 0 -1 1370
box -8 -3 104 105
use BUFX2  BUFX2_85
timestamp 1680363874
transform 1 0 3720 0 -1 1370
box -5 -3 28 105
use FILL  FILL_8408
timestamp 1680363874
transform 1 0 3744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8409
timestamp 1680363874
transform 1 0 3752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8410
timestamp 1680363874
transform 1 0 3760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8411
timestamp 1680363874
transform 1 0 3768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8413
timestamp 1680363874
transform 1 0 3776 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_504
timestamp 1680363874
transform 1 0 3784 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_430
timestamp 1680363874
transform -1 0 3896 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8418
timestamp 1680363874
transform 1 0 3896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8419
timestamp 1680363874
transform 1 0 3904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8420
timestamp 1680363874
transform 1 0 3912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8421
timestamp 1680363874
transform 1 0 3920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8423
timestamp 1680363874
transform 1 0 3928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8425
timestamp 1680363874
transform 1 0 3936 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_507
timestamp 1680363874
transform 1 0 3944 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8445
timestamp 1680363874
transform 1 0 3960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8446
timestamp 1680363874
transform 1 0 3968 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_432
timestamp 1680363874
transform -1 0 4072 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8447
timestamp 1680363874
transform 1 0 4072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8448
timestamp 1680363874
transform 1 0 4080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8449
timestamp 1680363874
transform 1 0 4088 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_433
timestamp 1680363874
transform 1 0 4096 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_434
timestamp 1680363874
transform 1 0 4192 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8450
timestamp 1680363874
transform 1 0 4288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8451
timestamp 1680363874
transform 1 0 4296 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_508
timestamp 1680363874
transform -1 0 4320 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8452
timestamp 1680363874
transform 1 0 4320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8454
timestamp 1680363874
transform 1 0 4328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8462
timestamp 1680363874
transform 1 0 4336 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_277
timestamp 1680363874
transform -1 0 4384 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8463
timestamp 1680363874
transform 1 0 4384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8465
timestamp 1680363874
transform 1 0 4392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8467
timestamp 1680363874
transform 1 0 4400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8469
timestamp 1680363874
transform 1 0 4408 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_435
timestamp 1680363874
transform 1 0 4416 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_509
timestamp 1680363874
transform -1 0 4528 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8480
timestamp 1680363874
transform 1 0 4528 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_510
timestamp 1680363874
transform 1 0 4536 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8481
timestamp 1680363874
transform 1 0 4552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8483
timestamp 1680363874
transform 1 0 4560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8486
timestamp 1680363874
transform 1 0 4568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8487
timestamp 1680363874
transform 1 0 4576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8488
timestamp 1680363874
transform 1 0 4584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8489
timestamp 1680363874
transform 1 0 4592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8490
timestamp 1680363874
transform 1 0 4600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8491
timestamp 1680363874
transform 1 0 4608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8492
timestamp 1680363874
transform 1 0 4616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8494
timestamp 1680363874
transform 1 0 4624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8496
timestamp 1680363874
transform 1 0 4632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8498
timestamp 1680363874
transform 1 0 4640 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_280
timestamp 1680363874
transform 1 0 4648 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8505
timestamp 1680363874
transform 1 0 4688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8507
timestamp 1680363874
transform 1 0 4696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8508
timestamp 1680363874
transform 1 0 4704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8509
timestamp 1680363874
transform 1 0 4712 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_511
timestamp 1680363874
transform 1 0 4720 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8510
timestamp 1680363874
transform 1 0 4736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8511
timestamp 1680363874
transform 1 0 4744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8512
timestamp 1680363874
transform 1 0 4752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8513
timestamp 1680363874
transform 1 0 4760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8514
timestamp 1680363874
transform 1 0 4768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8515
timestamp 1680363874
transform 1 0 4776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8516
timestamp 1680363874
transform 1 0 4784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8517
timestamp 1680363874
transform 1 0 4792 0 -1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_69
timestamp 1680363874
transform 1 0 4851 0 1 1270
box -10 -3 10 3
use M2_M1  M2_M1_7401
timestamp 1680363874
transform 1 0 76 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6790
timestamp 1680363874
transform 1 0 84 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7295
timestamp 1680363874
transform 1 0 100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7402
timestamp 1680363874
transform 1 0 100 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6755
timestamp 1680363874
transform 1 0 92 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7403
timestamp 1680363874
transform 1 0 116 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7296
timestamp 1680363874
transform 1 0 156 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6617
timestamp 1680363874
transform 1 0 188 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6632
timestamp 1680363874
transform 1 0 180 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7404
timestamp 1680363874
transform 1 0 172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6618
timestamp 1680363874
transform 1 0 212 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6633
timestamp 1680363874
transform 1 0 220 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6674
timestamp 1680363874
transform 1 0 292 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7297
timestamp 1680363874
transform 1 0 252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7298
timestamp 1680363874
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7405
timestamp 1680363874
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6756
timestamp 1680363874
transform 1 0 204 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6757
timestamp 1680363874
transform 1 0 276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6791
timestamp 1680363874
transform 1 0 196 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7406
timestamp 1680363874
transform 1 0 292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7283
timestamp 1680363874
transform 1 0 324 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6650
timestamp 1680363874
transform 1 0 340 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7299
timestamp 1680363874
transform 1 0 340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7407
timestamp 1680363874
transform 1 0 332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6738
timestamp 1680363874
transform 1 0 340 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6651
timestamp 1680363874
transform 1 0 372 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7284
timestamp 1680363874
transform 1 0 372 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6675
timestamp 1680363874
transform 1 0 380 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7300
timestamp 1680363874
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6739
timestamp 1680363874
transform 1 0 356 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7301
timestamp 1680363874
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7302
timestamp 1680363874
transform 1 0 412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7408
timestamp 1680363874
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7409
timestamp 1680363874
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6758
timestamp 1680363874
transform 1 0 372 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6759
timestamp 1680363874
transform 1 0 412 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6760
timestamp 1680363874
transform 1 0 460 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7303
timestamp 1680363874
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6740
timestamp 1680363874
transform 1 0 476 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7410
timestamp 1680363874
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6761
timestamp 1680363874
transform 1 0 492 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7411
timestamp 1680363874
transform 1 0 516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7285
timestamp 1680363874
transform 1 0 540 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7286
timestamp 1680363874
transform 1 0 548 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7287
timestamp 1680363874
transform 1 0 564 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7288
timestamp 1680363874
transform 1 0 588 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7412
timestamp 1680363874
transform 1 0 580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7289
timestamp 1680363874
transform 1 0 604 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7304
timestamp 1680363874
transform 1 0 596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7413
timestamp 1680363874
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6741
timestamp 1680363874
transform 1 0 620 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7414
timestamp 1680363874
transform 1 0 660 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6652
timestamp 1680363874
transform 1 0 692 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7290
timestamp 1680363874
transform 1 0 692 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7305
timestamp 1680363874
transform 1 0 684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7415
timestamp 1680363874
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6634
timestamp 1680363874
transform 1 0 788 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6653
timestamp 1680363874
transform 1 0 764 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6676
timestamp 1680363874
transform 1 0 820 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7306
timestamp 1680363874
transform 1 0 764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7307
timestamp 1680363874
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7416
timestamp 1680363874
transform 1 0 740 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6792
timestamp 1680363874
transform 1 0 740 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7417
timestamp 1680363874
transform 1 0 828 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6677
timestamp 1680363874
transform 1 0 892 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7308
timestamp 1680363874
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7309
timestamp 1680363874
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6635
timestamp 1680363874
transform 1 0 940 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6654
timestamp 1680363874
transform 1 0 972 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7310
timestamp 1680363874
transform 1 0 972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7311
timestamp 1680363874
transform 1 0 1004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7418
timestamp 1680363874
transform 1 0 924 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6762
timestamp 1680363874
transform 1 0 924 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7419
timestamp 1680363874
transform 1 0 1012 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6619
timestamp 1680363874
transform 1 0 1060 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6636
timestamp 1680363874
transform 1 0 1076 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6655
timestamp 1680363874
transform 1 0 1068 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6678
timestamp 1680363874
transform 1 0 1068 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6679
timestamp 1680363874
transform 1 0 1092 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7312
timestamp 1680363874
transform 1 0 1068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7313
timestamp 1680363874
transform 1 0 1076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7314
timestamp 1680363874
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7420
timestamp 1680363874
transform 1 0 1060 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6715
timestamp 1680363874
transform 1 0 1100 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7421
timestamp 1680363874
transform 1 0 1084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7422
timestamp 1680363874
transform 1 0 1100 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6620
timestamp 1680363874
transform 1 0 1172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6680
timestamp 1680363874
transform 1 0 1204 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6637
timestamp 1680363874
transform 1 0 1228 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7315
timestamp 1680363874
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7316
timestamp 1680363874
transform 1 0 1220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7317
timestamp 1680363874
transform 1 0 1228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7423
timestamp 1680363874
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6763
timestamp 1680363874
transform 1 0 1140 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6764
timestamp 1680363874
transform 1 0 1188 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6638
timestamp 1680363874
transform 1 0 1292 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7318
timestamp 1680363874
transform 1 0 1276 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6716
timestamp 1680363874
transform 1 0 1284 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7319
timestamp 1680363874
transform 1 0 1292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7424
timestamp 1680363874
transform 1 0 1252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7425
timestamp 1680363874
transform 1 0 1268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7426
timestamp 1680363874
transform 1 0 1284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7427
timestamp 1680363874
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6765
timestamp 1680363874
transform 1 0 1268 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6615
timestamp 1680363874
transform 1 0 1308 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6656
timestamp 1680363874
transform 1 0 1300 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7428
timestamp 1680363874
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6657
timestamp 1680363874
transform 1 0 1340 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6681
timestamp 1680363874
transform 1 0 1332 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7320
timestamp 1680363874
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7321
timestamp 1680363874
transform 1 0 1356 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6717
timestamp 1680363874
transform 1 0 1364 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7429
timestamp 1680363874
transform 1 0 1348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7430
timestamp 1680363874
transform 1 0 1364 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6793
timestamp 1680363874
transform 1 0 1340 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7322
timestamp 1680363874
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7431
timestamp 1680363874
transform 1 0 1396 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6766
timestamp 1680363874
transform 1 0 1444 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6794
timestamp 1680363874
transform 1 0 1444 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6767
timestamp 1680363874
transform 1 0 1524 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6718
timestamp 1680363874
transform 1 0 1540 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7432
timestamp 1680363874
transform 1 0 1532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7323
timestamp 1680363874
transform 1 0 1620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7433
timestamp 1680363874
transform 1 0 1636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6658
timestamp 1680363874
transform 1 0 1700 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6621
timestamp 1680363874
transform 1 0 1764 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6682
timestamp 1680363874
transform 1 0 1748 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7324
timestamp 1680363874
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7325
timestamp 1680363874
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7326
timestamp 1680363874
transform 1 0 1764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7434
timestamp 1680363874
transform 1 0 1732 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7435
timestamp 1680363874
transform 1 0 1740 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6795
timestamp 1680363874
transform 1 0 1748 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7436
timestamp 1680363874
transform 1 0 1772 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7282
timestamp 1680363874
transform 1 0 1812 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_7291
timestamp 1680363874
transform 1 0 1796 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6683
timestamp 1680363874
transform 1 0 1804 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7327
timestamp 1680363874
transform 1 0 1804 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6719
timestamp 1680363874
transform 1 0 1820 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7292
timestamp 1680363874
transform 1 0 1868 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6796
timestamp 1680363874
transform 1 0 1860 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6622
timestamp 1680363874
transform 1 0 1932 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7328
timestamp 1680363874
transform 1 0 1876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7329
timestamp 1680363874
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7437
timestamp 1680363874
transform 1 0 1956 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6768
timestamp 1680363874
transform 1 0 1932 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6623
timestamp 1680363874
transform 1 0 1980 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6684
timestamp 1680363874
transform 1 0 1972 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7438
timestamp 1680363874
transform 1 0 1972 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6685
timestamp 1680363874
transform 1 0 2004 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6720
timestamp 1680363874
transform 1 0 1996 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7330
timestamp 1680363874
transform 1 0 2004 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6721
timestamp 1680363874
transform 1 0 2012 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6659
timestamp 1680363874
transform 1 0 2036 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7439
timestamp 1680363874
transform 1 0 2012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7440
timestamp 1680363874
transform 1 0 2028 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7441
timestamp 1680363874
transform 1 0 2036 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6769
timestamp 1680363874
transform 1 0 2012 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7331
timestamp 1680363874
transform 1 0 2060 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6686
timestamp 1680363874
transform 1 0 2076 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6687
timestamp 1680363874
transform 1 0 2100 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7332
timestamp 1680363874
transform 1 0 2100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7442
timestamp 1680363874
transform 1 0 2076 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7333
timestamp 1680363874
transform 1 0 2172 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6660
timestamp 1680363874
transform 1 0 2268 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6688
timestamp 1680363874
transform 1 0 2236 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6689
timestamp 1680363874
transform 1 0 2276 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7334
timestamp 1680363874
transform 1 0 2236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7335
timestamp 1680363874
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7336
timestamp 1680363874
transform 1 0 2276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7443
timestamp 1680363874
transform 1 0 2188 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6639
timestamp 1680363874
transform 1 0 2300 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6661
timestamp 1680363874
transform 1 0 2316 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6690
timestamp 1680363874
transform 1 0 2324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6624
timestamp 1680363874
transform 1 0 2372 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6625
timestamp 1680363874
transform 1 0 2404 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6626
timestamp 1680363874
transform 1 0 2428 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6640
timestamp 1680363874
transform 1 0 2364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6662
timestamp 1680363874
transform 1 0 2364 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7293
timestamp 1680363874
transform 1 0 2340 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7337
timestamp 1680363874
transform 1 0 2324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7444
timestamp 1680363874
transform 1 0 2308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7445
timestamp 1680363874
transform 1 0 2316 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6797
timestamp 1680363874
transform 1 0 2308 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6641
timestamp 1680363874
transform 1 0 2396 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6663
timestamp 1680363874
transform 1 0 2428 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6664
timestamp 1680363874
transform 1 0 2444 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7294
timestamp 1680363874
transform 1 0 2412 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6691
timestamp 1680363874
transform 1 0 2428 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7338
timestamp 1680363874
transform 1 0 2348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7339
timestamp 1680363874
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7340
timestamp 1680363874
transform 1 0 2380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7446
timestamp 1680363874
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6722
timestamp 1680363874
transform 1 0 2388 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7341
timestamp 1680363874
transform 1 0 2396 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6723
timestamp 1680363874
transform 1 0 2412 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7342
timestamp 1680363874
transform 1 0 2428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7447
timestamp 1680363874
transform 1 0 2372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7448
timestamp 1680363874
transform 1 0 2404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7449
timestamp 1680363874
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7343
timestamp 1680363874
transform 1 0 2444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7450
timestamp 1680363874
transform 1 0 2436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7451
timestamp 1680363874
transform 1 0 2444 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6770
timestamp 1680363874
transform 1 0 2436 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6665
timestamp 1680363874
transform 1 0 2476 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6692
timestamp 1680363874
transform 1 0 2468 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7344
timestamp 1680363874
transform 1 0 2468 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6642
timestamp 1680363874
transform 1 0 2492 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7345
timestamp 1680363874
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7452
timestamp 1680363874
transform 1 0 2476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7453
timestamp 1680363874
transform 1 0 2484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6771
timestamp 1680363874
transform 1 0 2492 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6798
timestamp 1680363874
transform 1 0 2468 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6799
timestamp 1680363874
transform 1 0 2484 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7346
timestamp 1680363874
transform 1 0 2556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7454
timestamp 1680363874
transform 1 0 2580 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6772
timestamp 1680363874
transform 1 0 2516 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7347
timestamp 1680363874
transform 1 0 2668 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6616
timestamp 1680363874
transform 1 0 2708 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6643
timestamp 1680363874
transform 1 0 2700 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6666
timestamp 1680363874
transform 1 0 2684 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7348
timestamp 1680363874
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6627
timestamp 1680363874
transform 1 0 2764 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7349
timestamp 1680363874
transform 1 0 2764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7455
timestamp 1680363874
transform 1 0 2756 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6773
timestamp 1680363874
transform 1 0 2772 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6724
timestamp 1680363874
transform 1 0 2796 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7350
timestamp 1680363874
transform 1 0 2804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7351
timestamp 1680363874
transform 1 0 2820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7352
timestamp 1680363874
transform 1 0 2836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7456
timestamp 1680363874
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7457
timestamp 1680363874
transform 1 0 2844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6774
timestamp 1680363874
transform 1 0 2812 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6775
timestamp 1680363874
transform 1 0 2844 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6693
timestamp 1680363874
transform 1 0 2860 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7353
timestamp 1680363874
transform 1 0 2860 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6667
timestamp 1680363874
transform 1 0 2932 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6694
timestamp 1680363874
transform 1 0 2972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6695
timestamp 1680363874
transform 1 0 3028 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7354
timestamp 1680363874
transform 1 0 2964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7355
timestamp 1680363874
transform 1 0 3020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7356
timestamp 1680363874
transform 1 0 3028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7458
timestamp 1680363874
transform 1 0 2940 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6742
timestamp 1680363874
transform 1 0 3004 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6725
timestamp 1680363874
transform 1 0 3052 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6696
timestamp 1680363874
transform 1 0 3092 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7357
timestamp 1680363874
transform 1 0 3076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7358
timestamp 1680363874
transform 1 0 3092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7459
timestamp 1680363874
transform 1 0 3068 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7460
timestamp 1680363874
transform 1 0 3084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7461
timestamp 1680363874
transform 1 0 3236 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6800
timestamp 1680363874
transform 1 0 3244 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6644
timestamp 1680363874
transform 1 0 3260 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6743
timestamp 1680363874
transform 1 0 3268 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7359
timestamp 1680363874
transform 1 0 3348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6668
timestamp 1680363874
transform 1 0 3412 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7360
timestamp 1680363874
transform 1 0 3444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7462
timestamp 1680363874
transform 1 0 3476 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6628
timestamp 1680363874
transform 1 0 3500 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7361
timestamp 1680363874
transform 1 0 3508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7463
timestamp 1680363874
transform 1 0 3500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7464
timestamp 1680363874
transform 1 0 3532 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6629
timestamp 1680363874
transform 1 0 3564 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6669
timestamp 1680363874
transform 1 0 3556 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7362
timestamp 1680363874
transform 1 0 3548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7363
timestamp 1680363874
transform 1 0 3556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7364
timestamp 1680363874
transform 1 0 3572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7465
timestamp 1680363874
transform 1 0 3564 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6744
timestamp 1680363874
transform 1 0 3572 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7466
timestamp 1680363874
transform 1 0 3580 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6745
timestamp 1680363874
transform 1 0 3588 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7467
timestamp 1680363874
transform 1 0 3596 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6776
timestamp 1680363874
transform 1 0 3564 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7365
timestamp 1680363874
transform 1 0 3604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7366
timestamp 1680363874
transform 1 0 3652 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6726
timestamp 1680363874
transform 1 0 3660 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6777
timestamp 1680363874
transform 1 0 3652 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7468
timestamp 1680363874
transform 1 0 3668 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6778
timestamp 1680363874
transform 1 0 3668 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6697
timestamp 1680363874
transform 1 0 3684 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7367
timestamp 1680363874
transform 1 0 3676 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7368
timestamp 1680363874
transform 1 0 3684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7369
timestamp 1680363874
transform 1 0 3708 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6698
timestamp 1680363874
transform 1 0 3724 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7370
timestamp 1680363874
transform 1 0 3740 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6727
timestamp 1680363874
transform 1 0 3748 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7371
timestamp 1680363874
transform 1 0 3756 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6699
timestamp 1680363874
transform 1 0 3780 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7372
timestamp 1680363874
transform 1 0 3804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7469
timestamp 1680363874
transform 1 0 3796 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6746
timestamp 1680363874
transform 1 0 3804 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7470
timestamp 1680363874
transform 1 0 3812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7471
timestamp 1680363874
transform 1 0 3828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7472
timestamp 1680363874
transform 1 0 3836 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6779
timestamp 1680363874
transform 1 0 3836 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6645
timestamp 1680363874
transform 1 0 3852 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6646
timestamp 1680363874
transform 1 0 3876 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7373
timestamp 1680363874
transform 1 0 3860 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6728
timestamp 1680363874
transform 1 0 3868 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6700
timestamp 1680363874
transform 1 0 3908 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7374
timestamp 1680363874
transform 1 0 3876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7375
timestamp 1680363874
transform 1 0 3892 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6801
timestamp 1680363874
transform 1 0 3860 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6729
timestamp 1680363874
transform 1 0 3900 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7376
timestamp 1680363874
transform 1 0 3908 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6747
timestamp 1680363874
transform 1 0 3876 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7473
timestamp 1680363874
transform 1 0 3900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7474
timestamp 1680363874
transform 1 0 3908 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6802
timestamp 1680363874
transform 1 0 3892 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6647
timestamp 1680363874
transform 1 0 3948 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6701
timestamp 1680363874
transform 1 0 3956 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6702
timestamp 1680363874
transform 1 0 3996 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7377
timestamp 1680363874
transform 1 0 3956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7378
timestamp 1680363874
transform 1 0 3964 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6730
timestamp 1680363874
transform 1 0 3972 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7379
timestamp 1680363874
transform 1 0 3996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7475
timestamp 1680363874
transform 1 0 4044 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6731
timestamp 1680363874
transform 1 0 4068 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6748
timestamp 1680363874
transform 1 0 4076 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6703
timestamp 1680363874
transform 1 0 4092 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7476
timestamp 1680363874
transform 1 0 4092 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7477
timestamp 1680363874
transform 1 0 4108 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6780
timestamp 1680363874
transform 1 0 4108 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6670
timestamp 1680363874
transform 1 0 4172 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6704
timestamp 1680363874
transform 1 0 4156 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7380
timestamp 1680363874
transform 1 0 4132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7381
timestamp 1680363874
transform 1 0 4140 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6732
timestamp 1680363874
transform 1 0 4148 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7382
timestamp 1680363874
transform 1 0 4156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7383
timestamp 1680363874
transform 1 0 4172 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6749
timestamp 1680363874
transform 1 0 4140 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7478
timestamp 1680363874
transform 1 0 4148 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6781
timestamp 1680363874
transform 1 0 4148 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7479
timestamp 1680363874
transform 1 0 4180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7384
timestamp 1680363874
transform 1 0 4188 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6733
timestamp 1680363874
transform 1 0 4196 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6782
timestamp 1680363874
transform 1 0 4188 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7385
timestamp 1680363874
transform 1 0 4228 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6734
timestamp 1680363874
transform 1 0 4236 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7480
timestamp 1680363874
transform 1 0 4204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7481
timestamp 1680363874
transform 1 0 4220 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6750
timestamp 1680363874
transform 1 0 4228 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7482
timestamp 1680363874
transform 1 0 4236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7483
timestamp 1680363874
transform 1 0 4244 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6783
timestamp 1680363874
transform 1 0 4236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6705
timestamp 1680363874
transform 1 0 4260 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6706
timestamp 1680363874
transform 1 0 4300 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7386
timestamp 1680363874
transform 1 0 4260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7387
timestamp 1680363874
transform 1 0 4268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7388
timestamp 1680363874
transform 1 0 4300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7484
timestamp 1680363874
transform 1 0 4348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6784
timestamp 1680363874
transform 1 0 4268 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6803
timestamp 1680363874
transform 1 0 4348 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6648
timestamp 1680363874
transform 1 0 4436 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6649
timestamp 1680363874
transform 1 0 4476 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6671
timestamp 1680363874
transform 1 0 4452 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6707
timestamp 1680363874
transform 1 0 4420 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6708
timestamp 1680363874
transform 1 0 4460 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7389
timestamp 1680363874
transform 1 0 4420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7390
timestamp 1680363874
transform 1 0 4452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7391
timestamp 1680363874
transform 1 0 4460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7485
timestamp 1680363874
transform 1 0 4372 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6785
timestamp 1680363874
transform 1 0 4444 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7392
timestamp 1680363874
transform 1 0 4476 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6672
timestamp 1680363874
transform 1 0 4492 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6709
timestamp 1680363874
transform 1 0 4500 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7393
timestamp 1680363874
transform 1 0 4500 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6673
timestamp 1680363874
transform 1 0 4524 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6735
timestamp 1680363874
transform 1 0 4532 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7486
timestamp 1680363874
transform 1 0 4484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7487
timestamp 1680363874
transform 1 0 4492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7488
timestamp 1680363874
transform 1 0 4508 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7489
timestamp 1680363874
transform 1 0 4516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7490
timestamp 1680363874
transform 1 0 4524 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6710
timestamp 1680363874
transform 1 0 4564 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6630
timestamp 1680363874
transform 1 0 4652 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6711
timestamp 1680363874
transform 1 0 4596 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6712
timestamp 1680363874
transform 1 0 4628 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7394
timestamp 1680363874
transform 1 0 4548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7395
timestamp 1680363874
transform 1 0 4564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7396
timestamp 1680363874
transform 1 0 4580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7397
timestamp 1680363874
transform 1 0 4612 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6736
timestamp 1680363874
transform 1 0 4628 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7491
timestamp 1680363874
transform 1 0 4556 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6751
timestamp 1680363874
transform 1 0 4564 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7492
timestamp 1680363874
transform 1 0 4572 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6752
timestamp 1680363874
transform 1 0 4580 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7493
timestamp 1680363874
transform 1 0 4660 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6786
timestamp 1680363874
transform 1 0 4556 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6787
timestamp 1680363874
transform 1 0 4572 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6737
timestamp 1680363874
transform 1 0 4676 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7494
timestamp 1680363874
transform 1 0 4676 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6788
timestamp 1680363874
transform 1 0 4676 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6631
timestamp 1680363874
transform 1 0 4716 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6713
timestamp 1680363874
transform 1 0 4692 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6714
timestamp 1680363874
transform 1 0 4740 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7398
timestamp 1680363874
transform 1 0 4692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7399
timestamp 1680363874
transform 1 0 4700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7400
timestamp 1680363874
transform 1 0 4732 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6753
timestamp 1680363874
transform 1 0 4692 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6754
timestamp 1680363874
transform 1 0 4732 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7495
timestamp 1680363874
transform 1 0 4780 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6789
timestamp 1680363874
transform 1 0 4700 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6804
timestamp 1680363874
transform 1 0 4780 0 1 1185
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_70
timestamp 1680363874
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_8518
timestamp 1680363874
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_8520
timestamp 1680363874
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_8521
timestamp 1680363874
transform 1 0 88 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_512
timestamp 1680363874
transform 1 0 96 0 1 1170
box -9 -3 26 105
use FILL  FILL_8522
timestamp 1680363874
transform 1 0 112 0 1 1170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_1
timestamp 1680363874
transform 1 0 120 0 1 1170
box -8 -3 64 105
use FILL  FILL_8523
timestamp 1680363874
transform 1 0 176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8525
timestamp 1680363874
transform 1 0 184 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_438
timestamp 1680363874
transform 1 0 192 0 1 1170
box -8 -3 104 105
use FILL  FILL_8526
timestamp 1680363874
transform 1 0 288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8529
timestamp 1680363874
transform 1 0 296 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_49
timestamp 1680363874
transform 1 0 304 0 1 1170
box -8 -3 32 105
use FILL  FILL_8531
timestamp 1680363874
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8532
timestamp 1680363874
transform 1 0 336 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_149
timestamp 1680363874
transform 1 0 344 0 1 1170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_440
timestamp 1680363874
transform -1 0 472 0 1 1170
box -8 -3 104 105
use FILL  FILL_8533
timestamp 1680363874
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_8545
timestamp 1680363874
transform 1 0 480 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_151
timestamp 1680363874
transform 1 0 488 0 1 1170
box -8 -3 34 105
use FILL  FILL_8546
timestamp 1680363874
transform 1 0 520 0 1 1170
box -8 -3 16 105
use FILL  FILL_8547
timestamp 1680363874
transform 1 0 528 0 1 1170
box -8 -3 16 105
use FILL  FILL_8548
timestamp 1680363874
transform 1 0 536 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1680363874
transform -1 0 568 0 1 1170
box -8 -3 32 105
use FILL  FILL_8549
timestamp 1680363874
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_8550
timestamp 1680363874
transform 1 0 576 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_51
timestamp 1680363874
transform -1 0 608 0 1 1170
box -8 -3 32 105
use FILL  FILL_8551
timestamp 1680363874
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_8552
timestamp 1680363874
transform 1 0 616 0 1 1170
box -8 -3 16 105
use FILL  FILL_8553
timestamp 1680363874
transform 1 0 624 0 1 1170
box -8 -3 16 105
use FILL  FILL_8554
timestamp 1680363874
transform 1 0 632 0 1 1170
box -8 -3 16 105
use FILL  FILL_8559
timestamp 1680363874
transform 1 0 640 0 1 1170
box -8 -3 16 105
use FILL  FILL_8561
timestamp 1680363874
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8563
timestamp 1680363874
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8565
timestamp 1680363874
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8566
timestamp 1680363874
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8567
timestamp 1680363874
transform 1 0 680 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_52
timestamp 1680363874
transform -1 0 712 0 1 1170
box -8 -3 32 105
use FILL  FILL_8568
timestamp 1680363874
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_8569
timestamp 1680363874
transform 1 0 720 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_442
timestamp 1680363874
transform 1 0 728 0 1 1170
box -8 -3 104 105
use FILL  FILL_8571
timestamp 1680363874
transform 1 0 824 0 1 1170
box -8 -3 16 105
use FILL  FILL_8572
timestamp 1680363874
transform 1 0 832 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6805
timestamp 1680363874
transform 1 0 876 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_7
timestamp 1680363874
transform 1 0 840 0 1 1170
box -8 -3 64 105
use FILL  FILL_8573
timestamp 1680363874
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_8584
timestamp 1680363874
transform 1 0 904 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_444
timestamp 1680363874
transform 1 0 912 0 1 1170
box -8 -3 104 105
use FILL  FILL_8586
timestamp 1680363874
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6806
timestamp 1680363874
transform 1 0 1044 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_513
timestamp 1680363874
transform 1 0 1016 0 1 1170
box -9 -3 26 105
use FILL  FILL_8587
timestamp 1680363874
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_8588
timestamp 1680363874
transform 1 0 1040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8589
timestamp 1680363874
transform 1 0 1048 0 1 1170
box -8 -3 16 105
use FILL  FILL_8590
timestamp 1680363874
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_323
timestamp 1680363874
transform 1 0 1064 0 1 1170
box -8 -3 46 105
use FILL  FILL_8591
timestamp 1680363874
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8592
timestamp 1680363874
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8593
timestamp 1680363874
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6807
timestamp 1680363874
transform 1 0 1140 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_447
timestamp 1680363874
transform 1 0 1128 0 1 1170
box -8 -3 104 105
use FILL  FILL_8595
timestamp 1680363874
transform 1 0 1224 0 1 1170
box -8 -3 16 105
use FILL  FILL_8596
timestamp 1680363874
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use FILL  FILL_8597
timestamp 1680363874
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_324
timestamp 1680363874
transform 1 0 1248 0 1 1170
box -8 -3 46 105
use FILL  FILL_8598
timestamp 1680363874
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8599
timestamp 1680363874
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8600
timestamp 1680363874
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_8601
timestamp 1680363874
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use FILL  FILL_8602
timestamp 1680363874
transform 1 0 1320 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_326
timestamp 1680363874
transform 1 0 1328 0 1 1170
box -8 -3 46 105
use FILL  FILL_8614
timestamp 1680363874
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_8615
timestamp 1680363874
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6808
timestamp 1680363874
transform 1 0 1396 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_448
timestamp 1680363874
transform 1 0 1384 0 1 1170
box -8 -3 104 105
use FILL  FILL_8616
timestamp 1680363874
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_8625
timestamp 1680363874
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_8627
timestamp 1680363874
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_515
timestamp 1680363874
transform 1 0 1504 0 1 1170
box -9 -3 26 105
use FILL  FILL_8629
timestamp 1680363874
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_8630
timestamp 1680363874
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6809
timestamp 1680363874
transform 1 0 1548 0 1 1175
box -3 -3 3 3
use FILL  FILL_8631
timestamp 1680363874
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_8632
timestamp 1680363874
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_8634
timestamp 1680363874
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_8636
timestamp 1680363874
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_8638
timestamp 1680363874
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use FILL  FILL_8640
timestamp 1680363874
transform 1 0 1576 0 1 1170
box -8 -3 16 105
use FILL  FILL_8642
timestamp 1680363874
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use FILL  FILL_8643
timestamp 1680363874
transform 1 0 1592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8644
timestamp 1680363874
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use FILL  FILL_8645
timestamp 1680363874
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_8646
timestamp 1680363874
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_8647
timestamp 1680363874
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_8649
timestamp 1680363874
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_8651
timestamp 1680363874
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6810
timestamp 1680363874
transform 1 0 1668 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_516
timestamp 1680363874
transform 1 0 1648 0 1 1170
box -9 -3 26 105
use FILL  FILL_8653
timestamp 1680363874
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8654
timestamp 1680363874
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8655
timestamp 1680363874
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_8656
timestamp 1680363874
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_8657
timestamp 1680363874
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_8658
timestamp 1680363874
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_8662
timestamp 1680363874
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_8664
timestamp 1680363874
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_283
timestamp 1680363874
transform 1 0 1728 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_6811
timestamp 1680363874
transform 1 0 1780 0 1 1175
box -3 -3 3 3
use FILL  FILL_8666
timestamp 1680363874
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8667
timestamp 1680363874
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8668
timestamp 1680363874
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1680363874
transform 1 0 1792 0 1 1170
box -8 -3 40 105
use FILL  FILL_8672
timestamp 1680363874
transform 1 0 1824 0 1 1170
box -8 -3 16 105
use FILL  FILL_8676
timestamp 1680363874
transform 1 0 1832 0 1 1170
box -8 -3 16 105
use FILL  FILL_8678
timestamp 1680363874
transform 1 0 1840 0 1 1170
box -8 -3 16 105
use FILL  FILL_8680
timestamp 1680363874
transform 1 0 1848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8682
timestamp 1680363874
transform 1 0 1856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8683
timestamp 1680363874
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6812
timestamp 1680363874
transform 1 0 1972 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_450
timestamp 1680363874
transform -1 0 1968 0 1 1170
box -8 -3 104 105
use FILL  FILL_8684
timestamp 1680363874
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_8688
timestamp 1680363874
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_8689
timestamp 1680363874
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6813
timestamp 1680363874
transform 1 0 2004 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6814
timestamp 1680363874
transform 1 0 2020 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_330
timestamp 1680363874
transform -1 0 2032 0 1 1170
box -8 -3 46 105
use FILL  FILL_8690
timestamp 1680363874
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_8697
timestamp 1680363874
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8699
timestamp 1680363874
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_8701
timestamp 1680363874
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_452
timestamp 1680363874
transform 1 0 2064 0 1 1170
box -8 -3 104 105
use FILL  FILL_8703
timestamp 1680363874
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8712
timestamp 1680363874
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6815
timestamp 1680363874
transform 1 0 2196 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6816
timestamp 1680363874
transform 1 0 2220 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_453
timestamp 1680363874
transform 1 0 2176 0 1 1170
box -8 -3 104 105
use FILL  FILL_8714
timestamp 1680363874
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_519
timestamp 1680363874
transform -1 0 2296 0 1 1170
box -9 -3 26 105
use FILL  FILL_8715
timestamp 1680363874
transform 1 0 2296 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6817
timestamp 1680363874
transform 1 0 2316 0 1 1175
box -3 -3 3 3
use FILL  FILL_8726
timestamp 1680363874
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_154
timestamp 1680363874
transform 1 0 2312 0 1 1170
box -8 -3 34 105
use AND2X2  AND2X2_57
timestamp 1680363874
transform -1 0 2376 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_58
timestamp 1680363874
transform -1 0 2408 0 1 1170
box -8 -3 40 105
use M3_M2  M3_M2_6818
timestamp 1680363874
transform 1 0 2444 0 1 1175
box -3 -3 3 3
use OAI21X1  OAI21X1_155
timestamp 1680363874
transform -1 0 2440 0 1 1170
box -8 -3 34 105
use FILL  FILL_8728
timestamp 1680363874
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_285
timestamp 1680363874
transform -1 0 2488 0 1 1170
box -8 -3 46 105
use FILL  FILL_8729
timestamp 1680363874
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6819
timestamp 1680363874
transform 1 0 2580 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_454
timestamp 1680363874
transform -1 0 2592 0 1 1170
box -8 -3 104 105
use FILL  FILL_8730
timestamp 1680363874
transform 1 0 2592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8750
timestamp 1680363874
transform 1 0 2600 0 1 1170
box -8 -3 16 105
use FILL  FILL_8752
timestamp 1680363874
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_8754
timestamp 1680363874
transform 1 0 2616 0 1 1170
box -8 -3 16 105
use FILL  FILL_8755
timestamp 1680363874
transform 1 0 2624 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6820
timestamp 1680363874
transform 1 0 2644 0 1 1175
box -3 -3 3 3
use FILL  FILL_8756
timestamp 1680363874
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use FILL  FILL_8757
timestamp 1680363874
transform 1 0 2640 0 1 1170
box -8 -3 16 105
use FILL  FILL_8758
timestamp 1680363874
transform 1 0 2648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8759
timestamp 1680363874
transform 1 0 2656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8760
timestamp 1680363874
transform 1 0 2664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8763
timestamp 1680363874
transform 1 0 2672 0 1 1170
box -8 -3 16 105
use AND2X2  AND2X2_59
timestamp 1680363874
transform -1 0 2712 0 1 1170
box -8 -3 40 105
use FILL  FILL_8764
timestamp 1680363874
transform 1 0 2712 0 1 1170
box -8 -3 16 105
use FILL  FILL_8765
timestamp 1680363874
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_8766
timestamp 1680363874
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_8767
timestamp 1680363874
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use FILL  FILL_8768
timestamp 1680363874
transform 1 0 2744 0 1 1170
box -8 -3 16 105
use AND2X2  AND2X2_60
timestamp 1680363874
transform 1 0 2752 0 1 1170
box -8 -3 40 105
use FILL  FILL_8769
timestamp 1680363874
transform 1 0 2784 0 1 1170
box -8 -3 16 105
use FILL  FILL_8770
timestamp 1680363874
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_8771
timestamp 1680363874
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_8777
timestamp 1680363874
transform 1 0 2808 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6821
timestamp 1680363874
transform 1 0 2844 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_287
timestamp 1680363874
transform 1 0 2816 0 1 1170
box -8 -3 46 105
use FILL  FILL_8779
timestamp 1680363874
transform 1 0 2856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8784
timestamp 1680363874
transform 1 0 2864 0 1 1170
box -8 -3 16 105
use FILL  FILL_8786
timestamp 1680363874
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use FILL  FILL_8788
timestamp 1680363874
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6822
timestamp 1680363874
transform 1 0 2900 0 1 1175
box -3 -3 3 3
use FILL  FILL_8789
timestamp 1680363874
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_8790
timestamp 1680363874
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_8791
timestamp 1680363874
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_8792
timestamp 1680363874
transform 1 0 2912 0 1 1170
box -8 -3 16 105
use FILL  FILL_8793
timestamp 1680363874
transform 1 0 2920 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_457
timestamp 1680363874
transform 1 0 2928 0 1 1170
box -8 -3 104 105
use FILL  FILL_8795
timestamp 1680363874
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_8796
timestamp 1680363874
transform 1 0 3032 0 1 1170
box -8 -3 16 105
use FILL  FILL_8797
timestamp 1680363874
transform 1 0 3040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8808
timestamp 1680363874
transform 1 0 3048 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_289
timestamp 1680363874
transform -1 0 3096 0 1 1170
box -8 -3 46 105
use FILL  FILL_8809
timestamp 1680363874
transform 1 0 3096 0 1 1170
box -8 -3 16 105
use FILL  FILL_8810
timestamp 1680363874
transform 1 0 3104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8811
timestamp 1680363874
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8812
timestamp 1680363874
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_8813
timestamp 1680363874
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_8814
timestamp 1680363874
transform 1 0 3136 0 1 1170
box -8 -3 16 105
use FILL  FILL_8815
timestamp 1680363874
transform 1 0 3144 0 1 1170
box -8 -3 16 105
use FILL  FILL_8816
timestamp 1680363874
transform 1 0 3152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8817
timestamp 1680363874
transform 1 0 3160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8818
timestamp 1680363874
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8819
timestamp 1680363874
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8820
timestamp 1680363874
transform 1 0 3184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8821
timestamp 1680363874
transform 1 0 3192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8822
timestamp 1680363874
transform 1 0 3200 0 1 1170
box -8 -3 16 105
use FILL  FILL_8823
timestamp 1680363874
transform 1 0 3208 0 1 1170
box -8 -3 16 105
use FILL  FILL_8824
timestamp 1680363874
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_8825
timestamp 1680363874
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_8826
timestamp 1680363874
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_8827
timestamp 1680363874
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_8828
timestamp 1680363874
transform 1 0 3248 0 1 1170
box -8 -3 16 105
use FILL  FILL_8833
timestamp 1680363874
transform 1 0 3256 0 1 1170
box -8 -3 16 105
use FILL  FILL_8835
timestamp 1680363874
transform 1 0 3264 0 1 1170
box -8 -3 16 105
use FILL  FILL_8837
timestamp 1680363874
transform 1 0 3272 0 1 1170
box -8 -3 16 105
use FILL  FILL_8839
timestamp 1680363874
transform 1 0 3280 0 1 1170
box -8 -3 16 105
use FILL  FILL_8840
timestamp 1680363874
transform 1 0 3288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8841
timestamp 1680363874
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8842
timestamp 1680363874
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_8845
timestamp 1680363874
transform 1 0 3312 0 1 1170
box -8 -3 16 105
use FILL  FILL_8847
timestamp 1680363874
transform 1 0 3320 0 1 1170
box -8 -3 16 105
use FILL  FILL_8849
timestamp 1680363874
transform 1 0 3328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8851
timestamp 1680363874
transform 1 0 3336 0 1 1170
box -8 -3 16 105
use FILL  FILL_8853
timestamp 1680363874
transform 1 0 3344 0 1 1170
box -8 -3 16 105
use FILL  FILL_8854
timestamp 1680363874
transform 1 0 3352 0 1 1170
box -8 -3 16 105
use FILL  FILL_8855
timestamp 1680363874
transform 1 0 3360 0 1 1170
box -8 -3 16 105
use FILL  FILL_8856
timestamp 1680363874
transform 1 0 3368 0 1 1170
box -8 -3 16 105
use FILL  FILL_8857
timestamp 1680363874
transform 1 0 3376 0 1 1170
box -8 -3 16 105
use FILL  FILL_8858
timestamp 1680363874
transform 1 0 3384 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_459
timestamp 1680363874
transform -1 0 3488 0 1 1170
box -8 -3 104 105
use FILL  FILL_8859
timestamp 1680363874
transform 1 0 3488 0 1 1170
box -8 -3 16 105
use AND2X2  AND2X2_61
timestamp 1680363874
transform 1 0 3496 0 1 1170
box -8 -3 40 105
use FILL  FILL_8860
timestamp 1680363874
transform 1 0 3528 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6823
timestamp 1680363874
transform 1 0 3548 0 1 1175
box -3 -3 3 3
use FILL  FILL_8861
timestamp 1680363874
transform 1 0 3536 0 1 1170
box -8 -3 16 105
use FILL  FILL_8862
timestamp 1680363874
transform 1 0 3544 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6824
timestamp 1680363874
transform 1 0 3564 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_291
timestamp 1680363874
transform 1 0 3552 0 1 1170
box -8 -3 46 105
use FILL  FILL_8863
timestamp 1680363874
transform 1 0 3592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8864
timestamp 1680363874
transform 1 0 3600 0 1 1170
box -8 -3 16 105
use FILL  FILL_8865
timestamp 1680363874
transform 1 0 3608 0 1 1170
box -8 -3 16 105
use FILL  FILL_8866
timestamp 1680363874
transform 1 0 3616 0 1 1170
box -8 -3 16 105
use FILL  FILL_8867
timestamp 1680363874
transform 1 0 3624 0 1 1170
box -8 -3 16 105
use FILL  FILL_8868
timestamp 1680363874
transform 1 0 3632 0 1 1170
box -8 -3 16 105
use FILL  FILL_8869
timestamp 1680363874
transform 1 0 3640 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_523
timestamp 1680363874
transform 1 0 3648 0 1 1170
box -9 -3 26 105
use FILL  FILL_8870
timestamp 1680363874
transform 1 0 3664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8871
timestamp 1680363874
transform 1 0 3672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8872
timestamp 1680363874
transform 1 0 3680 0 1 1170
box -8 -3 16 105
use FILL  FILL_8873
timestamp 1680363874
transform 1 0 3688 0 1 1170
box -8 -3 16 105
use FILL  FILL_8887
timestamp 1680363874
transform 1 0 3696 0 1 1170
box -8 -3 16 105
use FILL  FILL_8889
timestamp 1680363874
transform 1 0 3704 0 1 1170
box -8 -3 16 105
use FILL  FILL_8891
timestamp 1680363874
transform 1 0 3712 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_293
timestamp 1680363874
transform 1 0 3720 0 1 1170
box -8 -3 46 105
use FILL  FILL_8892
timestamp 1680363874
transform 1 0 3760 0 1 1170
box -8 -3 16 105
use FILL  FILL_8895
timestamp 1680363874
transform 1 0 3768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8897
timestamp 1680363874
transform 1 0 3776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8899
timestamp 1680363874
transform 1 0 3784 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_335
timestamp 1680363874
transform -1 0 3832 0 1 1170
box -8 -3 46 105
use FILL  FILL_8900
timestamp 1680363874
transform 1 0 3832 0 1 1170
box -8 -3 16 105
use FILL  FILL_8906
timestamp 1680363874
transform 1 0 3840 0 1 1170
box -8 -3 16 105
use FILL  FILL_8908
timestamp 1680363874
transform 1 0 3848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8910
timestamp 1680363874
transform 1 0 3856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8911
timestamp 1680363874
transform 1 0 3864 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_295
timestamp 1680363874
transform 1 0 3872 0 1 1170
box -8 -3 46 105
use INVX2  INVX2_527
timestamp 1680363874
transform 1 0 3912 0 1 1170
box -9 -3 26 105
use FILL  FILL_8912
timestamp 1680363874
transform 1 0 3928 0 1 1170
box -8 -3 16 105
use FILL  FILL_8918
timestamp 1680363874
transform 1 0 3936 0 1 1170
box -8 -3 16 105
use FILL  FILL_8919
timestamp 1680363874
transform 1 0 3944 0 1 1170
box -8 -3 16 105
use FILL  FILL_8920
timestamp 1680363874
transform 1 0 3952 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_461
timestamp 1680363874
transform -1 0 4056 0 1 1170
box -8 -3 104 105
use FILL  FILL_8921
timestamp 1680363874
transform 1 0 4056 0 1 1170
box -8 -3 16 105
use FILL  FILL_8931
timestamp 1680363874
transform 1 0 4064 0 1 1170
box -8 -3 16 105
use FILL  FILL_8932
timestamp 1680363874
transform 1 0 4072 0 1 1170
box -8 -3 16 105
use FILL  FILL_8933
timestamp 1680363874
transform 1 0 4080 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_529
timestamp 1680363874
transform 1 0 4088 0 1 1170
box -9 -3 26 105
use FILL  FILL_8934
timestamp 1680363874
transform 1 0 4104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8936
timestamp 1680363874
transform 1 0 4112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8938
timestamp 1680363874
transform 1 0 4120 0 1 1170
box -8 -3 16 105
use FILL  FILL_8940
timestamp 1680363874
transform 1 0 4128 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_298
timestamp 1680363874
transform 1 0 4136 0 1 1170
box -8 -3 46 105
use FILL  FILL_8942
timestamp 1680363874
transform 1 0 4176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8943
timestamp 1680363874
transform 1 0 4184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8946
timestamp 1680363874
transform 1 0 4192 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_338
timestamp 1680363874
transform 1 0 4200 0 1 1170
box -8 -3 46 105
use INVX2  INVX2_530
timestamp 1680363874
transform 1 0 4240 0 1 1170
box -9 -3 26 105
use FILL  FILL_8948
timestamp 1680363874
transform 1 0 4256 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_462
timestamp 1680363874
transform -1 0 4360 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_463
timestamp 1680363874
transform 1 0 4360 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_531
timestamp 1680363874
transform -1 0 4472 0 1 1170
box -9 -3 26 105
use FILL  FILL_8949
timestamp 1680363874
transform 1 0 4472 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6825
timestamp 1680363874
transform 1 0 4508 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_299
timestamp 1680363874
transform -1 0 4520 0 1 1170
box -8 -3 46 105
use FILL  FILL_8950
timestamp 1680363874
transform 1 0 4520 0 1 1170
box -8 -3 16 105
use FILL  FILL_8973
timestamp 1680363874
transform 1 0 4528 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6826
timestamp 1680363874
transform 1 0 4572 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_339
timestamp 1680363874
transform 1 0 4536 0 1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_465
timestamp 1680363874
transform -1 0 4672 0 1 1170
box -8 -3 104 105
use FILL  FILL_8974
timestamp 1680363874
transform 1 0 4672 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_534
timestamp 1680363874
transform 1 0 4680 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_466
timestamp 1680363874
transform -1 0 4792 0 1 1170
box -8 -3 104 105
use FILL  FILL_8987
timestamp 1680363874
transform 1 0 4792 0 1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_71
timestamp 1680363874
transform 1 0 4827 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_6835
timestamp 1680363874
transform 1 0 116 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7502
timestamp 1680363874
transform 1 0 92 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7598
timestamp 1680363874
transform 1 0 116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7599
timestamp 1680363874
transform 1 0 180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7600
timestamp 1680363874
transform 1 0 188 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6914
timestamp 1680363874
transform 1 0 188 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7503
timestamp 1680363874
transform 1 0 276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7601
timestamp 1680363874
transform 1 0 252 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7504
timestamp 1680363874
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6915
timestamp 1680363874
transform 1 0 292 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7496
timestamp 1680363874
transform 1 0 324 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6853
timestamp 1680363874
transform 1 0 332 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6854
timestamp 1680363874
transform 1 0 356 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6878
timestamp 1680363874
transform 1 0 348 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7505
timestamp 1680363874
transform 1 0 356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7602
timestamp 1680363874
transform 1 0 348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7603
timestamp 1680363874
transform 1 0 356 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6916
timestamp 1680363874
transform 1 0 356 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6956
timestamp 1680363874
transform 1 0 348 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7497
timestamp 1680363874
transform 1 0 388 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6836
timestamp 1680363874
transform 1 0 404 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7506
timestamp 1680363874
transform 1 0 404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7604
timestamp 1680363874
transform 1 0 396 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6957
timestamp 1680363874
transform 1 0 396 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7507
timestamp 1680363874
transform 1 0 420 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6879
timestamp 1680363874
transform 1 0 460 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7699
timestamp 1680363874
transform 1 0 452 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7508
timestamp 1680363874
transform 1 0 476 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6995
timestamp 1680363874
transform 1 0 476 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6837
timestamp 1680363874
transform 1 0 540 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7509
timestamp 1680363874
transform 1 0 492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7605
timestamp 1680363874
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6996
timestamp 1680363874
transform 1 0 500 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7606
timestamp 1680363874
transform 1 0 580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7700
timestamp 1680363874
transform 1 0 596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7510
timestamp 1680363874
transform 1 0 604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7498
timestamp 1680363874
transform 1 0 636 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7607
timestamp 1680363874
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6890
timestamp 1680363874
transform 1 0 628 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7511
timestamp 1680363874
transform 1 0 644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7512
timestamp 1680363874
transform 1 0 668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7513
timestamp 1680363874
transform 1 0 692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7701
timestamp 1680363874
transform 1 0 684 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7514
timestamp 1680363874
transform 1 0 716 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6891
timestamp 1680363874
transform 1 0 700 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7608
timestamp 1680363874
transform 1 0 708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7515
timestamp 1680363874
transform 1 0 756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7609
timestamp 1680363874
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7610
timestamp 1680363874
transform 1 0 836 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6855
timestamp 1680363874
transform 1 0 884 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7516
timestamp 1680363874
transform 1 0 924 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6880
timestamp 1680363874
transform 1 0 972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6838
timestamp 1680363874
transform 1 0 1020 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6839
timestamp 1680363874
transform 1 0 1044 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6856
timestamp 1680363874
transform 1 0 1036 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6857
timestamp 1680363874
transform 1 0 1068 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7517
timestamp 1680363874
transform 1 0 1020 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6881
timestamp 1680363874
transform 1 0 1084 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7611
timestamp 1680363874
transform 1 0 972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7612
timestamp 1680363874
transform 1 0 1004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7613
timestamp 1680363874
transform 1 0 1068 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6840
timestamp 1680363874
transform 1 0 1116 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6841
timestamp 1680363874
transform 1 0 1132 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7518
timestamp 1680363874
transform 1 0 1132 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6858
timestamp 1680363874
transform 1 0 1156 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6859
timestamp 1680363874
transform 1 0 1180 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7519
timestamp 1680363874
transform 1 0 1156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7520
timestamp 1680363874
transform 1 0 1172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7521
timestamp 1680363874
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7614
timestamp 1680363874
transform 1 0 1132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6892
timestamp 1680363874
transform 1 0 1140 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7615
timestamp 1680363874
transform 1 0 1148 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6917
timestamp 1680363874
transform 1 0 1140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6893
timestamp 1680363874
transform 1 0 1180 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7616
timestamp 1680363874
transform 1 0 1188 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6958
timestamp 1680363874
transform 1 0 1172 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6894
timestamp 1680363874
transform 1 0 1196 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6918
timestamp 1680363874
transform 1 0 1204 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7617
timestamp 1680363874
transform 1 0 1212 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6860
timestamp 1680363874
transform 1 0 1228 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7618
timestamp 1680363874
transform 1 0 1236 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6919
timestamp 1680363874
transform 1 0 1236 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6959
timestamp 1680363874
transform 1 0 1236 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6997
timestamp 1680363874
transform 1 0 1236 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7522
timestamp 1680363874
transform 1 0 1268 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6979
timestamp 1680363874
transform 1 0 1260 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6842
timestamp 1680363874
transform 1 0 1284 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7619
timestamp 1680363874
transform 1 0 1284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6895
timestamp 1680363874
transform 1 0 1292 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7620
timestamp 1680363874
transform 1 0 1300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7702
timestamp 1680363874
transform 1 0 1292 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6920
timestamp 1680363874
transform 1 0 1300 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6960
timestamp 1680363874
transform 1 0 1292 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7706
timestamp 1680363874
transform 1 0 1308 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6980
timestamp 1680363874
transform 1 0 1292 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7703
timestamp 1680363874
transform 1 0 1324 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6961
timestamp 1680363874
transform 1 0 1332 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7523
timestamp 1680363874
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7524
timestamp 1680363874
transform 1 0 1452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7621
timestamp 1680363874
transform 1 0 1404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7622
timestamp 1680363874
transform 1 0 1436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7623
timestamp 1680363874
transform 1 0 1444 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6921
timestamp 1680363874
transform 1 0 1404 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6981
timestamp 1680363874
transform 1 0 1444 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6998
timestamp 1680363874
transform 1 0 1452 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7525
timestamp 1680363874
transform 1 0 1492 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6922
timestamp 1680363874
transform 1 0 1484 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7526
timestamp 1680363874
transform 1 0 1524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7527
timestamp 1680363874
transform 1 0 1540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7624
timestamp 1680363874
transform 1 0 1532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7625
timestamp 1680363874
transform 1 0 1580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7528
timestamp 1680363874
transform 1 0 1596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7529
timestamp 1680363874
transform 1 0 1620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7626
timestamp 1680363874
transform 1 0 1604 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6827
timestamp 1680363874
transform 1 0 1636 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7627
timestamp 1680363874
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6982
timestamp 1680363874
transform 1 0 1644 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6861
timestamp 1680363874
transform 1 0 1708 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7530
timestamp 1680363874
transform 1 0 1660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7531
timestamp 1680363874
transform 1 0 1668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7532
timestamp 1680363874
transform 1 0 1684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7533
timestamp 1680363874
transform 1 0 1700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7628
timestamp 1680363874
transform 1 0 1676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7629
timestamp 1680363874
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6923
timestamp 1680363874
transform 1 0 1668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6924
timestamp 1680363874
transform 1 0 1724 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6828
timestamp 1680363874
transform 1 0 1764 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6843
timestamp 1680363874
transform 1 0 1756 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7534
timestamp 1680363874
transform 1 0 1748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7535
timestamp 1680363874
transform 1 0 1764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7536
timestamp 1680363874
transform 1 0 1780 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6925
timestamp 1680363874
transform 1 0 1740 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7630
timestamp 1680363874
transform 1 0 1772 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6926
timestamp 1680363874
transform 1 0 1772 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7631
timestamp 1680363874
transform 1 0 1788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7537
timestamp 1680363874
transform 1 0 1804 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6962
timestamp 1680363874
transform 1 0 1820 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6963
timestamp 1680363874
transform 1 0 1844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6983
timestamp 1680363874
transform 1 0 1844 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6862
timestamp 1680363874
transform 1 0 1868 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7538
timestamp 1680363874
transform 1 0 1868 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6896
timestamp 1680363874
transform 1 0 1892 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7632
timestamp 1680363874
transform 1 0 1916 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6927
timestamp 1680363874
transform 1 0 1916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6863
timestamp 1680363874
transform 1 0 1956 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6897
timestamp 1680363874
transform 1 0 2028 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7704
timestamp 1680363874
transform 1 0 2020 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6928
timestamp 1680363874
transform 1 0 2028 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7633
timestamp 1680363874
transform 1 0 2052 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6999
timestamp 1680363874
transform 1 0 2044 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6898
timestamp 1680363874
transform 1 0 2060 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6864
timestamp 1680363874
transform 1 0 2076 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7539
timestamp 1680363874
transform 1 0 2100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7634
timestamp 1680363874
transform 1 0 2092 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6899
timestamp 1680363874
transform 1 0 2100 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7540
timestamp 1680363874
transform 1 0 2116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7635
timestamp 1680363874
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7499
timestamp 1680363874
transform 1 0 2188 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6964
timestamp 1680363874
transform 1 0 2180 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7541
timestamp 1680363874
transform 1 0 2212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7636
timestamp 1680363874
transform 1 0 2204 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6984
timestamp 1680363874
transform 1 0 2212 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7500
timestamp 1680363874
transform 1 0 2236 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6900
timestamp 1680363874
transform 1 0 2236 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6929
timestamp 1680363874
transform 1 0 2236 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7637
timestamp 1680363874
transform 1 0 2268 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6930
timestamp 1680363874
transform 1 0 2260 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6829
timestamp 1680363874
transform 1 0 2420 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6865
timestamp 1680363874
transform 1 0 2372 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6866
timestamp 1680363874
transform 1 0 2420 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7542
timestamp 1680363874
transform 1 0 2420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7638
timestamp 1680363874
transform 1 0 2340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7639
timestamp 1680363874
transform 1 0 2396 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6931
timestamp 1680363874
transform 1 0 2396 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6965
timestamp 1680363874
transform 1 0 2372 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6966
timestamp 1680363874
transform 1 0 2420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6985
timestamp 1680363874
transform 1 0 2404 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7000
timestamp 1680363874
transform 1 0 2380 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7543
timestamp 1680363874
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6967
timestamp 1680363874
transform 1 0 2452 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6932
timestamp 1680363874
transform 1 0 2468 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6830
timestamp 1680363874
transform 1 0 2484 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7640
timestamp 1680363874
transform 1 0 2500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6933
timestamp 1680363874
transform 1 0 2492 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7641
timestamp 1680363874
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6831
timestamp 1680363874
transform 1 0 2564 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7501
timestamp 1680363874
transform 1 0 2564 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6867
timestamp 1680363874
transform 1 0 2588 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7642
timestamp 1680363874
transform 1 0 2604 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6968
timestamp 1680363874
transform 1 0 2604 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7544
timestamp 1680363874
transform 1 0 2628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7545
timestamp 1680363874
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7643
timestamp 1680363874
transform 1 0 2644 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6934
timestamp 1680363874
transform 1 0 2636 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7546
timestamp 1680363874
transform 1 0 2676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7644
timestamp 1680363874
transform 1 0 2684 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6844
timestamp 1680363874
transform 1 0 2716 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6845
timestamp 1680363874
transform 1 0 2796 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7547
timestamp 1680363874
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7645
timestamp 1680363874
transform 1 0 2764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7646
timestamp 1680363874
transform 1 0 2796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7647
timestamp 1680363874
transform 1 0 2804 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6935
timestamp 1680363874
transform 1 0 2716 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6936
timestamp 1680363874
transform 1 0 2748 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6937
timestamp 1680363874
transform 1 0 2764 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6938
timestamp 1680363874
transform 1 0 2804 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7648
timestamp 1680363874
transform 1 0 2844 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6846
timestamp 1680363874
transform 1 0 2908 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7548
timestamp 1680363874
transform 1 0 2884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7549
timestamp 1680363874
transform 1 0 2892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7550
timestamp 1680363874
transform 1 0 2908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7551
timestamp 1680363874
transform 1 0 2916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7649
timestamp 1680363874
transform 1 0 2900 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6868
timestamp 1680363874
transform 1 0 2932 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7650
timestamp 1680363874
transform 1 0 2948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7552
timestamp 1680363874
transform 1 0 2988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7553
timestamp 1680363874
transform 1 0 3020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7651
timestamp 1680363874
transform 1 0 3012 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6901
timestamp 1680363874
transform 1 0 3020 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7652
timestamp 1680363874
transform 1 0 3028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6939
timestamp 1680363874
transform 1 0 3012 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6986
timestamp 1680363874
transform 1 0 3028 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7554
timestamp 1680363874
transform 1 0 3060 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6902
timestamp 1680363874
transform 1 0 3060 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7555
timestamp 1680363874
transform 1 0 3068 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6832
timestamp 1680363874
transform 1 0 3092 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6869
timestamp 1680363874
transform 1 0 3124 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6870
timestamp 1680363874
transform 1 0 3148 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7556
timestamp 1680363874
transform 1 0 3092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7557
timestamp 1680363874
transform 1 0 3108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7558
timestamp 1680363874
transform 1 0 3124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7653
timestamp 1680363874
transform 1 0 3084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7654
timestamp 1680363874
transform 1 0 3100 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6940
timestamp 1680363874
transform 1 0 3084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6987
timestamp 1680363874
transform 1 0 3100 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6882
timestamp 1680363874
transform 1 0 3172 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7559
timestamp 1680363874
transform 1 0 3212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7560
timestamp 1680363874
transform 1 0 3236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7561
timestamp 1680363874
transform 1 0 3244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7655
timestamp 1680363874
transform 1 0 3172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7656
timestamp 1680363874
transform 1 0 3204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7657
timestamp 1680363874
transform 1 0 3212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7658
timestamp 1680363874
transform 1 0 3228 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6941
timestamp 1680363874
transform 1 0 3228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6969
timestamp 1680363874
transform 1 0 3156 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6970
timestamp 1680363874
transform 1 0 3212 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6988
timestamp 1680363874
transform 1 0 3140 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6989
timestamp 1680363874
transform 1 0 3220 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6883
timestamp 1680363874
transform 1 0 3252 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7659
timestamp 1680363874
transform 1 0 3252 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6903
timestamp 1680363874
transform 1 0 3268 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7562
timestamp 1680363874
transform 1 0 3300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7660
timestamp 1680363874
transform 1 0 3308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6942
timestamp 1680363874
transform 1 0 3300 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6847
timestamp 1680363874
transform 1 0 3348 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7563
timestamp 1680363874
transform 1 0 3348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7564
timestamp 1680363874
transform 1 0 3364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7661
timestamp 1680363874
transform 1 0 3372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6943
timestamp 1680363874
transform 1 0 3372 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6833
timestamp 1680363874
transform 1 0 3420 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7565
timestamp 1680363874
transform 1 0 3420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7662
timestamp 1680363874
transform 1 0 3444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7566
timestamp 1680363874
transform 1 0 3468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7567
timestamp 1680363874
transform 1 0 3476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7568
timestamp 1680363874
transform 1 0 3492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7663
timestamp 1680363874
transform 1 0 3460 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6944
timestamp 1680363874
transform 1 0 3452 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6904
timestamp 1680363874
transform 1 0 3468 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7664
timestamp 1680363874
transform 1 0 3500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6945
timestamp 1680363874
transform 1 0 3500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6971
timestamp 1680363874
transform 1 0 3484 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6848
timestamp 1680363874
transform 1 0 3540 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6849
timestamp 1680363874
transform 1 0 3564 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6871
timestamp 1680363874
transform 1 0 3532 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6884
timestamp 1680363874
transform 1 0 3524 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6834
timestamp 1680363874
transform 1 0 3580 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7569
timestamp 1680363874
transform 1 0 3532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7570
timestamp 1680363874
transform 1 0 3540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7571
timestamp 1680363874
transform 1 0 3556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7572
timestamp 1680363874
transform 1 0 3564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7665
timestamp 1680363874
transform 1 0 3516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7001
timestamp 1680363874
transform 1 0 3524 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6905
timestamp 1680363874
transform 1 0 3540 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7666
timestamp 1680363874
transform 1 0 3548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6972
timestamp 1680363874
transform 1 0 3548 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6885
timestamp 1680363874
transform 1 0 3572 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6872
timestamp 1680363874
transform 1 0 3596 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7573
timestamp 1680363874
transform 1 0 3580 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6906
timestamp 1680363874
transform 1 0 3580 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7574
timestamp 1680363874
transform 1 0 3676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7667
timestamp 1680363874
transform 1 0 3588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7668
timestamp 1680363874
transform 1 0 3596 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6907
timestamp 1680363874
transform 1 0 3612 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7669
timestamp 1680363874
transform 1 0 3628 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6946
timestamp 1680363874
transform 1 0 3588 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6947
timestamp 1680363874
transform 1 0 3628 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6850
timestamp 1680363874
transform 1 0 3692 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7670
timestamp 1680363874
transform 1 0 3692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6973
timestamp 1680363874
transform 1 0 3692 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6990
timestamp 1680363874
transform 1 0 3644 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6991
timestamp 1680363874
transform 1 0 3684 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7575
timestamp 1680363874
transform 1 0 3708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7576
timestamp 1680363874
transform 1 0 3740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7577
timestamp 1680363874
transform 1 0 3748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7671
timestamp 1680363874
transform 1 0 3732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7672
timestamp 1680363874
transform 1 0 3748 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6948
timestamp 1680363874
transform 1 0 3748 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6992
timestamp 1680363874
transform 1 0 3740 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7002
timestamp 1680363874
transform 1 0 3748 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6993
timestamp 1680363874
transform 1 0 3764 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7673
timestamp 1680363874
transform 1 0 3836 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6994
timestamp 1680363874
transform 1 0 3828 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6851
timestamp 1680363874
transform 1 0 3852 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7578
timestamp 1680363874
transform 1 0 3868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7579
timestamp 1680363874
transform 1 0 3884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7580
timestamp 1680363874
transform 1 0 3900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7674
timestamp 1680363874
transform 1 0 3876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7675
timestamp 1680363874
transform 1 0 3892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7676
timestamp 1680363874
transform 1 0 3908 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6949
timestamp 1680363874
transform 1 0 3908 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6852
timestamp 1680363874
transform 1 0 3972 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6873
timestamp 1680363874
transform 1 0 3964 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6874
timestamp 1680363874
transform 1 0 3980 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6886
timestamp 1680363874
transform 1 0 3948 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7581
timestamp 1680363874
transform 1 0 3972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7582
timestamp 1680363874
transform 1 0 3980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7677
timestamp 1680363874
transform 1 0 3948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7678
timestamp 1680363874
transform 1 0 3964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7679
timestamp 1680363874
transform 1 0 3980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7680
timestamp 1680363874
transform 1 0 3988 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6950
timestamp 1680363874
transform 1 0 3956 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6951
timestamp 1680363874
transform 1 0 3988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6974
timestamp 1680363874
transform 1 0 3980 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7681
timestamp 1680363874
transform 1 0 4044 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6975
timestamp 1680363874
transform 1 0 4044 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7583
timestamp 1680363874
transform 1 0 4068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7584
timestamp 1680363874
transform 1 0 4092 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6908
timestamp 1680363874
transform 1 0 4068 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6887
timestamp 1680363874
transform 1 0 4100 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7682
timestamp 1680363874
transform 1 0 4084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7683
timestamp 1680363874
transform 1 0 4100 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6909
timestamp 1680363874
transform 1 0 4108 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6976
timestamp 1680363874
transform 1 0 4116 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6875
timestamp 1680363874
transform 1 0 4156 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7585
timestamp 1680363874
transform 1 0 4164 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6888
timestamp 1680363874
transform 1 0 4172 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7586
timestamp 1680363874
transform 1 0 4180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7684
timestamp 1680363874
transform 1 0 4148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7685
timestamp 1680363874
transform 1 0 4172 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6910
timestamp 1680363874
transform 1 0 4180 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6952
timestamp 1680363874
transform 1 0 4172 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6889
timestamp 1680363874
transform 1 0 4220 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7686
timestamp 1680363874
transform 1 0 4220 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6953
timestamp 1680363874
transform 1 0 4228 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7587
timestamp 1680363874
transform 1 0 4236 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6876
timestamp 1680363874
transform 1 0 4268 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7588
timestamp 1680363874
transform 1 0 4268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7589
timestamp 1680363874
transform 1 0 4292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7687
timestamp 1680363874
transform 1 0 4244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7688
timestamp 1680363874
transform 1 0 4260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7689
timestamp 1680363874
transform 1 0 4276 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7690
timestamp 1680363874
transform 1 0 4284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6977
timestamp 1680363874
transform 1 0 4244 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6911
timestamp 1680363874
transform 1 0 4292 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7003
timestamp 1680363874
transform 1 0 4308 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7590
timestamp 1680363874
transform 1 0 4356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7691
timestamp 1680363874
transform 1 0 4388 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7004
timestamp 1680363874
transform 1 0 4348 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7591
timestamp 1680363874
transform 1 0 4460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7705
timestamp 1680363874
transform 1 0 4476 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7692
timestamp 1680363874
transform 1 0 4492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7592
timestamp 1680363874
transform 1 0 4516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7693
timestamp 1680363874
transform 1 0 4572 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6877
timestamp 1680363874
transform 1 0 4612 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7593
timestamp 1680363874
transform 1 0 4612 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6954
timestamp 1680363874
transform 1 0 4628 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7594
timestamp 1680363874
transform 1 0 4644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7595
timestamp 1680363874
transform 1 0 4660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7596
timestamp 1680363874
transform 1 0 4668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7694
timestamp 1680363874
transform 1 0 4652 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6912
timestamp 1680363874
transform 1 0 4660 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7695
timestamp 1680363874
transform 1 0 4668 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6955
timestamp 1680363874
transform 1 0 4652 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6913
timestamp 1680363874
transform 1 0 4676 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7597
timestamp 1680363874
transform 1 0 4780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7696
timestamp 1680363874
transform 1 0 4692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7697
timestamp 1680363874
transform 1 0 4700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7698
timestamp 1680363874
transform 1 0 4740 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6978
timestamp 1680363874
transform 1 0 4668 0 1 1105
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_72
timestamp 1680363874
transform 1 0 24 0 1 1070
box -10 -3 10 3
use FILL  FILL_8519
timestamp 1680363874
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_437
timestamp 1680363874
transform 1 0 80 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8524
timestamp 1680363874
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8527
timestamp 1680363874
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_439
timestamp 1680363874
transform -1 0 288 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8528
timestamp 1680363874
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8530
timestamp 1680363874
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8534
timestamp 1680363874
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8535
timestamp 1680363874
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use OR2X1  OR2X1_1
timestamp 1680363874
transform 1 0 320 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8536
timestamp 1680363874
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8537
timestamp 1680363874
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_101
timestamp 1680363874
transform -1 0 392 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8538
timestamp 1680363874
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8539
timestamp 1680363874
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8540
timestamp 1680363874
transform 1 0 408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8541
timestamp 1680363874
transform 1 0 416 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_150
timestamp 1680363874
transform 1 0 424 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8542
timestamp 1680363874
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8543
timestamp 1680363874
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8544
timestamp 1680363874
transform 1 0 472 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_441
timestamp 1680363874
transform 1 0 480 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8555
timestamp 1680363874
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8556
timestamp 1680363874
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8557
timestamp 1680363874
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_152
timestamp 1680363874
transform -1 0 632 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8558
timestamp 1680363874
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8560
timestamp 1680363874
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8562
timestamp 1680363874
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8564
timestamp 1680363874
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_53
timestamp 1680363874
transform 1 0 664 0 -1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_153
timestamp 1680363874
transform -1 0 720 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8570
timestamp 1680363874
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8574
timestamp 1680363874
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8575
timestamp 1680363874
transform 1 0 736 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_443
timestamp 1680363874
transform 1 0 744 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8576
timestamp 1680363874
transform 1 0 840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8577
timestamp 1680363874
transform 1 0 848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8578
timestamp 1680363874
transform 1 0 856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8579
timestamp 1680363874
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8580
timestamp 1680363874
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8581
timestamp 1680363874
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8582
timestamp 1680363874
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8583
timestamp 1680363874
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8585
timestamp 1680363874
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_445
timestamp 1680363874
transform 1 0 912 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_446
timestamp 1680363874
transform 1 0 1008 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_514
timestamp 1680363874
transform 1 0 1104 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8594
timestamp 1680363874
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8603
timestamp 1680363874
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_325
timestamp 1680363874
transform -1 0 1176 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8604
timestamp 1680363874
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8605
timestamp 1680363874
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8606
timestamp 1680363874
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8607
timestamp 1680363874
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8608
timestamp 1680363874
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_281
timestamp 1680363874
transform -1 0 1256 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8609
timestamp 1680363874
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8610
timestamp 1680363874
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8611
timestamp 1680363874
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8612
timestamp 1680363874
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_63
timestamp 1680363874
transform 1 0 1288 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8613
timestamp 1680363874
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8617
timestamp 1680363874
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8618
timestamp 1680363874
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_449
timestamp 1680363874
transform 1 0 1344 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8619
timestamp 1680363874
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8620
timestamp 1680363874
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8621
timestamp 1680363874
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8622
timestamp 1680363874
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8623
timestamp 1680363874
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8624
timestamp 1680363874
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8626
timestamp 1680363874
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8628
timestamp 1680363874
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_327
timestamp 1680363874
transform 1 0 1504 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8633
timestamp 1680363874
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8635
timestamp 1680363874
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8637
timestamp 1680363874
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8639
timestamp 1680363874
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8641
timestamp 1680363874
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_282
timestamp 1680363874
transform 1 0 1584 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8648
timestamp 1680363874
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8650
timestamp 1680363874
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8652
timestamp 1680363874
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8659
timestamp 1680363874
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8660
timestamp 1680363874
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_328
timestamp 1680363874
transform -1 0 1704 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8661
timestamp 1680363874
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8663
timestamp 1680363874
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8665
timestamp 1680363874
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8669
timestamp 1680363874
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8670
timestamp 1680363874
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_329
timestamp 1680363874
transform 1 0 1744 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8671
timestamp 1680363874
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8673
timestamp 1680363874
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8674
timestamp 1680363874
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_517
timestamp 1680363874
transform 1 0 1808 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8675
timestamp 1680363874
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8677
timestamp 1680363874
transform 1 0 1832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8679
timestamp 1680363874
transform 1 0 1840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8681
timestamp 1680363874
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_451
timestamp 1680363874
transform 1 0 1856 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8685
timestamp 1680363874
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8686
timestamp 1680363874
transform 1 0 1960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8687
timestamp 1680363874
transform 1 0 1968 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_518
timestamp 1680363874
transform 1 0 1976 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8691
timestamp 1680363874
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8692
timestamp 1680363874
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8693
timestamp 1680363874
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8694
timestamp 1680363874
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8695
timestamp 1680363874
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8696
timestamp 1680363874
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8698
timestamp 1680363874
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8700
timestamp 1680363874
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8702
timestamp 1680363874
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8704
timestamp 1680363874
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_284
timestamp 1680363874
transform -1 0 2112 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8705
timestamp 1680363874
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8706
timestamp 1680363874
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8707
timestamp 1680363874
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8708
timestamp 1680363874
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8709
timestamp 1680363874
transform 1 0 2144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8710
timestamp 1680363874
transform 1 0 2152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8711
timestamp 1680363874
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8713
timestamp 1680363874
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8716
timestamp 1680363874
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_102
timestamp 1680363874
transform 1 0 2184 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8717
timestamp 1680363874
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8718
timestamp 1680363874
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8719
timestamp 1680363874
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_103
timestamp 1680363874
transform 1 0 2232 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8720
timestamp 1680363874
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8721
timestamp 1680363874
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8722
timestamp 1680363874
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8723
timestamp 1680363874
transform 1 0 2280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8724
timestamp 1680363874
transform 1 0 2288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8725
timestamp 1680363874
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8727
timestamp 1680363874
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8731
timestamp 1680363874
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8732
timestamp 1680363874
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8733
timestamp 1680363874
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_455
timestamp 1680363874
transform -1 0 2432 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8734
timestamp 1680363874
transform 1 0 2432 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7005
timestamp 1680363874
transform 1 0 2452 0 1 1075
box -3 -3 3 3
use FILL  FILL_8735
timestamp 1680363874
transform 1 0 2440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8736
timestamp 1680363874
transform 1 0 2448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8737
timestamp 1680363874
transform 1 0 2456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8738
timestamp 1680363874
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8739
timestamp 1680363874
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8740
timestamp 1680363874
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8741
timestamp 1680363874
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8742
timestamp 1680363874
transform 1 0 2496 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_104
timestamp 1680363874
transform -1 0 2528 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8743
timestamp 1680363874
transform 1 0 2528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8744
timestamp 1680363874
transform 1 0 2536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8745
timestamp 1680363874
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8746
timestamp 1680363874
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8747
timestamp 1680363874
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_520
timestamp 1680363874
transform -1 0 2584 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8748
timestamp 1680363874
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8749
timestamp 1680363874
transform 1 0 2592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8751
timestamp 1680363874
transform 1 0 2600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8753
timestamp 1680363874
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8761
timestamp 1680363874
transform 1 0 2616 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_286
timestamp 1680363874
transform -1 0 2664 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8762
timestamp 1680363874
transform 1 0 2664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8772
timestamp 1680363874
transform 1 0 2672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8773
timestamp 1680363874
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8774
timestamp 1680363874
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8775
timestamp 1680363874
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_456
timestamp 1680363874
transform 1 0 2704 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8776
timestamp 1680363874
transform 1 0 2800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8778
timestamp 1680363874
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8780
timestamp 1680363874
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8781
timestamp 1680363874
transform 1 0 2824 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_521
timestamp 1680363874
transform -1 0 2848 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8782
timestamp 1680363874
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8783
timestamp 1680363874
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8785
timestamp 1680363874
transform 1 0 2864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8787
timestamp 1680363874
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_288
timestamp 1680363874
transform 1 0 2880 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8794
timestamp 1680363874
transform 1 0 2920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8798
timestamp 1680363874
transform 1 0 2928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8799
timestamp 1680363874
transform 1 0 2936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8800
timestamp 1680363874
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7006
timestamp 1680363874
transform 1 0 2964 0 1 1075
box -3 -3 3 3
use FILL  FILL_8801
timestamp 1680363874
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8802
timestamp 1680363874
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8803
timestamp 1680363874
transform 1 0 2968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8804
timestamp 1680363874
transform 1 0 2976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8805
timestamp 1680363874
transform 1 0 2984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8806
timestamp 1680363874
transform 1 0 2992 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_331
timestamp 1680363874
transform -1 0 3040 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8807
timestamp 1680363874
transform 1 0 3040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8829
timestamp 1680363874
transform 1 0 3048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8830
timestamp 1680363874
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8831
timestamp 1680363874
transform 1 0 3064 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_332
timestamp 1680363874
transform -1 0 3112 0 -1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_458
timestamp 1680363874
transform 1 0 3112 0 -1 1170
box -8 -3 104 105
use AOI22X1  AOI22X1_290
timestamp 1680363874
transform -1 0 3248 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8832
timestamp 1680363874
transform 1 0 3248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8834
timestamp 1680363874
transform 1 0 3256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8836
timestamp 1680363874
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8838
timestamp 1680363874
transform 1 0 3272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8843
timestamp 1680363874
transform 1 0 3280 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7007
timestamp 1680363874
transform 1 0 3300 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_522
timestamp 1680363874
transform -1 0 3304 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8844
timestamp 1680363874
transform 1 0 3304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8846
timestamp 1680363874
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8848
timestamp 1680363874
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8850
timestamp 1680363874
transform 1 0 3328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8852
timestamp 1680363874
transform 1 0 3336 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_333
timestamp 1680363874
transform 1 0 3344 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8874
timestamp 1680363874
transform 1 0 3384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8875
timestamp 1680363874
transform 1 0 3392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8876
timestamp 1680363874
transform 1 0 3400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8877
timestamp 1680363874
transform 1 0 3408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8878
timestamp 1680363874
transform 1 0 3416 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_524
timestamp 1680363874
transform -1 0 3440 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8879
timestamp 1680363874
transform 1 0 3440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8880
timestamp 1680363874
transform 1 0 3448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8881
timestamp 1680363874
transform 1 0 3456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8882
timestamp 1680363874
transform 1 0 3464 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_334
timestamp 1680363874
transform 1 0 3472 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8883
timestamp 1680363874
transform 1 0 3512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8884
timestamp 1680363874
transform 1 0 3520 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_292
timestamp 1680363874
transform -1 0 3568 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8885
timestamp 1680363874
transform 1 0 3568 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_525
timestamp 1680363874
transform 1 0 3576 0 -1 1170
box -9 -3 26 105
use M3_M2  M3_M2_7008
timestamp 1680363874
transform 1 0 3676 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_460
timestamp 1680363874
transform -1 0 3688 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8886
timestamp 1680363874
transform 1 0 3688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8888
timestamp 1680363874
transform 1 0 3696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8890
timestamp 1680363874
transform 1 0 3704 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7009
timestamp 1680363874
transform 1 0 3748 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_294
timestamp 1680363874
transform 1 0 3712 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8893
timestamp 1680363874
transform 1 0 3752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8894
timestamp 1680363874
transform 1 0 3760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8896
timestamp 1680363874
transform 1 0 3768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8898
timestamp 1680363874
transform 1 0 3776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8901
timestamp 1680363874
transform 1 0 3784 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_526
timestamp 1680363874
transform 1 0 3792 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8902
timestamp 1680363874
transform 1 0 3808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8903
timestamp 1680363874
transform 1 0 3816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8904
timestamp 1680363874
transform 1 0 3824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8905
timestamp 1680363874
transform 1 0 3832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8907
timestamp 1680363874
transform 1 0 3840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8909
timestamp 1680363874
transform 1 0 3848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8913
timestamp 1680363874
transform 1 0 3856 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_336
timestamp 1680363874
transform -1 0 3904 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8914
timestamp 1680363874
transform 1 0 3904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8915
timestamp 1680363874
transform 1 0 3912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8916
timestamp 1680363874
transform 1 0 3920 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7010
timestamp 1680363874
transform 1 0 3940 0 1 1075
box -3 -3 3 3
use FILL  FILL_8917
timestamp 1680363874
transform 1 0 3928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8922
timestamp 1680363874
transform 1 0 3936 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_296
timestamp 1680363874
transform -1 0 3984 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8923
timestamp 1680363874
transform 1 0 3984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8924
timestamp 1680363874
transform 1 0 3992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8925
timestamp 1680363874
transform 1 0 4000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8926
timestamp 1680363874
transform 1 0 4008 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_528
timestamp 1680363874
transform 1 0 4016 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8927
timestamp 1680363874
transform 1 0 4032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8928
timestamp 1680363874
transform 1 0 4040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8929
timestamp 1680363874
transform 1 0 4048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8930
timestamp 1680363874
transform 1 0 4056 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_297
timestamp 1680363874
transform 1 0 4064 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8935
timestamp 1680363874
transform 1 0 4104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8937
timestamp 1680363874
transform 1 0 4112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8939
timestamp 1680363874
transform 1 0 4120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8941
timestamp 1680363874
transform 1 0 4128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8944
timestamp 1680363874
transform 1 0 4136 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_337
timestamp 1680363874
transform 1 0 4144 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8945
timestamp 1680363874
transform 1 0 4184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8947
timestamp 1680363874
transform 1 0 4192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8951
timestamp 1680363874
transform 1 0 4200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8952
timestamp 1680363874
transform 1 0 4208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8953
timestamp 1680363874
transform 1 0 4216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8954
timestamp 1680363874
transform 1 0 4224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8955
timestamp 1680363874
transform 1 0 4232 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_300
timestamp 1680363874
transform -1 0 4280 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8956
timestamp 1680363874
transform 1 0 4280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8957
timestamp 1680363874
transform 1 0 4288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8958
timestamp 1680363874
transform 1 0 4296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8959
timestamp 1680363874
transform 1 0 4304 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7011
timestamp 1680363874
transform 1 0 4340 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_532
timestamp 1680363874
transform 1 0 4312 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8960
timestamp 1680363874
transform 1 0 4328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8961
timestamp 1680363874
transform 1 0 4336 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_464
timestamp 1680363874
transform 1 0 4344 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8962
timestamp 1680363874
transform 1 0 4440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8963
timestamp 1680363874
transform 1 0 4448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8964
timestamp 1680363874
transform 1 0 4456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8965
timestamp 1680363874
transform 1 0 4464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8966
timestamp 1680363874
transform 1 0 4472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8967
timestamp 1680363874
transform 1 0 4480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8968
timestamp 1680363874
transform 1 0 4488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8969
timestamp 1680363874
transform 1 0 4496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8970
timestamp 1680363874
transform 1 0 4504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8971
timestamp 1680363874
transform 1 0 4512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8972
timestamp 1680363874
transform 1 0 4520 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_533
timestamp 1680363874
transform 1 0 4528 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8975
timestamp 1680363874
transform 1 0 4544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8976
timestamp 1680363874
transform 1 0 4552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8977
timestamp 1680363874
transform 1 0 4560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8978
timestamp 1680363874
transform 1 0 4568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8979
timestamp 1680363874
transform 1 0 4576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8980
timestamp 1680363874
transform 1 0 4584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8981
timestamp 1680363874
transform 1 0 4592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8982
timestamp 1680363874
transform 1 0 4600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8983
timestamp 1680363874
transform 1 0 4608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8984
timestamp 1680363874
transform 1 0 4616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8985
timestamp 1680363874
transform 1 0 4624 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_301
timestamp 1680363874
transform 1 0 4632 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8986
timestamp 1680363874
transform 1 0 4672 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_535
timestamp 1680363874
transform 1 0 4680 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_467
timestamp 1680363874
transform -1 0 4792 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8988
timestamp 1680363874
transform 1 0 4792 0 -1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_73
timestamp 1680363874
transform 1 0 4851 0 1 1070
box -10 -3 10 3
use M2_M1  M2_M1_7724
timestamp 1680363874
transform 1 0 116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7831
timestamp 1680363874
transform 1 0 92 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7712
timestamp 1680363874
transform 1 0 196 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7725
timestamp 1680363874
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7726
timestamp 1680363874
transform 1 0 196 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7094
timestamp 1680363874
transform 1 0 220 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7832
timestamp 1680363874
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7915
timestamp 1680363874
transform 1 0 220 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7713
timestamp 1680363874
transform 1 0 244 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7059
timestamp 1680363874
transform 1 0 252 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7727
timestamp 1680363874
transform 1 0 236 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7095
timestamp 1680363874
transform 1 0 244 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7833
timestamp 1680363874
transform 1 0 244 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7046
timestamp 1680363874
transform 1 0 276 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7714
timestamp 1680363874
transform 1 0 276 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7728
timestamp 1680363874
transform 1 0 268 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7142
timestamp 1680363874
transform 1 0 268 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7729
timestamp 1680363874
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7047
timestamp 1680363874
transform 1 0 308 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7060
timestamp 1680363874
transform 1 0 332 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7730
timestamp 1680363874
transform 1 0 332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7731
timestamp 1680363874
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7834
timestamp 1680363874
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7835
timestamp 1680363874
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7143
timestamp 1680363874
transform 1 0 292 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7715
timestamp 1680363874
transform 1 0 404 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7061
timestamp 1680363874
transform 1 0 444 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7732
timestamp 1680363874
transform 1 0 452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7836
timestamp 1680363874
transform 1 0 444 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7124
timestamp 1680363874
transform 1 0 452 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7062
timestamp 1680363874
transform 1 0 556 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7096
timestamp 1680363874
transform 1 0 476 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7733
timestamp 1680363874
transform 1 0 500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7734
timestamp 1680363874
transform 1 0 556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7837
timestamp 1680363874
transform 1 0 476 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7125
timestamp 1680363874
transform 1 0 564 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7097
timestamp 1680363874
transform 1 0 580 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7063
timestamp 1680363874
transform 1 0 668 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7735
timestamp 1680363874
transform 1 0 604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7736
timestamp 1680363874
transform 1 0 660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7838
timestamp 1680363874
transform 1 0 580 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7048
timestamp 1680363874
transform 1 0 716 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7064
timestamp 1680363874
transform 1 0 764 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7098
timestamp 1680363874
transform 1 0 684 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7737
timestamp 1680363874
transform 1 0 708 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7099
timestamp 1680363874
transform 1 0 732 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7738
timestamp 1680363874
transform 1 0 764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7839
timestamp 1680363874
transform 1 0 684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7840
timestamp 1680363874
transform 1 0 772 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7841
timestamp 1680363874
transform 1 0 788 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7065
timestamp 1680363874
transform 1 0 828 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7739
timestamp 1680363874
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7740
timestamp 1680363874
transform 1 0 820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7842
timestamp 1680363874
transform 1 0 812 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7126
timestamp 1680363874
transform 1 0 820 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7843
timestamp 1680363874
transform 1 0 828 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7844
timestamp 1680363874
transform 1 0 836 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7049
timestamp 1680363874
transform 1 0 948 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7066
timestamp 1680363874
transform 1 0 860 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7067
timestamp 1680363874
transform 1 0 924 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7741
timestamp 1680363874
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7127
timestamp 1680363874
transform 1 0 844 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7845
timestamp 1680363874
transform 1 0 852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7742
timestamp 1680363874
transform 1 0 860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7743
timestamp 1680363874
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7744
timestamp 1680363874
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7846
timestamp 1680363874
transform 1 0 948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7847
timestamp 1680363874
transform 1 0 964 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7144
timestamp 1680363874
transform 1 0 964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7169
timestamp 1680363874
transform 1 0 932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7170
timestamp 1680363874
transform 1 0 972 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7745
timestamp 1680363874
transform 1 0 996 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7128
timestamp 1680363874
transform 1 0 996 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7746
timestamp 1680363874
transform 1 0 1068 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7848
timestamp 1680363874
transform 1 0 1020 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7145
timestamp 1680363874
transform 1 0 1020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7146
timestamp 1680363874
transform 1 0 1068 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7171
timestamp 1680363874
transform 1 0 1012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7172
timestamp 1680363874
transform 1 0 1052 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7849
timestamp 1680363874
transform 1 0 1132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7068
timestamp 1680363874
transform 1 0 1188 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7747
timestamp 1680363874
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7100
timestamp 1680363874
transform 1 0 1164 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7748
timestamp 1680363874
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7749
timestamp 1680363874
transform 1 0 1188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7850
timestamp 1680363874
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7129
timestamp 1680363874
transform 1 0 1188 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7851
timestamp 1680363874
transform 1 0 1196 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7147
timestamp 1680363874
transform 1 0 1180 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7173
timestamp 1680363874
transform 1 0 1164 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7750
timestamp 1680363874
transform 1 0 1212 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7174
timestamp 1680363874
transform 1 0 1204 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7101
timestamp 1680363874
transform 1 0 1220 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7852
timestamp 1680363874
transform 1 0 1236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7751
timestamp 1680363874
transform 1 0 1268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7752
timestamp 1680363874
transform 1 0 1284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7853
timestamp 1680363874
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7854
timestamp 1680363874
transform 1 0 1276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7855
timestamp 1680363874
transform 1 0 1300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7148
timestamp 1680363874
transform 1 0 1308 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7856
timestamp 1680363874
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7149
timestamp 1680363874
transform 1 0 1324 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7753
timestamp 1680363874
transform 1 0 1420 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7130
timestamp 1680363874
transform 1 0 1420 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7857
timestamp 1680363874
transform 1 0 1428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7858
timestamp 1680363874
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7131
timestamp 1680363874
transform 1 0 1452 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7069
timestamp 1680363874
transform 1 0 1492 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7754
timestamp 1680363874
transform 1 0 1460 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7102
timestamp 1680363874
transform 1 0 1468 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7755
timestamp 1680363874
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7756
timestamp 1680363874
transform 1 0 1492 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7103
timestamp 1680363874
transform 1 0 1508 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7859
timestamp 1680363874
transform 1 0 1484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7860
timestamp 1680363874
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7861
timestamp 1680363874
transform 1 0 1508 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7150
timestamp 1680363874
transform 1 0 1484 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7151
timestamp 1680363874
transform 1 0 1516 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7033
timestamp 1680363874
transform 1 0 1548 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7070
timestamp 1680363874
transform 1 0 1564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7757
timestamp 1680363874
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7758
timestamp 1680363874
transform 1 0 1564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7759
timestamp 1680363874
transform 1 0 1580 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7132
timestamp 1680363874
transform 1 0 1564 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7862
timestamp 1680363874
transform 1 0 1572 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7050
timestamp 1680363874
transform 1 0 1604 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7716
timestamp 1680363874
transform 1 0 1604 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7104
timestamp 1680363874
transform 1 0 1596 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7012
timestamp 1680363874
transform 1 0 1644 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7034
timestamp 1680363874
transform 1 0 1636 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7709
timestamp 1680363874
transform 1 0 1644 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_7071
timestamp 1680363874
transform 1 0 1636 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7035
timestamp 1680363874
transform 1 0 1660 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7717
timestamp 1680363874
transform 1 0 1652 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7105
timestamp 1680363874
transform 1 0 1628 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7760
timestamp 1680363874
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7152
timestamp 1680363874
transform 1 0 1620 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7020
timestamp 1680363874
transform 1 0 1748 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7021
timestamp 1680363874
transform 1 0 1780 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7036
timestamp 1680363874
transform 1 0 1700 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7037
timestamp 1680363874
transform 1 0 1748 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7072
timestamp 1680363874
transform 1 0 1692 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7106
timestamp 1680363874
transform 1 0 1708 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7107
timestamp 1680363874
transform 1 0 1732 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7761
timestamp 1680363874
transform 1 0 1756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7863
timestamp 1680363874
transform 1 0 1708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7153
timestamp 1680363874
transform 1 0 1708 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7175
timestamp 1680363874
transform 1 0 1748 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7176
timestamp 1680363874
transform 1 0 1780 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7718
timestamp 1680363874
transform 1 0 1796 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7762
timestamp 1680363874
transform 1 0 1804 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7154
timestamp 1680363874
transform 1 0 1804 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7038
timestamp 1680363874
transform 1 0 1836 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7051
timestamp 1680363874
transform 1 0 1836 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7710
timestamp 1680363874
transform 1 0 1844 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_7719
timestamp 1680363874
transform 1 0 1852 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7763
timestamp 1680363874
transform 1 0 1836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7764
timestamp 1680363874
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7765
timestamp 1680363874
transform 1 0 1916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7766
timestamp 1680363874
transform 1 0 1932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7864
timestamp 1680363874
transform 1 0 1892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7865
timestamp 1680363874
transform 1 0 1908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7866
timestamp 1680363874
transform 1 0 1924 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7155
timestamp 1680363874
transform 1 0 1924 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7867
timestamp 1680363874
transform 1 0 1972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7767
timestamp 1680363874
transform 1 0 1988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7868
timestamp 1680363874
transform 1 0 2004 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7073
timestamp 1680363874
transform 1 0 2036 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7768
timestamp 1680363874
transform 1 0 2020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7769
timestamp 1680363874
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7869
timestamp 1680363874
transform 1 0 2028 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7133
timestamp 1680363874
transform 1 0 2036 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7870
timestamp 1680363874
transform 1 0 2052 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7156
timestamp 1680363874
transform 1 0 2044 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7720
timestamp 1680363874
transform 1 0 2068 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7013
timestamp 1680363874
transform 1 0 2116 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7039
timestamp 1680363874
transform 1 0 2108 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7711
timestamp 1680363874
transform 1 0 2108 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_7770
timestamp 1680363874
transform 1 0 2100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7721
timestamp 1680363874
transform 1 0 2124 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7771
timestamp 1680363874
transform 1 0 2124 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7134
timestamp 1680363874
transform 1 0 2124 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7772
timestamp 1680363874
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7108
timestamp 1680363874
transform 1 0 2188 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7871
timestamp 1680363874
transform 1 0 2180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7177
timestamp 1680363874
transform 1 0 2188 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7135
timestamp 1680363874
transform 1 0 2244 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7722
timestamp 1680363874
transform 1 0 2260 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7872
timestamp 1680363874
transform 1 0 2268 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7052
timestamp 1680363874
transform 1 0 2284 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7773
timestamp 1680363874
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7136
timestamp 1680363874
transform 1 0 2300 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7774
timestamp 1680363874
transform 1 0 2324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7873
timestamp 1680363874
transform 1 0 2340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7775
timestamp 1680363874
transform 1 0 2356 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7178
timestamp 1680363874
transform 1 0 2348 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7022
timestamp 1680363874
transform 1 0 2396 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7776
timestamp 1680363874
transform 1 0 2420 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7023
timestamp 1680363874
transform 1 0 2460 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7040
timestamp 1680363874
transform 1 0 2436 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7074
timestamp 1680363874
transform 1 0 2444 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7777
timestamp 1680363874
transform 1 0 2444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7778
timestamp 1680363874
transform 1 0 2460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7779
timestamp 1680363874
transform 1 0 2468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7874
timestamp 1680363874
transform 1 0 2452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7875
timestamp 1680363874
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7075
timestamp 1680363874
transform 1 0 2492 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7876
timestamp 1680363874
transform 1 0 2492 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7137
timestamp 1680363874
transform 1 0 2516 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7780
timestamp 1680363874
transform 1 0 2532 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7024
timestamp 1680363874
transform 1 0 2588 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7025
timestamp 1680363874
transform 1 0 2644 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7041
timestamp 1680363874
transform 1 0 2660 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7076
timestamp 1680363874
transform 1 0 2620 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7077
timestamp 1680363874
transform 1 0 2660 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7781
timestamp 1680363874
transform 1 0 2620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7782
timestamp 1680363874
transform 1 0 2660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7877
timestamp 1680363874
transform 1 0 2644 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7179
timestamp 1680363874
transform 1 0 2652 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7042
timestamp 1680363874
transform 1 0 2692 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7878
timestamp 1680363874
transform 1 0 2708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7180
timestamp 1680363874
transform 1 0 2700 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7181
timestamp 1680363874
transform 1 0 2724 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7043
timestamp 1680363874
transform 1 0 2812 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7078
timestamp 1680363874
transform 1 0 2804 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7783
timestamp 1680363874
transform 1 0 2796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7784
timestamp 1680363874
transform 1 0 2804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7785
timestamp 1680363874
transform 1 0 2820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7879
timestamp 1680363874
transform 1 0 2804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7880
timestamp 1680363874
transform 1 0 2812 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7079
timestamp 1680363874
transform 1 0 2844 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7080
timestamp 1680363874
transform 1 0 2860 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7786
timestamp 1680363874
transform 1 0 2860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7881
timestamp 1680363874
transform 1 0 2860 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7014
timestamp 1680363874
transform 1 0 2876 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7787
timestamp 1680363874
transform 1 0 2876 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7109
timestamp 1680363874
transform 1 0 2884 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7882
timestamp 1680363874
transform 1 0 2884 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7157
timestamp 1680363874
transform 1 0 2892 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7026
timestamp 1680363874
transform 1 0 2924 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7723
timestamp 1680363874
transform 1 0 2924 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7788
timestamp 1680363874
transform 1 0 2916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7883
timestamp 1680363874
transform 1 0 2908 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7044
timestamp 1680363874
transform 1 0 2956 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7138
timestamp 1680363874
transform 1 0 2948 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7045
timestamp 1680363874
transform 1 0 2972 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7081
timestamp 1680363874
transform 1 0 2996 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7789
timestamp 1680363874
transform 1 0 2964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7790
timestamp 1680363874
transform 1 0 2980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7791
timestamp 1680363874
transform 1 0 2996 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7884
timestamp 1680363874
transform 1 0 2964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7885
timestamp 1680363874
transform 1 0 2972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7886
timestamp 1680363874
transform 1 0 2988 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7015
timestamp 1680363874
transform 1 0 3012 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7707
timestamp 1680363874
transform 1 0 3012 0 1 1055
box -2 -2 2 2
use M3_M2  M3_M2_7027
timestamp 1680363874
transform 1 0 3028 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7708
timestamp 1680363874
transform 1 0 3036 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_7916
timestamp 1680363874
transform 1 0 3044 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7887
timestamp 1680363874
transform 1 0 3068 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7110
timestamp 1680363874
transform 1 0 3108 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7917
timestamp 1680363874
transform 1 0 3108 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7918
timestamp 1680363874
transform 1 0 3116 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7792
timestamp 1680363874
transform 1 0 3156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7793
timestamp 1680363874
transform 1 0 3172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7794
timestamp 1680363874
transform 1 0 3188 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7182
timestamp 1680363874
transform 1 0 3188 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7795
timestamp 1680363874
transform 1 0 3244 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7111
timestamp 1680363874
transform 1 0 3252 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7888
timestamp 1680363874
transform 1 0 3228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7889
timestamp 1680363874
transform 1 0 3236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7890
timestamp 1680363874
transform 1 0 3252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7891
timestamp 1680363874
transform 1 0 3260 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7158
timestamp 1680363874
transform 1 0 3236 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7796
timestamp 1680363874
transform 1 0 3276 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7139
timestamp 1680363874
transform 1 0 3276 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7053
timestamp 1680363874
transform 1 0 3308 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7082
timestamp 1680363874
transform 1 0 3308 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7797
timestamp 1680363874
transform 1 0 3308 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7054
timestamp 1680363874
transform 1 0 3364 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7083
timestamp 1680363874
transform 1 0 3356 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7798
timestamp 1680363874
transform 1 0 3324 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7112
timestamp 1680363874
transform 1 0 3332 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7799
timestamp 1680363874
transform 1 0 3356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7892
timestamp 1680363874
transform 1 0 3404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7084
timestamp 1680363874
transform 1 0 3428 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7055
timestamp 1680363874
transform 1 0 3556 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7085
timestamp 1680363874
transform 1 0 3460 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7086
timestamp 1680363874
transform 1 0 3524 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7087
timestamp 1680363874
transform 1 0 3564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7800
timestamp 1680363874
transform 1 0 3428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7801
timestamp 1680363874
transform 1 0 3452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7802
timestamp 1680363874
transform 1 0 3468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7803
timestamp 1680363874
transform 1 0 3524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7893
timestamp 1680363874
transform 1 0 3420 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7113
timestamp 1680363874
transform 1 0 3548 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7804
timestamp 1680363874
transform 1 0 3564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7894
timestamp 1680363874
transform 1 0 3444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7895
timestamp 1680363874
transform 1 0 3460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7896
timestamp 1680363874
transform 1 0 3548 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7159
timestamp 1680363874
transform 1 0 3460 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7183
timestamp 1680363874
transform 1 0 3436 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7184
timestamp 1680363874
transform 1 0 3548 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7028
timestamp 1680363874
transform 1 0 3588 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7056
timestamp 1680363874
transform 1 0 3580 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7805
timestamp 1680363874
transform 1 0 3588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7897
timestamp 1680363874
transform 1 0 3588 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7029
timestamp 1680363874
transform 1 0 3604 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7016
timestamp 1680363874
transform 1 0 3644 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7806
timestamp 1680363874
transform 1 0 3612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7807
timestamp 1680363874
transform 1 0 3628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7808
timestamp 1680363874
transform 1 0 3636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7898
timestamp 1680363874
transform 1 0 3604 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7160
timestamp 1680363874
transform 1 0 3636 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7899
timestamp 1680363874
transform 1 0 3652 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7017
timestamp 1680363874
transform 1 0 3692 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7030
timestamp 1680363874
transform 1 0 3676 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7809
timestamp 1680363874
transform 1 0 3724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7900
timestamp 1680363874
transform 1 0 3748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7810
timestamp 1680363874
transform 1 0 3764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7811
timestamp 1680363874
transform 1 0 3836 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7114
timestamp 1680363874
transform 1 0 3884 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7812
timestamp 1680363874
transform 1 0 3900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7813
timestamp 1680363874
transform 1 0 3956 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7901
timestamp 1680363874
transform 1 0 3884 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7161
timestamp 1680363874
transform 1 0 3844 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7162
timestamp 1680363874
transform 1 0 3868 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7115
timestamp 1680363874
transform 1 0 3980 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7902
timestamp 1680363874
transform 1 0 3980 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7031
timestamp 1680363874
transform 1 0 4100 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7088
timestamp 1680363874
transform 1 0 4060 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7089
timestamp 1680363874
transform 1 0 4100 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7116
timestamp 1680363874
transform 1 0 4012 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7814
timestamp 1680363874
transform 1 0 4060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7815
timestamp 1680363874
transform 1 0 4092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7816
timestamp 1680363874
transform 1 0 4100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7903
timestamp 1680363874
transform 1 0 4012 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7904
timestamp 1680363874
transform 1 0 4100 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7163
timestamp 1680363874
transform 1 0 4012 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7185
timestamp 1680363874
transform 1 0 4012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7186
timestamp 1680363874
transform 1 0 4036 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7817
timestamp 1680363874
transform 1 0 4116 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7117
timestamp 1680363874
transform 1 0 4132 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7032
timestamp 1680363874
transform 1 0 4196 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7090
timestamp 1680363874
transform 1 0 4196 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7118
timestamp 1680363874
transform 1 0 4172 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7818
timestamp 1680363874
transform 1 0 4180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7819
timestamp 1680363874
transform 1 0 4196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7820
timestamp 1680363874
transform 1 0 4204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7905
timestamp 1680363874
transform 1 0 4172 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7187
timestamp 1680363874
transform 1 0 4172 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7821
timestamp 1680363874
transform 1 0 4284 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7119
timestamp 1680363874
transform 1 0 4308 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7906
timestamp 1680363874
transform 1 0 4308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7188
timestamp 1680363874
transform 1 0 4276 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7018
timestamp 1680363874
transform 1 0 4340 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7120
timestamp 1680363874
transform 1 0 4356 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7164
timestamp 1680363874
transform 1 0 4372 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7019
timestamp 1680363874
transform 1 0 4396 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7822
timestamp 1680363874
transform 1 0 4388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7823
timestamp 1680363874
transform 1 0 4460 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7091
timestamp 1680363874
transform 1 0 4476 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7092
timestamp 1680363874
transform 1 0 4500 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7121
timestamp 1680363874
transform 1 0 4476 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7824
timestamp 1680363874
transform 1 0 4484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7825
timestamp 1680363874
transform 1 0 4500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7907
timestamp 1680363874
transform 1 0 4468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7908
timestamp 1680363874
transform 1 0 4476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7909
timestamp 1680363874
transform 1 0 4492 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7165
timestamp 1680363874
transform 1 0 4468 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7166
timestamp 1680363874
transform 1 0 4484 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7826
timestamp 1680363874
transform 1 0 4548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7827
timestamp 1680363874
transform 1 0 4588 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7140
timestamp 1680363874
transform 1 0 4564 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7910
timestamp 1680363874
transform 1 0 4580 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7141
timestamp 1680363874
transform 1 0 4588 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7057
timestamp 1680363874
transform 1 0 4604 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7093
timestamp 1680363874
transform 1 0 4612 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7828
timestamp 1680363874
transform 1 0 4612 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7189
timestamp 1680363874
transform 1 0 4612 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7058
timestamp 1680363874
transform 1 0 4636 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7829
timestamp 1680363874
transform 1 0 4652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7830
timestamp 1680363874
transform 1 0 4668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7911
timestamp 1680363874
transform 1 0 4636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7912
timestamp 1680363874
transform 1 0 4644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7913
timestamp 1680363874
transform 1 0 4660 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7167
timestamp 1680363874
transform 1 0 4636 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7168
timestamp 1680363874
transform 1 0 4660 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7190
timestamp 1680363874
transform 1 0 4644 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7122
timestamp 1680363874
transform 1 0 4676 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7914
timestamp 1680363874
transform 1 0 4700 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7123
timestamp 1680363874
transform 1 0 4748 0 1 1015
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_74
timestamp 1680363874
transform 1 0 48 0 1 970
box -10 -3 10 3
use FILL  FILL_8989
timestamp 1680363874
transform 1 0 72 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_468
timestamp 1680363874
transform 1 0 80 0 1 970
box -8 -3 104 105
use FILL  FILL_8990
timestamp 1680363874
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_8993
timestamp 1680363874
transform 1 0 184 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_54
timestamp 1680363874
transform -1 0 216 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1680363874
transform 1 0 216 0 1 970
box -8 -3 32 105
use FILL  FILL_8995
timestamp 1680363874
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_8996
timestamp 1680363874
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_8997
timestamp 1680363874
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_8998
timestamp 1680363874
transform 1 0 264 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_55
timestamp 1680363874
transform -1 0 296 0 1 970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_470
timestamp 1680363874
transform 1 0 296 0 1 970
box -8 -3 104 105
use FILL  FILL_8999
timestamp 1680363874
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_9000
timestamp 1680363874
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_9001
timestamp 1680363874
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_9002
timestamp 1680363874
transform 1 0 416 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_56
timestamp 1680363874
transform -1 0 448 0 1 970
box -8 -3 32 105
use FILL  FILL_9003
timestamp 1680363874
transform 1 0 448 0 1 970
box -8 -3 16 105
use FILL  FILL_9004
timestamp 1680363874
transform 1 0 456 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_471
timestamp 1680363874
transform 1 0 464 0 1 970
box -8 -3 104 105
use FILL  FILL_9005
timestamp 1680363874
transform 1 0 560 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_472
timestamp 1680363874
transform 1 0 568 0 1 970
box -8 -3 104 105
use FILL  FILL_9006
timestamp 1680363874
transform 1 0 664 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_473
timestamp 1680363874
transform 1 0 672 0 1 970
box -8 -3 104 105
use FILL  FILL_9007
timestamp 1680363874
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_9008
timestamp 1680363874
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_9009
timestamp 1680363874
transform 1 0 784 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_340
timestamp 1680363874
transform 1 0 792 0 1 970
box -8 -3 46 105
use INVX2  INVX2_536
timestamp 1680363874
transform 1 0 832 0 1 970
box -9 -3 26 105
use INVX2  INVX2_537
timestamp 1680363874
transform 1 0 848 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_474
timestamp 1680363874
transform -1 0 960 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7191
timestamp 1680363874
transform 1 0 972 0 1 975
box -3 -3 3 3
use INVX2  INVX2_538
timestamp 1680363874
transform 1 0 960 0 1 970
box -9 -3 26 105
use FILL  FILL_9010
timestamp 1680363874
transform 1 0 976 0 1 970
box -8 -3 16 105
use FILL  FILL_9011
timestamp 1680363874
transform 1 0 984 0 1 970
box -8 -3 16 105
use FILL  FILL_9012
timestamp 1680363874
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_9013
timestamp 1680363874
transform 1 0 1000 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_475
timestamp 1680363874
transform 1 0 1008 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7192
timestamp 1680363874
transform 1 0 1116 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7193
timestamp 1680363874
transform 1 0 1132 0 1 975
box -3 -3 3 3
use INVX2  INVX2_539
timestamp 1680363874
transform 1 0 1104 0 1 970
box -9 -3 26 105
use FILL  FILL_9014
timestamp 1680363874
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_9015
timestamp 1680363874
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_9016
timestamp 1680363874
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_9017
timestamp 1680363874
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_9018
timestamp 1680363874
transform 1 0 1152 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_341
timestamp 1680363874
transform -1 0 1200 0 1 970
box -8 -3 46 105
use FILL  FILL_9019
timestamp 1680363874
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_9020
timestamp 1680363874
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_9021
timestamp 1680363874
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_9022
timestamp 1680363874
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_9023
timestamp 1680363874
transform 1 0 1232 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_342
timestamp 1680363874
transform 1 0 1240 0 1 970
box -8 -3 46 105
use FILL  FILL_9024
timestamp 1680363874
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_9046
timestamp 1680363874
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_9048
timestamp 1680363874
transform 1 0 1296 0 1 970
box -8 -3 16 105
use INVX2  INVX2_544
timestamp 1680363874
transform 1 0 1304 0 1 970
box -9 -3 26 105
use FILL  FILL_9050
timestamp 1680363874
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_9051
timestamp 1680363874
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_9052
timestamp 1680363874
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_9053
timestamp 1680363874
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_9054
timestamp 1680363874
transform 1 0 1352 0 1 970
box -8 -3 16 105
use INVX2  INVX2_545
timestamp 1680363874
transform 1 0 1360 0 1 970
box -9 -3 26 105
use FILL  FILL_9055
timestamp 1680363874
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_9056
timestamp 1680363874
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_9057
timestamp 1680363874
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_9058
timestamp 1680363874
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_9059
timestamp 1680363874
transform 1 0 1408 0 1 970
box -8 -3 16 105
use FILL  FILL_9062
timestamp 1680363874
transform 1 0 1416 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7194
timestamp 1680363874
transform 1 0 1444 0 1 975
box -3 -3 3 3
use INVX2  INVX2_546
timestamp 1680363874
transform 1 0 1424 0 1 970
box -9 -3 26 105
use FILL  FILL_9064
timestamp 1680363874
transform 1 0 1440 0 1 970
box -8 -3 16 105
use FILL  FILL_9065
timestamp 1680363874
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_9066
timestamp 1680363874
transform 1 0 1456 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_346
timestamp 1680363874
transform -1 0 1504 0 1 970
box -8 -3 46 105
use FILL  FILL_9067
timestamp 1680363874
transform 1 0 1504 0 1 970
box -8 -3 16 105
use FILL  FILL_9068
timestamp 1680363874
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_9069
timestamp 1680363874
transform 1 0 1520 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7195
timestamp 1680363874
transform 1 0 1540 0 1 975
box -3 -3 3 3
use FILL  FILL_9070
timestamp 1680363874
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_9071
timestamp 1680363874
transform 1 0 1536 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_302
timestamp 1680363874
transform -1 0 1584 0 1 970
box -8 -3 46 105
use FILL  FILL_9072
timestamp 1680363874
transform 1 0 1584 0 1 970
box -8 -3 16 105
use FILL  FILL_9073
timestamp 1680363874
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_9074
timestamp 1680363874
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_9081
timestamp 1680363874
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_9082
timestamp 1680363874
transform 1 0 1616 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_65
timestamp 1680363874
transform 1 0 1624 0 1 970
box -8 -3 40 105
use FILL  FILL_9083
timestamp 1680363874
transform 1 0 1656 0 1 970
box -8 -3 16 105
use FILL  FILL_9086
timestamp 1680363874
transform 1 0 1664 0 1 970
box -8 -3 16 105
use FILL  FILL_9088
timestamp 1680363874
transform 1 0 1672 0 1 970
box -8 -3 16 105
use FILL  FILL_9090
timestamp 1680363874
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_9092
timestamp 1680363874
transform 1 0 1688 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7196
timestamp 1680363874
transform 1 0 1716 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7197
timestamp 1680363874
transform 1 0 1740 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_485
timestamp 1680363874
transform 1 0 1696 0 1 970
box -8 -3 104 105
use FILL  FILL_9093
timestamp 1680363874
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_9101
timestamp 1680363874
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_9102
timestamp 1680363874
transform 1 0 1808 0 1 970
box -8 -3 16 105
use FILL  FILL_9103
timestamp 1680363874
transform 1 0 1816 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_66
timestamp 1680363874
transform 1 0 1824 0 1 970
box -8 -3 40 105
use FILL  FILL_9104
timestamp 1680363874
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_9105
timestamp 1680363874
transform 1 0 1864 0 1 970
box -8 -3 16 105
use FILL  FILL_9106
timestamp 1680363874
transform 1 0 1872 0 1 970
box -8 -3 16 105
use FILL  FILL_9112
timestamp 1680363874
transform 1 0 1880 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_350
timestamp 1680363874
transform 1 0 1888 0 1 970
box -8 -3 46 105
use FILL  FILL_9113
timestamp 1680363874
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_9114
timestamp 1680363874
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_9115
timestamp 1680363874
transform 1 0 1944 0 1 970
box -8 -3 16 105
use INVX2  INVX2_549
timestamp 1680363874
transform -1 0 1968 0 1 970
box -9 -3 26 105
use FILL  FILL_9116
timestamp 1680363874
transform 1 0 1968 0 1 970
box -8 -3 16 105
use FILL  FILL_9117
timestamp 1680363874
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_9119
timestamp 1680363874
transform 1 0 1984 0 1 970
box -8 -3 16 105
use FILL  FILL_9121
timestamp 1680363874
transform 1 0 1992 0 1 970
box -8 -3 16 105
use FILL  FILL_9123
timestamp 1680363874
transform 1 0 2000 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_351
timestamp 1680363874
transform -1 0 2048 0 1 970
box -8 -3 46 105
use FILL  FILL_9124
timestamp 1680363874
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_9127
timestamp 1680363874
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_9129
timestamp 1680363874
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_9131
timestamp 1680363874
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_9133
timestamp 1680363874
transform 1 0 2080 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_67
timestamp 1680363874
transform 1 0 2088 0 1 970
box -8 -3 40 105
use FILL  FILL_9135
timestamp 1680363874
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_9136
timestamp 1680363874
transform 1 0 2128 0 1 970
box -8 -3 16 105
use FILL  FILL_9137
timestamp 1680363874
transform 1 0 2136 0 1 970
box -8 -3 16 105
use INVX2  INVX2_550
timestamp 1680363874
transform -1 0 2160 0 1 970
box -9 -3 26 105
use FILL  FILL_9138
timestamp 1680363874
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_9139
timestamp 1680363874
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_9140
timestamp 1680363874
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_9141
timestamp 1680363874
transform 1 0 2184 0 1 970
box -8 -3 16 105
use FILL  FILL_9143
timestamp 1680363874
transform 1 0 2192 0 1 970
box -8 -3 16 105
use FILL  FILL_9144
timestamp 1680363874
transform 1 0 2200 0 1 970
box -8 -3 16 105
use FILL  FILL_9145
timestamp 1680363874
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_9146
timestamp 1680363874
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_9147
timestamp 1680363874
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_9148
timestamp 1680363874
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_9151
timestamp 1680363874
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_9153
timestamp 1680363874
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_9155
timestamp 1680363874
transform 1 0 2256 0 1 970
box -8 -3 16 105
use FILL  FILL_9157
timestamp 1680363874
transform 1 0 2264 0 1 970
box -8 -3 16 105
use FILL  FILL_9158
timestamp 1680363874
transform 1 0 2272 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_157
timestamp 1680363874
transform -1 0 2312 0 1 970
box -8 -3 34 105
use FILL  FILL_9159
timestamp 1680363874
transform 1 0 2312 0 1 970
box -8 -3 16 105
use FILL  FILL_9160
timestamp 1680363874
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_9161
timestamp 1680363874
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_9162
timestamp 1680363874
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_9163
timestamp 1680363874
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_9164
timestamp 1680363874
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_9165
timestamp 1680363874
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_9166
timestamp 1680363874
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_9167
timestamp 1680363874
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_9168
timestamp 1680363874
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_9169
timestamp 1680363874
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_9170
timestamp 1680363874
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_9173
timestamp 1680363874
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_9175
timestamp 1680363874
transform 1 0 2416 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_303
timestamp 1680363874
transform -1 0 2464 0 1 970
box -8 -3 46 105
use FILL  FILL_9177
timestamp 1680363874
transform 1 0 2464 0 1 970
box -8 -3 16 105
use FILL  FILL_9179
timestamp 1680363874
transform 1 0 2472 0 1 970
box -8 -3 16 105
use INVX2  INVX2_553
timestamp 1680363874
transform -1 0 2496 0 1 970
box -9 -3 26 105
use FILL  FILL_9180
timestamp 1680363874
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_9181
timestamp 1680363874
transform 1 0 2504 0 1 970
box -8 -3 16 105
use FILL  FILL_9182
timestamp 1680363874
transform 1 0 2512 0 1 970
box -8 -3 16 105
use FILL  FILL_9183
timestamp 1680363874
transform 1 0 2520 0 1 970
box -8 -3 16 105
use FILL  FILL_9184
timestamp 1680363874
transform 1 0 2528 0 1 970
box -8 -3 16 105
use FILL  FILL_9189
timestamp 1680363874
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_9190
timestamp 1680363874
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_9191
timestamp 1680363874
transform 1 0 2552 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_489
timestamp 1680363874
transform -1 0 2656 0 1 970
box -8 -3 104 105
use INVX2  INVX2_554
timestamp 1680363874
transform -1 0 2672 0 1 970
box -9 -3 26 105
use FILL  FILL_9192
timestamp 1680363874
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_9201
timestamp 1680363874
transform 1 0 2680 0 1 970
box -8 -3 16 105
use FILL  FILL_9202
timestamp 1680363874
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_9203
timestamp 1680363874
transform 1 0 2696 0 1 970
box -8 -3 16 105
use FILL  FILL_9204
timestamp 1680363874
transform 1 0 2704 0 1 970
box -8 -3 16 105
use FILL  FILL_9205
timestamp 1680363874
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_9206
timestamp 1680363874
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_9207
timestamp 1680363874
transform 1 0 2728 0 1 970
box -8 -3 16 105
use FILL  FILL_9210
timestamp 1680363874
transform 1 0 2736 0 1 970
box -8 -3 16 105
use INVX2  INVX2_556
timestamp 1680363874
transform -1 0 2760 0 1 970
box -9 -3 26 105
use FILL  FILL_9211
timestamp 1680363874
transform 1 0 2760 0 1 970
box -8 -3 16 105
use FILL  FILL_9212
timestamp 1680363874
transform 1 0 2768 0 1 970
box -8 -3 16 105
use FILL  FILL_9213
timestamp 1680363874
transform 1 0 2776 0 1 970
box -8 -3 16 105
use FILL  FILL_9214
timestamp 1680363874
transform 1 0 2784 0 1 970
box -8 -3 16 105
use FILL  FILL_9215
timestamp 1680363874
transform 1 0 2792 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_307
timestamp 1680363874
transform 1 0 2800 0 1 970
box -8 -3 46 105
use FILL  FILL_9216
timestamp 1680363874
transform 1 0 2840 0 1 970
box -8 -3 16 105
use FILL  FILL_9217
timestamp 1680363874
transform 1 0 2848 0 1 970
box -8 -3 16 105
use FILL  FILL_9218
timestamp 1680363874
transform 1 0 2856 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_353
timestamp 1680363874
transform -1 0 2904 0 1 970
box -8 -3 46 105
use FILL  FILL_9219
timestamp 1680363874
transform 1 0 2904 0 1 970
box -8 -3 16 105
use FILL  FILL_9220
timestamp 1680363874
transform 1 0 2912 0 1 970
box -8 -3 16 105
use FILL  FILL_9221
timestamp 1680363874
transform 1 0 2920 0 1 970
box -8 -3 16 105
use FILL  FILL_9222
timestamp 1680363874
transform 1 0 2928 0 1 970
box -8 -3 16 105
use INVX2  INVX2_557
timestamp 1680363874
transform -1 0 2952 0 1 970
box -9 -3 26 105
use FILL  FILL_9223
timestamp 1680363874
transform 1 0 2952 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_308
timestamp 1680363874
transform 1 0 2960 0 1 970
box -8 -3 46 105
use FILL  FILL_9224
timestamp 1680363874
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_9233
timestamp 1680363874
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_9235
timestamp 1680363874
transform 1 0 3016 0 1 970
box -8 -3 16 105
use FILL  FILL_9237
timestamp 1680363874
transform 1 0 3024 0 1 970
box -8 -3 16 105
use FILL  FILL_9238
timestamp 1680363874
transform 1 0 3032 0 1 970
box -8 -3 16 105
use FILL  FILL_9239
timestamp 1680363874
transform 1 0 3040 0 1 970
box -8 -3 16 105
use FILL  FILL_9240
timestamp 1680363874
transform 1 0 3048 0 1 970
box -8 -3 16 105
use FILL  FILL_9241
timestamp 1680363874
transform 1 0 3056 0 1 970
box -8 -3 16 105
use FILL  FILL_9242
timestamp 1680363874
transform 1 0 3064 0 1 970
box -8 -3 16 105
use FILL  FILL_9243
timestamp 1680363874
transform 1 0 3072 0 1 970
box -8 -3 16 105
use FILL  FILL_9244
timestamp 1680363874
transform 1 0 3080 0 1 970
box -8 -3 16 105
use FILL  FILL_9245
timestamp 1680363874
transform 1 0 3088 0 1 970
box -8 -3 16 105
use FILL  FILL_9246
timestamp 1680363874
transform 1 0 3096 0 1 970
box -8 -3 16 105
use FILL  FILL_9247
timestamp 1680363874
transform 1 0 3104 0 1 970
box -8 -3 16 105
use FILL  FILL_9248
timestamp 1680363874
transform 1 0 3112 0 1 970
box -8 -3 16 105
use FILL  FILL_9249
timestamp 1680363874
transform 1 0 3120 0 1 970
box -8 -3 16 105
use FILL  FILL_9250
timestamp 1680363874
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_9251
timestamp 1680363874
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_9252
timestamp 1680363874
transform 1 0 3144 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7198
timestamp 1680363874
transform 1 0 3164 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7199
timestamp 1680363874
transform 1 0 3188 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_309
timestamp 1680363874
transform -1 0 3192 0 1 970
box -8 -3 46 105
use FILL  FILL_9253
timestamp 1680363874
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_9254
timestamp 1680363874
transform 1 0 3200 0 1 970
box -8 -3 16 105
use FILL  FILL_9255
timestamp 1680363874
transform 1 0 3208 0 1 970
box -8 -3 16 105
use FILL  FILL_9256
timestamp 1680363874
transform 1 0 3216 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_310
timestamp 1680363874
transform 1 0 3224 0 1 970
box -8 -3 46 105
use FILL  FILL_9257
timestamp 1680363874
transform 1 0 3264 0 1 970
box -8 -3 16 105
use FILL  FILL_9258
timestamp 1680363874
transform 1 0 3272 0 1 970
box -8 -3 16 105
use INVX2  INVX2_559
timestamp 1680363874
transform 1 0 3280 0 1 970
box -9 -3 26 105
use FILL  FILL_9259
timestamp 1680363874
transform 1 0 3296 0 1 970
box -8 -3 16 105
use FILL  FILL_9260
timestamp 1680363874
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_9266
timestamp 1680363874
transform 1 0 3312 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7200
timestamp 1680363874
transform 1 0 3404 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_494
timestamp 1680363874
transform -1 0 3416 0 1 970
box -8 -3 104 105
use FILL  FILL_9267
timestamp 1680363874
transform 1 0 3416 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7201
timestamp 1680363874
transform 1 0 3444 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_354
timestamp 1680363874
transform 1 0 3424 0 1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_495
timestamp 1680363874
transform -1 0 3560 0 1 970
box -8 -3 104 105
use INVX2  INVX2_561
timestamp 1680363874
transform -1 0 3576 0 1 970
box -9 -3 26 105
use FILL  FILL_9268
timestamp 1680363874
transform 1 0 3576 0 1 970
box -8 -3 16 105
use FILL  FILL_9269
timestamp 1680363874
transform 1 0 3584 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_312
timestamp 1680363874
transform -1 0 3632 0 1 970
box -8 -3 46 105
use FILL  FILL_9270
timestamp 1680363874
transform 1 0 3632 0 1 970
box -8 -3 16 105
use FILL  FILL_9291
timestamp 1680363874
transform 1 0 3640 0 1 970
box -8 -3 16 105
use FILL  FILL_9293
timestamp 1680363874
transform 1 0 3648 0 1 970
box -8 -3 16 105
use FILL  FILL_9294
timestamp 1680363874
transform 1 0 3656 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7202
timestamp 1680363874
transform 1 0 3716 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7203
timestamp 1680363874
transform 1 0 3740 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_497
timestamp 1680363874
transform -1 0 3760 0 1 970
box -8 -3 104 105
use FILL  FILL_9295
timestamp 1680363874
transform 1 0 3760 0 1 970
box -8 -3 16 105
use FILL  FILL_9296
timestamp 1680363874
transform 1 0 3768 0 1 970
box -8 -3 16 105
use FILL  FILL_9297
timestamp 1680363874
transform 1 0 3776 0 1 970
box -8 -3 16 105
use FILL  FILL_9308
timestamp 1680363874
transform 1 0 3784 0 1 970
box -8 -3 16 105
use FILL  FILL_9310
timestamp 1680363874
transform 1 0 3792 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_498
timestamp 1680363874
transform -1 0 3896 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7204
timestamp 1680363874
transform 1 0 3996 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_499
timestamp 1680363874
transform -1 0 3992 0 1 970
box -8 -3 104 105
use FILL  FILL_9311
timestamp 1680363874
transform 1 0 3992 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7205
timestamp 1680363874
transform 1 0 4020 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_501
timestamp 1680363874
transform 1 0 4000 0 1 970
box -8 -3 104 105
use INVX2  INVX2_566
timestamp 1680363874
transform 1 0 4096 0 1 970
box -9 -3 26 105
use FILL  FILL_9318
timestamp 1680363874
transform 1 0 4112 0 1 970
box -8 -3 16 105
use FILL  FILL_9319
timestamp 1680363874
transform 1 0 4120 0 1 970
box -8 -3 16 105
use FILL  FILL_9320
timestamp 1680363874
transform 1 0 4128 0 1 970
box -8 -3 16 105
use FILL  FILL_9321
timestamp 1680363874
transform 1 0 4136 0 1 970
box -8 -3 16 105
use FILL  FILL_9322
timestamp 1680363874
transform 1 0 4144 0 1 970
box -8 -3 16 105
use FILL  FILL_9323
timestamp 1680363874
transform 1 0 4152 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_314
timestamp 1680363874
transform 1 0 4160 0 1 970
box -8 -3 46 105
use FILL  FILL_9324
timestamp 1680363874
transform 1 0 4200 0 1 970
box -8 -3 16 105
use FILL  FILL_9325
timestamp 1680363874
transform 1 0 4208 0 1 970
box -8 -3 16 105
use FILL  FILL_9326
timestamp 1680363874
transform 1 0 4216 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_502
timestamp 1680363874
transform -1 0 4320 0 1 970
box -8 -3 104 105
use FILL  FILL_9327
timestamp 1680363874
transform 1 0 4320 0 1 970
box -8 -3 16 105
use FILL  FILL_9328
timestamp 1680363874
transform 1 0 4328 0 1 970
box -8 -3 16 105
use FILL  FILL_9329
timestamp 1680363874
transform 1 0 4336 0 1 970
box -8 -3 16 105
use FILL  FILL_9330
timestamp 1680363874
transform 1 0 4344 0 1 970
box -8 -3 16 105
use FILL  FILL_9331
timestamp 1680363874
transform 1 0 4352 0 1 970
box -8 -3 16 105
use FILL  FILL_9332
timestamp 1680363874
transform 1 0 4360 0 1 970
box -8 -3 16 105
use FILL  FILL_9333
timestamp 1680363874
transform 1 0 4368 0 1 970
box -8 -3 16 105
use FILL  FILL_9334
timestamp 1680363874
transform 1 0 4376 0 1 970
box -8 -3 16 105
use INVX2  INVX2_567
timestamp 1680363874
transform -1 0 4400 0 1 970
box -9 -3 26 105
use FILL  FILL_9335
timestamp 1680363874
transform 1 0 4400 0 1 970
box -8 -3 16 105
use FILL  FILL_9350
timestamp 1680363874
transform 1 0 4408 0 1 970
box -8 -3 16 105
use FILL  FILL_9352
timestamp 1680363874
transform 1 0 4416 0 1 970
box -8 -3 16 105
use FILL  FILL_9353
timestamp 1680363874
transform 1 0 4424 0 1 970
box -8 -3 16 105
use FILL  FILL_9354
timestamp 1680363874
transform 1 0 4432 0 1 970
box -8 -3 16 105
use FILL  FILL_9355
timestamp 1680363874
transform 1 0 4440 0 1 970
box -8 -3 16 105
use FILL  FILL_9358
timestamp 1680363874
transform 1 0 4448 0 1 970
box -8 -3 16 105
use FILL  FILL_9360
timestamp 1680363874
transform 1 0 4456 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_315
timestamp 1680363874
transform 1 0 4464 0 1 970
box -8 -3 46 105
use FILL  FILL_9362
timestamp 1680363874
transform 1 0 4504 0 1 970
box -8 -3 16 105
use FILL  FILL_9364
timestamp 1680363874
transform 1 0 4512 0 1 970
box -8 -3 16 105
use FILL  FILL_9366
timestamp 1680363874
transform 1 0 4520 0 1 970
box -8 -3 16 105
use FILL  FILL_9368
timestamp 1680363874
transform 1 0 4528 0 1 970
box -8 -3 16 105
use FILL  FILL_9370
timestamp 1680363874
transform 1 0 4536 0 1 970
box -8 -3 16 105
use FILL  FILL_9371
timestamp 1680363874
transform 1 0 4544 0 1 970
box -8 -3 16 105
use FILL  FILL_9372
timestamp 1680363874
transform 1 0 4552 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_358
timestamp 1680363874
transform 1 0 4560 0 1 970
box -8 -3 46 105
use FILL  FILL_9373
timestamp 1680363874
transform 1 0 4600 0 1 970
box -8 -3 16 105
use FILL  FILL_9374
timestamp 1680363874
transform 1 0 4608 0 1 970
box -8 -3 16 105
use FILL  FILL_9375
timestamp 1680363874
transform 1 0 4616 0 1 970
box -8 -3 16 105
use FILL  FILL_9376
timestamp 1680363874
transform 1 0 4624 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_317
timestamp 1680363874
transform 1 0 4632 0 1 970
box -8 -3 46 105
use FILL  FILL_9377
timestamp 1680363874
transform 1 0 4672 0 1 970
box -8 -3 16 105
use FILL  FILL_9384
timestamp 1680363874
transform 1 0 4680 0 1 970
box -8 -3 16 105
use FILL  FILL_9386
timestamp 1680363874
transform 1 0 4688 0 1 970
box -8 -3 16 105
use FILL  FILL_9387
timestamp 1680363874
transform 1 0 4696 0 1 970
box -8 -3 16 105
use FILL  FILL_9388
timestamp 1680363874
transform 1 0 4704 0 1 970
box -8 -3 16 105
use FILL  FILL_9389
timestamp 1680363874
transform 1 0 4712 0 1 970
box -8 -3 16 105
use FILL  FILL_9390
timestamp 1680363874
transform 1 0 4720 0 1 970
box -8 -3 16 105
use FILL  FILL_9391
timestamp 1680363874
transform 1 0 4728 0 1 970
box -8 -3 16 105
use FILL  FILL_9392
timestamp 1680363874
transform 1 0 4736 0 1 970
box -8 -3 16 105
use FILL  FILL_9393
timestamp 1680363874
transform 1 0 4744 0 1 970
box -8 -3 16 105
use FILL  FILL_9394
timestamp 1680363874
transform 1 0 4752 0 1 970
box -8 -3 16 105
use FILL  FILL_9395
timestamp 1680363874
transform 1 0 4760 0 1 970
box -8 -3 16 105
use FILL  FILL_9396
timestamp 1680363874
transform 1 0 4768 0 1 970
box -8 -3 16 105
use FILL  FILL_9397
timestamp 1680363874
transform 1 0 4776 0 1 970
box -8 -3 16 105
use FILL  FILL_9398
timestamp 1680363874
transform 1 0 4784 0 1 970
box -8 -3 16 105
use FILL  FILL_9399
timestamp 1680363874
transform 1 0 4792 0 1 970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_75
timestamp 1680363874
transform 1 0 4827 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_7270
timestamp 1680363874
transform 1 0 68 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8019
timestamp 1680363874
transform 1 0 68 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7392
timestamp 1680363874
transform 1 0 4 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7921
timestamp 1680363874
transform 1 0 164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8020
timestamp 1680363874
transform 1 0 124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8021
timestamp 1680363874
transform 1 0 196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7919
timestamp 1680363874
transform 1 0 212 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7271
timestamp 1680363874
transform 1 0 212 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7922
timestamp 1680363874
transform 1 0 220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8022
timestamp 1680363874
transform 1 0 220 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7229
timestamp 1680363874
transform 1 0 236 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7923
timestamp 1680363874
transform 1 0 244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8023
timestamp 1680363874
transform 1 0 236 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7272
timestamp 1680363874
transform 1 0 268 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8024
timestamp 1680363874
transform 1 0 260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8025
timestamp 1680363874
transform 1 0 268 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7352
timestamp 1680363874
transform 1 0 260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7377
timestamp 1680363874
transform 1 0 284 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7924
timestamp 1680363874
transform 1 0 292 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7230
timestamp 1680363874
transform 1 0 316 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7925
timestamp 1680363874
transform 1 0 316 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7231
timestamp 1680363874
transform 1 0 420 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7926
timestamp 1680363874
transform 1 0 420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8026
timestamp 1680363874
transform 1 0 316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8027
timestamp 1680363874
transform 1 0 324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8028
timestamp 1680363874
transform 1 0 340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8029
timestamp 1680363874
transform 1 0 372 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7312
timestamp 1680363874
transform 1 0 324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7286
timestamp 1680363874
transform 1 0 420 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7232
timestamp 1680363874
transform 1 0 476 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7233
timestamp 1680363874
transform 1 0 516 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7927
timestamp 1680363874
transform 1 0 516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8030
timestamp 1680363874
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8031
timestamp 1680363874
transform 1 0 468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8133
timestamp 1680363874
transform 1 0 332 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7313
timestamp 1680363874
transform 1 0 372 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7353
timestamp 1680363874
transform 1 0 332 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7378
timestamp 1680363874
transform 1 0 396 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7393
timestamp 1680363874
transform 1 0 404 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7394
timestamp 1680363874
transform 1 0 508 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7215
timestamp 1680363874
transform 1 0 636 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7234
timestamp 1680363874
transform 1 0 596 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7235
timestamp 1680363874
transform 1 0 652 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7928
timestamp 1680363874
transform 1 0 548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7929
timestamp 1680363874
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7930
timestamp 1680363874
transform 1 0 652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7931
timestamp 1680363874
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7932
timestamp 1680363874
transform 1 0 676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8032
timestamp 1680363874
transform 1 0 596 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7287
timestamp 1680363874
transform 1 0 628 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8033
timestamp 1680363874
transform 1 0 636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8034
timestamp 1680363874
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8035
timestamp 1680363874
transform 1 0 660 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7314
timestamp 1680363874
transform 1 0 636 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7395
timestamp 1680363874
transform 1 0 548 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7288
timestamp 1680363874
transform 1 0 668 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7354
timestamp 1680363874
transform 1 0 660 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7315
timestamp 1680363874
transform 1 0 676 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7379
timestamp 1680363874
transform 1 0 644 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7380
timestamp 1680363874
transform 1 0 668 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7216
timestamp 1680363874
transform 1 0 772 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7217
timestamp 1680363874
transform 1 0 796 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7236
timestamp 1680363874
transform 1 0 732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7237
timestamp 1680363874
transform 1 0 756 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7238
timestamp 1680363874
transform 1 0 780 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8036
timestamp 1680363874
transform 1 0 708 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7355
timestamp 1680363874
transform 1 0 708 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7933
timestamp 1680363874
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8037
timestamp 1680363874
transform 1 0 780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7356
timestamp 1680363874
transform 1 0 772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7396
timestamp 1680363874
transform 1 0 764 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7239
timestamp 1680363874
transform 1 0 852 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7934
timestamp 1680363874
transform 1 0 836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7935
timestamp 1680363874
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8038
timestamp 1680363874
transform 1 0 828 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8039
timestamp 1680363874
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8040
timestamp 1680363874
transform 1 0 860 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7397
timestamp 1680363874
transform 1 0 836 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7936
timestamp 1680363874
transform 1 0 876 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7937
timestamp 1680363874
transform 1 0 884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7938
timestamp 1680363874
transform 1 0 916 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7939
timestamp 1680363874
transform 1 0 932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8041
timestamp 1680363874
transform 1 0 924 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7398
timestamp 1680363874
transform 1 0 932 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7206
timestamp 1680363874
transform 1 0 1020 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7940
timestamp 1680363874
transform 1 0 964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8042
timestamp 1680363874
transform 1 0 988 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7357
timestamp 1680363874
transform 1 0 956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7358
timestamp 1680363874
transform 1 0 988 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7399
timestamp 1680363874
transform 1 0 988 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8043
timestamp 1680363874
transform 1 0 1052 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7207
timestamp 1680363874
transform 1 0 1076 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7941
timestamp 1680363874
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8044
timestamp 1680363874
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8045
timestamp 1680363874
transform 1 0 1156 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7359
timestamp 1680363874
transform 1 0 1068 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7360
timestamp 1680363874
transform 1 0 1100 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7361
timestamp 1680363874
transform 1 0 1124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7400
timestamp 1680363874
transform 1 0 1076 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7240
timestamp 1680363874
transform 1 0 1172 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7208
timestamp 1680363874
transform 1 0 1196 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7209
timestamp 1680363874
transform 1 0 1268 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7241
timestamp 1680363874
transform 1 0 1236 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7942
timestamp 1680363874
transform 1 0 1188 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7273
timestamp 1680363874
transform 1 0 1236 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7274
timestamp 1680363874
transform 1 0 1260 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8046
timestamp 1680363874
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7316
timestamp 1680363874
transform 1 0 1188 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7317
timestamp 1680363874
transform 1 0 1236 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7362
timestamp 1680363874
transform 1 0 1180 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7289
timestamp 1680363874
transform 1 0 1276 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8047
timestamp 1680363874
transform 1 0 1300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8048
timestamp 1680363874
transform 1 0 1308 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7218
timestamp 1680363874
transform 1 0 1380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7242
timestamp 1680363874
transform 1 0 1372 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7943
timestamp 1680363874
transform 1 0 1396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8049
timestamp 1680363874
transform 1 0 1372 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7318
timestamp 1680363874
transform 1 0 1396 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7944
timestamp 1680363874
transform 1 0 1412 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7290
timestamp 1680363874
transform 1 0 1412 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7243
timestamp 1680363874
transform 1 0 1460 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7945
timestamp 1680363874
transform 1 0 1460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7946
timestamp 1680363874
transform 1 0 1476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8050
timestamp 1680363874
transform 1 0 1452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8051
timestamp 1680363874
transform 1 0 1468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7363
timestamp 1680363874
transform 1 0 1468 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7920
timestamp 1680363874
transform 1 0 1500 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7219
timestamp 1680363874
transform 1 0 1548 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7244
timestamp 1680363874
transform 1 0 1564 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7947
timestamp 1680363874
transform 1 0 1516 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7275
timestamp 1680363874
transform 1 0 1596 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8052
timestamp 1680363874
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7319
timestamp 1680363874
transform 1 0 1516 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7401
timestamp 1680363874
transform 1 0 1572 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7276
timestamp 1680363874
transform 1 0 1612 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7220
timestamp 1680363874
transform 1 0 1652 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7245
timestamp 1680363874
transform 1 0 1636 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7948
timestamp 1680363874
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7277
timestamp 1680363874
transform 1 0 1628 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7949
timestamp 1680363874
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7950
timestamp 1680363874
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7951
timestamp 1680363874
transform 1 0 1660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8053
timestamp 1680363874
transform 1 0 1612 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7291
timestamp 1680363874
transform 1 0 1620 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8054
timestamp 1680363874
transform 1 0 1628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8055
timestamp 1680363874
transform 1 0 1644 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7320
timestamp 1680363874
transform 1 0 1612 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7364
timestamp 1680363874
transform 1 0 1644 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7321
timestamp 1680363874
transform 1 0 1660 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7278
timestamp 1680363874
transform 1 0 1692 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8056
timestamp 1680363874
transform 1 0 1692 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7210
timestamp 1680363874
transform 1 0 1724 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7952
timestamp 1680363874
transform 1 0 1748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7953
timestamp 1680363874
transform 1 0 1764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8057
timestamp 1680363874
transform 1 0 1740 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7365
timestamp 1680363874
transform 1 0 1740 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7402
timestamp 1680363874
transform 1 0 1732 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8058
timestamp 1680363874
transform 1 0 1772 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7279
timestamp 1680363874
transform 1 0 1788 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8059
timestamp 1680363874
transform 1 0 1788 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7322
timestamp 1680363874
transform 1 0 1788 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7954
timestamp 1680363874
transform 1 0 1804 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7292
timestamp 1680363874
transform 1 0 1804 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7211
timestamp 1680363874
transform 1 0 1820 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7955
timestamp 1680363874
transform 1 0 1820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7956
timestamp 1680363874
transform 1 0 1828 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7403
timestamp 1680363874
transform 1 0 1828 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7246
timestamp 1680363874
transform 1 0 1892 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7247
timestamp 1680363874
transform 1 0 1940 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7957
timestamp 1680363874
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8060
timestamp 1680363874
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7293
timestamp 1680363874
transform 1 0 1892 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8061
timestamp 1680363874
transform 1 0 1916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8062
timestamp 1680363874
transform 1 0 1972 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7323
timestamp 1680363874
transform 1 0 1876 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7324
timestamp 1680363874
transform 1 0 1956 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7366
timestamp 1680363874
transform 1 0 1868 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7404
timestamp 1680363874
transform 1 0 1980 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7958
timestamp 1680363874
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7248
timestamp 1680363874
transform 1 0 2028 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7959
timestamp 1680363874
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7960
timestamp 1680363874
transform 1 0 2044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8063
timestamp 1680363874
transform 1 0 2012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8064
timestamp 1680363874
transform 1 0 2036 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7367
timestamp 1680363874
transform 1 0 2012 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7961
timestamp 1680363874
transform 1 0 2076 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7221
timestamp 1680363874
transform 1 0 2140 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7249
timestamp 1680363874
transform 1 0 2124 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7962
timestamp 1680363874
transform 1 0 2100 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7294
timestamp 1680363874
transform 1 0 2100 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8065
timestamp 1680363874
transform 1 0 2124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8066
timestamp 1680363874
transform 1 0 2180 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7325
timestamp 1680363874
transform 1 0 2124 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7963
timestamp 1680363874
transform 1 0 2204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8134
timestamp 1680363874
transform 1 0 2204 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7326
timestamp 1680363874
transform 1 0 2228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7222
timestamp 1680363874
transform 1 0 2252 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8067
timestamp 1680363874
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8135
timestamp 1680363874
transform 1 0 2236 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7964
timestamp 1680363874
transform 1 0 2268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7965
timestamp 1680363874
transform 1 0 2284 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7966
timestamp 1680363874
transform 1 0 2372 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7295
timestamp 1680363874
transform 1 0 2276 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8068
timestamp 1680363874
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8069
timestamp 1680363874
transform 1 0 2348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8070
timestamp 1680363874
transform 1 0 2388 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7327
timestamp 1680363874
transform 1 0 2348 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7328
timestamp 1680363874
transform 1 0 2388 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7368
timestamp 1680363874
transform 1 0 2372 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7967
timestamp 1680363874
transform 1 0 2428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7968
timestamp 1680363874
transform 1 0 2436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7969
timestamp 1680363874
transform 1 0 2452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8071
timestamp 1680363874
transform 1 0 2428 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7296
timestamp 1680363874
transform 1 0 2436 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8072
timestamp 1680363874
transform 1 0 2444 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7297
timestamp 1680363874
transform 1 0 2452 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7381
timestamp 1680363874
transform 1 0 2428 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8136
timestamp 1680363874
transform 1 0 2476 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7223
timestamp 1680363874
transform 1 0 2492 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8073
timestamp 1680363874
transform 1 0 2492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7970
timestamp 1680363874
transform 1 0 2500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8074
timestamp 1680363874
transform 1 0 2516 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7250
timestamp 1680363874
transform 1 0 2532 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7971
timestamp 1680363874
transform 1 0 2532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7972
timestamp 1680363874
transform 1 0 2540 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7369
timestamp 1680363874
transform 1 0 2540 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7973
timestamp 1680363874
transform 1 0 2572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8075
timestamp 1680363874
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8137
timestamp 1680363874
transform 1 0 2580 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7382
timestamp 1680363874
transform 1 0 2580 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7974
timestamp 1680363874
transform 1 0 2612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7975
timestamp 1680363874
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8076
timestamp 1680363874
transform 1 0 2604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7298
timestamp 1680363874
transform 1 0 2612 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8077
timestamp 1680363874
transform 1 0 2620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7329
timestamp 1680363874
transform 1 0 2604 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7370
timestamp 1680363874
transform 1 0 2628 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7383
timestamp 1680363874
transform 1 0 2604 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7384
timestamp 1680363874
transform 1 0 2620 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7251
timestamp 1680363874
transform 1 0 2644 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7976
timestamp 1680363874
transform 1 0 2644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8078
timestamp 1680363874
transform 1 0 2660 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7299
timestamp 1680363874
transform 1 0 2676 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8079
timestamp 1680363874
transform 1 0 2684 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7330
timestamp 1680363874
transform 1 0 2684 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7977
timestamp 1680363874
transform 1 0 2716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7978
timestamp 1680363874
transform 1 0 2724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8080
timestamp 1680363874
transform 1 0 2708 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7300
timestamp 1680363874
transform 1 0 2716 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7224
timestamp 1680363874
transform 1 0 2788 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7979
timestamp 1680363874
transform 1 0 2772 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7301
timestamp 1680363874
transform 1 0 2772 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8081
timestamp 1680363874
transform 1 0 2796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8082
timestamp 1680363874
transform 1 0 2860 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7252
timestamp 1680363874
transform 1 0 2884 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7253
timestamp 1680363874
transform 1 0 2932 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7980
timestamp 1680363874
transform 1 0 2884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8083
timestamp 1680363874
transform 1 0 2916 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7331
timestamp 1680363874
transform 1 0 2932 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7405
timestamp 1680363874
transform 1 0 2884 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7981
timestamp 1680363874
transform 1 0 2972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8084
timestamp 1680363874
transform 1 0 2988 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7371
timestamp 1680363874
transform 1 0 3004 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8085
timestamp 1680363874
transform 1 0 3020 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7254
timestamp 1680363874
transform 1 0 3036 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7982
timestamp 1680363874
transform 1 0 3036 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7302
timestamp 1680363874
transform 1 0 3076 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8086
timestamp 1680363874
transform 1 0 3084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8087
timestamp 1680363874
transform 1 0 3116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8088
timestamp 1680363874
transform 1 0 3124 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7332
timestamp 1680363874
transform 1 0 3084 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7333
timestamp 1680363874
transform 1 0 3124 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7255
timestamp 1680363874
transform 1 0 3148 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7983
timestamp 1680363874
transform 1 0 3148 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7334
timestamp 1680363874
transform 1 0 3140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7385
timestamp 1680363874
transform 1 0 3132 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7256
timestamp 1680363874
transform 1 0 3172 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7984
timestamp 1680363874
transform 1 0 3236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8089
timestamp 1680363874
transform 1 0 3156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8090
timestamp 1680363874
transform 1 0 3212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7303
timestamp 1680363874
transform 1 0 3236 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7335
timestamp 1680363874
transform 1 0 3172 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7304
timestamp 1680363874
transform 1 0 3252 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7257
timestamp 1680363874
transform 1 0 3268 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7985
timestamp 1680363874
transform 1 0 3268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7986
timestamp 1680363874
transform 1 0 3292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7987
timestamp 1680363874
transform 1 0 3300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8091
timestamp 1680363874
transform 1 0 3268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8092
timestamp 1680363874
transform 1 0 3284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7305
timestamp 1680363874
transform 1 0 3292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8093
timestamp 1680363874
transform 1 0 3308 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7212
timestamp 1680363874
transform 1 0 3380 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7258
timestamp 1680363874
transform 1 0 3348 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7259
timestamp 1680363874
transform 1 0 3396 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7260
timestamp 1680363874
transform 1 0 3428 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7988
timestamp 1680363874
transform 1 0 3428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8094
timestamp 1680363874
transform 1 0 3340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8095
timestamp 1680363874
transform 1 0 3348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8096
timestamp 1680363874
transform 1 0 3388 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7336
timestamp 1680363874
transform 1 0 3340 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7406
timestamp 1680363874
transform 1 0 3332 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7306
timestamp 1680363874
transform 1 0 3428 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7337
timestamp 1680363874
transform 1 0 3388 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7386
timestamp 1680363874
transform 1 0 3364 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7387
timestamp 1680363874
transform 1 0 3388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7407
timestamp 1680363874
transform 1 0 3420 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7307
timestamp 1680363874
transform 1 0 3444 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7261
timestamp 1680363874
transform 1 0 3468 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8097
timestamp 1680363874
transform 1 0 3460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7262
timestamp 1680363874
transform 1 0 3524 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7989
timestamp 1680363874
transform 1 0 3516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7990
timestamp 1680363874
transform 1 0 3524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8098
timestamp 1680363874
transform 1 0 3524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8099
timestamp 1680363874
transform 1 0 3532 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7213
timestamp 1680363874
transform 1 0 3596 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7991
timestamp 1680363874
transform 1 0 3596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7992
timestamp 1680363874
transform 1 0 3612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8100
timestamp 1680363874
transform 1 0 3588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8101
timestamp 1680363874
transform 1 0 3604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7214
timestamp 1680363874
transform 1 0 3628 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8102
timestamp 1680363874
transform 1 0 3644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7993
timestamp 1680363874
transform 1 0 3668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8103
timestamp 1680363874
transform 1 0 3716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8104
timestamp 1680363874
transform 1 0 3724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7338
timestamp 1680363874
transform 1 0 3716 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7280
timestamp 1680363874
transform 1 0 3756 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8105
timestamp 1680363874
transform 1 0 3756 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7281
timestamp 1680363874
transform 1 0 3780 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8106
timestamp 1680363874
transform 1 0 3780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7225
timestamp 1680363874
transform 1 0 3820 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7263
timestamp 1680363874
transform 1 0 3812 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7994
timestamp 1680363874
transform 1 0 3812 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7388
timestamp 1680363874
transform 1 0 3804 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7339
timestamp 1680363874
transform 1 0 3820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7226
timestamp 1680363874
transform 1 0 3836 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7995
timestamp 1680363874
transform 1 0 3836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7996
timestamp 1680363874
transform 1 0 3844 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7282
timestamp 1680363874
transform 1 0 3860 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7227
timestamp 1680363874
transform 1 0 3940 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7264
timestamp 1680363874
transform 1 0 3948 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7265
timestamp 1680363874
transform 1 0 3972 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7997
timestamp 1680363874
transform 1 0 3868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7998
timestamp 1680363874
transform 1 0 3884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7999
timestamp 1680363874
transform 1 0 3972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8107
timestamp 1680363874
transform 1 0 3860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8108
timestamp 1680363874
transform 1 0 3876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8109
timestamp 1680363874
transform 1 0 3892 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8110
timestamp 1680363874
transform 1 0 3924 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7340
timestamp 1680363874
transform 1 0 3844 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7341
timestamp 1680363874
transform 1 0 3860 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7342
timestamp 1680363874
transform 1 0 3892 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7372
timestamp 1680363874
transform 1 0 3844 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7389
timestamp 1680363874
transform 1 0 3876 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8000
timestamp 1680363874
transform 1 0 3988 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7373
timestamp 1680363874
transform 1 0 3932 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7374
timestamp 1680363874
transform 1 0 3980 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7283
timestamp 1680363874
transform 1 0 3996 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8111
timestamp 1680363874
transform 1 0 3996 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7266
timestamp 1680363874
transform 1 0 4044 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8001
timestamp 1680363874
transform 1 0 4020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8002
timestamp 1680363874
transform 1 0 4036 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7308
timestamp 1680363874
transform 1 0 4020 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8112
timestamp 1680363874
transform 1 0 4028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8113
timestamp 1680363874
transform 1 0 4052 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7267
timestamp 1680363874
transform 1 0 4076 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7284
timestamp 1680363874
transform 1 0 4076 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8003
timestamp 1680363874
transform 1 0 4084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8004
timestamp 1680363874
transform 1 0 4124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8005
timestamp 1680363874
transform 1 0 4140 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7285
timestamp 1680363874
transform 1 0 4148 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8114
timestamp 1680363874
transform 1 0 4132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8115
timestamp 1680363874
transform 1 0 4148 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7343
timestamp 1680363874
transform 1 0 4132 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8006
timestamp 1680363874
transform 1 0 4164 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7228
timestamp 1680363874
transform 1 0 4204 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8007
timestamp 1680363874
transform 1 0 4204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8116
timestamp 1680363874
transform 1 0 4252 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7408
timestamp 1680363874
transform 1 0 4252 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8117
timestamp 1680363874
transform 1 0 4292 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7268
timestamp 1680363874
transform 1 0 4388 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8008
timestamp 1680363874
transform 1 0 4308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8118
timestamp 1680363874
transform 1 0 4356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8119
timestamp 1680363874
transform 1 0 4388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8120
timestamp 1680363874
transform 1 0 4396 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7344
timestamp 1680363874
transform 1 0 4356 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7409
timestamp 1680363874
transform 1 0 4316 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7345
timestamp 1680363874
transform 1 0 4396 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7390
timestamp 1680363874
transform 1 0 4396 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7269
timestamp 1680363874
transform 1 0 4492 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8009
timestamp 1680363874
transform 1 0 4460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8010
timestamp 1680363874
transform 1 0 4468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8011
timestamp 1680363874
transform 1 0 4476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8012
timestamp 1680363874
transform 1 0 4492 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7346
timestamp 1680363874
transform 1 0 4460 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8121
timestamp 1680363874
transform 1 0 4484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8122
timestamp 1680363874
transform 1 0 4500 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7347
timestamp 1680363874
transform 1 0 4484 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7375
timestamp 1680363874
transform 1 0 4476 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8123
timestamp 1680363874
transform 1 0 4524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8013
timestamp 1680363874
transform 1 0 4556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8124
timestamp 1680363874
transform 1 0 4548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8125
timestamp 1680363874
transform 1 0 4564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7391
timestamp 1680363874
transform 1 0 4564 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8014
timestamp 1680363874
transform 1 0 4588 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7309
timestamp 1680363874
transform 1 0 4588 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8126
timestamp 1680363874
transform 1 0 4596 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7376
timestamp 1680363874
transform 1 0 4596 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8015
timestamp 1680363874
transform 1 0 4612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8016
timestamp 1680363874
transform 1 0 4628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8017
timestamp 1680363874
transform 1 0 4636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8127
timestamp 1680363874
transform 1 0 4620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7310
timestamp 1680363874
transform 1 0 4628 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8128
timestamp 1680363874
transform 1 0 4636 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7348
timestamp 1680363874
transform 1 0 4620 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8129
timestamp 1680363874
transform 1 0 4652 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7349
timestamp 1680363874
transform 1 0 4644 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8018
timestamp 1680363874
transform 1 0 4780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8130
timestamp 1680363874
transform 1 0 4692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8131
timestamp 1680363874
transform 1 0 4700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7350
timestamp 1680363874
transform 1 0 4692 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7311
timestamp 1680363874
transform 1 0 4708 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8132
timestamp 1680363874
transform 1 0 4732 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7351
timestamp 1680363874
transform 1 0 4732 0 1 915
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_76
timestamp 1680363874
transform 1 0 24 0 1 870
box -10 -3 10 3
use FILL  FILL_8991
timestamp 1680363874
transform 1 0 72 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_469
timestamp 1680363874
transform -1 0 176 0 -1 970
box -8 -3 104 105
use FILL  FILL_8992
timestamp 1680363874
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_8994
timestamp 1680363874
transform 1 0 184 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_106
timestamp 1680363874
transform -1 0 216 0 -1 970
box -8 -3 32 105
use INVX2  INVX2_540
timestamp 1680363874
transform 1 0 216 0 -1 970
box -9 -3 26 105
use FILL  FILL_9025
timestamp 1680363874
transform 1 0 232 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_541
timestamp 1680363874
transform 1 0 240 0 -1 970
box -9 -3 26 105
use NAND2X1  NAND2X1_57
timestamp 1680363874
transform 1 0 256 0 -1 970
box -8 -3 32 105
use FILL  FILL_9026
timestamp 1680363874
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_9027
timestamp 1680363874
transform 1 0 288 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_542
timestamp 1680363874
transform 1 0 296 0 -1 970
box -9 -3 26 105
use NAND2X1  NAND2X1_58
timestamp 1680363874
transform 1 0 312 0 -1 970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_476
timestamp 1680363874
transform -1 0 432 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_477
timestamp 1680363874
transform -1 0 528 0 -1 970
box -8 -3 104 105
use FILL  FILL_9028
timestamp 1680363874
transform 1 0 528 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_478
timestamp 1680363874
transform 1 0 536 0 -1 970
box -8 -3 104 105
use OAI22X1  OAI22X1_343
timestamp 1680363874
transform 1 0 632 0 -1 970
box -8 -3 46 105
use FILL  FILL_9029
timestamp 1680363874
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9030
timestamp 1680363874
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_9031
timestamp 1680363874
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_9032
timestamp 1680363874
transform 1 0 696 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_543
timestamp 1680363874
transform 1 0 704 0 -1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_479
timestamp 1680363874
transform 1 0 720 0 -1 970
box -8 -3 104 105
use FILL  FILL_9033
timestamp 1680363874
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_9034
timestamp 1680363874
transform 1 0 824 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_344
timestamp 1680363874
transform -1 0 872 0 -1 970
box -8 -3 46 105
use FILL  FILL_9035
timestamp 1680363874
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_9036
timestamp 1680363874
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_9037
timestamp 1680363874
transform 1 0 888 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_345
timestamp 1680363874
transform 1 0 896 0 -1 970
box -8 -3 46 105
use FILL  FILL_9038
timestamp 1680363874
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_9039
timestamp 1680363874
transform 1 0 944 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_480
timestamp 1680363874
transform 1 0 952 0 -1 970
box -8 -3 104 105
use FILL  FILL_9040
timestamp 1680363874
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9041
timestamp 1680363874
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_481
timestamp 1680363874
transform 1 0 1064 0 -1 970
box -8 -3 104 105
use FILL  FILL_9042
timestamp 1680363874
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use FILL  FILL_9043
timestamp 1680363874
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7410
timestamp 1680363874
transform 1 0 1196 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7411
timestamp 1680363874
transform 1 0 1228 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_482
timestamp 1680363874
transform 1 0 1176 0 -1 970
box -8 -3 104 105
use FILL  FILL_9044
timestamp 1680363874
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_9045
timestamp 1680363874
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_9047
timestamp 1680363874
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_9049
timestamp 1680363874
transform 1 0 1296 0 -1 970
box -8 -3 16 105
use FILL  FILL_9060
timestamp 1680363874
transform 1 0 1304 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_483
timestamp 1680363874
transform -1 0 1408 0 -1 970
box -8 -3 104 105
use FILL  FILL_9061
timestamp 1680363874
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_9063
timestamp 1680363874
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_9075
timestamp 1680363874
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use FILL  FILL_9076
timestamp 1680363874
transform 1 0 1432 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_347
timestamp 1680363874
transform -1 0 1480 0 -1 970
box -8 -3 46 105
use FILL  FILL_9077
timestamp 1680363874
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_9078
timestamp 1680363874
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_9079
timestamp 1680363874
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_484
timestamp 1680363874
transform 1 0 1504 0 -1 970
box -8 -3 104 105
use FILL  FILL_9080
timestamp 1680363874
transform 1 0 1600 0 -1 970
box -8 -3 16 105
use FILL  FILL_9084
timestamp 1680363874
transform 1 0 1608 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_348
timestamp 1680363874
transform -1 0 1656 0 -1 970
box -8 -3 46 105
use FILL  FILL_9085
timestamp 1680363874
transform 1 0 1656 0 -1 970
box -8 -3 16 105
use FILL  FILL_9087
timestamp 1680363874
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9089
timestamp 1680363874
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9091
timestamp 1680363874
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_547
timestamp 1680363874
transform 1 0 1688 0 -1 970
box -9 -3 26 105
use FILL  FILL_9094
timestamp 1680363874
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_9095
timestamp 1680363874
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_9096
timestamp 1680363874
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_9097
timestamp 1680363874
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_9098
timestamp 1680363874
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_349
timestamp 1680363874
transform 1 0 1744 0 -1 970
box -8 -3 46 105
use FILL  FILL_9099
timestamp 1680363874
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_9100
timestamp 1680363874
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_9107
timestamp 1680363874
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_548
timestamp 1680363874
transform -1 0 1824 0 -1 970
box -9 -3 26 105
use FILL  FILL_9108
timestamp 1680363874
transform 1 0 1824 0 -1 970
box -8 -3 16 105
use FILL  FILL_9109
timestamp 1680363874
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use FILL  FILL_9110
timestamp 1680363874
transform 1 0 1840 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_86
timestamp 1680363874
transform -1 0 1872 0 -1 970
box -5 -3 28 105
use FILL  FILL_9111
timestamp 1680363874
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_486
timestamp 1680363874
transform 1 0 1880 0 -1 970
box -8 -3 104 105
use FILL  FILL_9118
timestamp 1680363874
transform 1 0 1976 0 -1 970
box -8 -3 16 105
use FILL  FILL_9120
timestamp 1680363874
transform 1 0 1984 0 -1 970
box -8 -3 16 105
use FILL  FILL_9122
timestamp 1680363874
transform 1 0 1992 0 -1 970
box -8 -3 16 105
use FILL  FILL_9125
timestamp 1680363874
transform 1 0 2000 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_352
timestamp 1680363874
transform 1 0 2008 0 -1 970
box -8 -3 46 105
use FILL  FILL_9126
timestamp 1680363874
transform 1 0 2048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9128
timestamp 1680363874
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_9130
timestamp 1680363874
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_9132
timestamp 1680363874
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_9134
timestamp 1680363874
transform 1 0 2080 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7412
timestamp 1680363874
transform 1 0 2108 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7413
timestamp 1680363874
transform 1 0 2164 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_487
timestamp 1680363874
transform 1 0 2088 0 -1 970
box -8 -3 104 105
use FILL  FILL_9142
timestamp 1680363874
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9149
timestamp 1680363874
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_156
timestamp 1680363874
transform -1 0 2232 0 -1 970
box -8 -3 34 105
use FILL  FILL_9150
timestamp 1680363874
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_9152
timestamp 1680363874
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_9154
timestamp 1680363874
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_9156
timestamp 1680363874
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9171
timestamp 1680363874
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_551
timestamp 1680363874
transform -1 0 2288 0 -1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_488
timestamp 1680363874
transform -1 0 2384 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_552
timestamp 1680363874
transform -1 0 2400 0 -1 970
box -9 -3 26 105
use FILL  FILL_9172
timestamp 1680363874
transform 1 0 2400 0 -1 970
box -8 -3 16 105
use FILL  FILL_9174
timestamp 1680363874
transform 1 0 2408 0 -1 970
box -8 -3 16 105
use FILL  FILL_9176
timestamp 1680363874
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_304
timestamp 1680363874
transform -1 0 2464 0 -1 970
box -8 -3 46 105
use FILL  FILL_9178
timestamp 1680363874
transform 1 0 2464 0 -1 970
box -8 -3 16 105
use FILL  FILL_9185
timestamp 1680363874
transform 1 0 2472 0 -1 970
box -8 -3 16 105
use FILL  FILL_9186
timestamp 1680363874
transform 1 0 2480 0 -1 970
box -8 -3 16 105
use FILL  FILL_9187
timestamp 1680363874
transform 1 0 2488 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_158
timestamp 1680363874
transform -1 0 2528 0 -1 970
box -8 -3 34 105
use FILL  FILL_9188
timestamp 1680363874
transform 1 0 2528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9193
timestamp 1680363874
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_87
timestamp 1680363874
transform -1 0 2568 0 -1 970
box -5 -3 28 105
use FILL  FILL_9194
timestamp 1680363874
transform 1 0 2568 0 -1 970
box -8 -3 16 105
use FILL  FILL_9195
timestamp 1680363874
transform 1 0 2576 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_305
timestamp 1680363874
transform -1 0 2624 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_555
timestamp 1680363874
transform 1 0 2624 0 -1 970
box -9 -3 26 105
use FILL  FILL_9196
timestamp 1680363874
transform 1 0 2640 0 -1 970
box -8 -3 16 105
use FILL  FILL_9197
timestamp 1680363874
transform 1 0 2648 0 -1 970
box -8 -3 16 105
use FILL  FILL_9198
timestamp 1680363874
transform 1 0 2656 0 -1 970
box -8 -3 16 105
use FILL  FILL_9199
timestamp 1680363874
transform 1 0 2664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9200
timestamp 1680363874
transform 1 0 2672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9208
timestamp 1680363874
transform 1 0 2680 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_306
timestamp 1680363874
transform -1 0 2728 0 -1 970
box -8 -3 46 105
use FILL  FILL_9209
timestamp 1680363874
transform 1 0 2728 0 -1 970
box -8 -3 16 105
use FILL  FILL_9225
timestamp 1680363874
transform 1 0 2736 0 -1 970
box -8 -3 16 105
use FILL  FILL_9226
timestamp 1680363874
transform 1 0 2744 0 -1 970
box -8 -3 16 105
use FILL  FILL_9227
timestamp 1680363874
transform 1 0 2752 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_490
timestamp 1680363874
transform 1 0 2760 0 -1 970
box -8 -3 104 105
use FILL  FILL_9228
timestamp 1680363874
transform 1 0 2856 0 -1 970
box -8 -3 16 105
use FILL  FILL_9229
timestamp 1680363874
transform 1 0 2864 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_491
timestamp 1680363874
transform 1 0 2872 0 -1 970
box -8 -3 104 105
use FILL  FILL_9230
timestamp 1680363874
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use FILL  FILL_9231
timestamp 1680363874
transform 1 0 2976 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_558
timestamp 1680363874
transform 1 0 2984 0 -1 970
box -9 -3 26 105
use FILL  FILL_9232
timestamp 1680363874
transform 1 0 3000 0 -1 970
box -8 -3 16 105
use FILL  FILL_9234
timestamp 1680363874
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use FILL  FILL_9236
timestamp 1680363874
transform 1 0 3016 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7414
timestamp 1680363874
transform 1 0 3060 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_492
timestamp 1680363874
transform 1 0 3024 0 -1 970
box -8 -3 104 105
use FILL  FILL_9261
timestamp 1680363874
transform 1 0 3120 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_560
timestamp 1680363874
transform -1 0 3144 0 -1 970
box -9 -3 26 105
use FILL  FILL_9262
timestamp 1680363874
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_493
timestamp 1680363874
transform -1 0 3248 0 -1 970
box -8 -3 104 105
use FILL  FILL_9263
timestamp 1680363874
transform 1 0 3248 0 -1 970
box -8 -3 16 105
use FILL  FILL_9264
timestamp 1680363874
transform 1 0 3256 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_311
timestamp 1680363874
transform -1 0 3304 0 -1 970
box -8 -3 46 105
use FILL  FILL_9265
timestamp 1680363874
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_9271
timestamp 1680363874
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_562
timestamp 1680363874
transform 1 0 3320 0 -1 970
box -9 -3 26 105
use FILL  FILL_9272
timestamp 1680363874
transform 1 0 3336 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7415
timestamp 1680363874
transform 1 0 3380 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_496
timestamp 1680363874
transform -1 0 3440 0 -1 970
box -8 -3 104 105
use FILL  FILL_9273
timestamp 1680363874
transform 1 0 3440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9274
timestamp 1680363874
transform 1 0 3448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9275
timestamp 1680363874
transform 1 0 3456 0 -1 970
box -8 -3 16 105
use FILL  FILL_9276
timestamp 1680363874
transform 1 0 3464 0 -1 970
box -8 -3 16 105
use FILL  FILL_9277
timestamp 1680363874
transform 1 0 3472 0 -1 970
box -8 -3 16 105
use FILL  FILL_9278
timestamp 1680363874
transform 1 0 3480 0 -1 970
box -8 -3 16 105
use FILL  FILL_9279
timestamp 1680363874
transform 1 0 3488 0 -1 970
box -8 -3 16 105
use FILL  FILL_9280
timestamp 1680363874
transform 1 0 3496 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_563
timestamp 1680363874
transform -1 0 3520 0 -1 970
box -9 -3 26 105
use FILL  FILL_9281
timestamp 1680363874
transform 1 0 3520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9282
timestamp 1680363874
transform 1 0 3528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9283
timestamp 1680363874
transform 1 0 3536 0 -1 970
box -8 -3 16 105
use FILL  FILL_9284
timestamp 1680363874
transform 1 0 3544 0 -1 970
box -8 -3 16 105
use FILL  FILL_9285
timestamp 1680363874
transform 1 0 3552 0 -1 970
box -8 -3 16 105
use FILL  FILL_9286
timestamp 1680363874
transform 1 0 3560 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_313
timestamp 1680363874
transform -1 0 3608 0 -1 970
box -8 -3 46 105
use FILL  FILL_9287
timestamp 1680363874
transform 1 0 3608 0 -1 970
box -8 -3 16 105
use FILL  FILL_9288
timestamp 1680363874
transform 1 0 3616 0 -1 970
box -8 -3 16 105
use FILL  FILL_9289
timestamp 1680363874
transform 1 0 3624 0 -1 970
box -8 -3 16 105
use FILL  FILL_9290
timestamp 1680363874
transform 1 0 3632 0 -1 970
box -8 -3 16 105
use FILL  FILL_9292
timestamp 1680363874
transform 1 0 3640 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_564
timestamp 1680363874
transform 1 0 3648 0 -1 970
box -9 -3 26 105
use FILL  FILL_9298
timestamp 1680363874
transform 1 0 3664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9299
timestamp 1680363874
transform 1 0 3672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9300
timestamp 1680363874
transform 1 0 3680 0 -1 970
box -8 -3 16 105
use FILL  FILL_9301
timestamp 1680363874
transform 1 0 3688 0 -1 970
box -8 -3 16 105
use FILL  FILL_9302
timestamp 1680363874
transform 1 0 3696 0 -1 970
box -8 -3 16 105
use FILL  FILL_9303
timestamp 1680363874
transform 1 0 3704 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_565
timestamp 1680363874
transform 1 0 3712 0 -1 970
box -9 -3 26 105
use FILL  FILL_9304
timestamp 1680363874
transform 1 0 3728 0 -1 970
box -8 -3 16 105
use FILL  FILL_9305
timestamp 1680363874
transform 1 0 3736 0 -1 970
box -8 -3 16 105
use FILL  FILL_9306
timestamp 1680363874
transform 1 0 3744 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_88
timestamp 1680363874
transform 1 0 3752 0 -1 970
box -5 -3 28 105
use FILL  FILL_9307
timestamp 1680363874
transform 1 0 3776 0 -1 970
box -8 -3 16 105
use FILL  FILL_9309
timestamp 1680363874
transform 1 0 3784 0 -1 970
box -8 -3 16 105
use FILL  FILL_9312
timestamp 1680363874
transform 1 0 3792 0 -1 970
box -8 -3 16 105
use FILL  FILL_9313
timestamp 1680363874
transform 1 0 3800 0 -1 970
box -8 -3 16 105
use FILL  FILL_9314
timestamp 1680363874
transform 1 0 3808 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_89
timestamp 1680363874
transform 1 0 3816 0 -1 970
box -5 -3 28 105
use FILL  FILL_9315
timestamp 1680363874
transform 1 0 3840 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_355
timestamp 1680363874
transform 1 0 3848 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_500
timestamp 1680363874
transform -1 0 3984 0 -1 970
box -8 -3 104 105
use FILL  FILL_9316
timestamp 1680363874
transform 1 0 3984 0 -1 970
box -8 -3 16 105
use FILL  FILL_9317
timestamp 1680363874
transform 1 0 3992 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_356
timestamp 1680363874
transform 1 0 4000 0 -1 970
box -8 -3 46 105
use FILL  FILL_9336
timestamp 1680363874
transform 1 0 4040 0 -1 970
box -8 -3 16 105
use FILL  FILL_9337
timestamp 1680363874
transform 1 0 4048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9338
timestamp 1680363874
transform 1 0 4056 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_90
timestamp 1680363874
transform 1 0 4064 0 -1 970
box -5 -3 28 105
use FILL  FILL_9339
timestamp 1680363874
transform 1 0 4088 0 -1 970
box -8 -3 16 105
use FILL  FILL_9340
timestamp 1680363874
transform 1 0 4096 0 -1 970
box -8 -3 16 105
use FILL  FILL_9341
timestamp 1680363874
transform 1 0 4104 0 -1 970
box -8 -3 16 105
use FILL  FILL_9342
timestamp 1680363874
transform 1 0 4112 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_357
timestamp 1680363874
transform -1 0 4160 0 -1 970
box -8 -3 46 105
use FILL  FILL_9343
timestamp 1680363874
transform 1 0 4160 0 -1 970
box -8 -3 16 105
use FILL  FILL_9344
timestamp 1680363874
transform 1 0 4168 0 -1 970
box -8 -3 16 105
use FILL  FILL_9345
timestamp 1680363874
transform 1 0 4176 0 -1 970
box -8 -3 16 105
use FILL  FILL_9346
timestamp 1680363874
transform 1 0 4184 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_503
timestamp 1680363874
transform 1 0 4192 0 -1 970
box -8 -3 104 105
use FILL  FILL_9347
timestamp 1680363874
transform 1 0 4288 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_504
timestamp 1680363874
transform 1 0 4296 0 -1 970
box -8 -3 104 105
use FILL  FILL_9348
timestamp 1680363874
transform 1 0 4392 0 -1 970
box -8 -3 16 105
use FILL  FILL_9349
timestamp 1680363874
transform 1 0 4400 0 -1 970
box -8 -3 16 105
use FILL  FILL_9351
timestamp 1680363874
transform 1 0 4408 0 -1 970
box -8 -3 16 105
use FILL  FILL_9356
timestamp 1680363874
transform 1 0 4416 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_568
timestamp 1680363874
transform -1 0 4440 0 -1 970
box -9 -3 26 105
use FILL  FILL_9357
timestamp 1680363874
transform 1 0 4440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9359
timestamp 1680363874
transform 1 0 4448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9361
timestamp 1680363874
transform 1 0 4456 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_316
timestamp 1680363874
transform 1 0 4464 0 -1 970
box -8 -3 46 105
use FILL  FILL_9363
timestamp 1680363874
transform 1 0 4504 0 -1 970
box -8 -3 16 105
use FILL  FILL_9365
timestamp 1680363874
transform 1 0 4512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9367
timestamp 1680363874
transform 1 0 4520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9369
timestamp 1680363874
transform 1 0 4528 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_359
timestamp 1680363874
transform 1 0 4536 0 -1 970
box -8 -3 46 105
use FILL  FILL_9378
timestamp 1680363874
transform 1 0 4576 0 -1 970
box -8 -3 16 105
use FILL  FILL_9379
timestamp 1680363874
transform 1 0 4584 0 -1 970
box -8 -3 16 105
use FILL  FILL_9380
timestamp 1680363874
transform 1 0 4592 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_318
timestamp 1680363874
transform 1 0 4600 0 -1 970
box -8 -3 46 105
use FILL  FILL_9381
timestamp 1680363874
transform 1 0 4640 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_569
timestamp 1680363874
transform 1 0 4648 0 -1 970
box -9 -3 26 105
use FILL  FILL_9382
timestamp 1680363874
transform 1 0 4664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9383
timestamp 1680363874
transform 1 0 4672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9385
timestamp 1680363874
transform 1 0 4680 0 -1 970
box -8 -3 16 105
use FILL  FILL_9400
timestamp 1680363874
transform 1 0 4688 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_505
timestamp 1680363874
transform -1 0 4792 0 -1 970
box -8 -3 104 105
use FILL  FILL_9401
timestamp 1680363874
transform 1 0 4792 0 -1 970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_77
timestamp 1680363874
transform 1 0 4851 0 1 870
box -10 -3 10 3
use M2_M1  M2_M1_8149
timestamp 1680363874
transform 1 0 76 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8150
timestamp 1680363874
transform 1 0 124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8281
timestamp 1680363874
transform 1 0 164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8282
timestamp 1680363874
transform 1 0 244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8140
timestamp 1680363874
transform 1 0 268 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7464
timestamp 1680363874
transform 1 0 316 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8151
timestamp 1680363874
transform 1 0 316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8283
timestamp 1680363874
transform 1 0 308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8141
timestamp 1680363874
transform 1 0 332 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7465
timestamp 1680363874
transform 1 0 356 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8152
timestamp 1680363874
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8284
timestamp 1680363874
transform 1 0 356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8389
timestamp 1680363874
transform 1 0 372 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_8153
timestamp 1680363874
transform 1 0 396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8285
timestamp 1680363874
transform 1 0 396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8286
timestamp 1680363874
transform 1 0 404 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7545
timestamp 1680363874
transform 1 0 396 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8154
timestamp 1680363874
transform 1 0 420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8155
timestamp 1680363874
transform 1 0 428 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7524
timestamp 1680363874
transform 1 0 420 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7525
timestamp 1680363874
transform 1 0 444 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7505
timestamp 1680363874
transform 1 0 476 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8156
timestamp 1680363874
transform 1 0 500 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7506
timestamp 1680363874
transform 1 0 548 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8287
timestamp 1680363874
transform 1 0 548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7546
timestamp 1680363874
transform 1 0 500 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8157
timestamp 1680363874
transform 1 0 620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8158
timestamp 1680363874
transform 1 0 676 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7507
timestamp 1680363874
transform 1 0 700 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8288
timestamp 1680363874
transform 1 0 700 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7547
timestamp 1680363874
transform 1 0 676 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8289
timestamp 1680363874
transform 1 0 716 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7445
timestamp 1680363874
transform 1 0 740 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7508
timestamp 1680363874
transform 1 0 732 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8159
timestamp 1680363874
transform 1 0 740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8160
timestamp 1680363874
transform 1 0 756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8290
timestamp 1680363874
transform 1 0 748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8291
timestamp 1680363874
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8292
timestamp 1680363874
transform 1 0 772 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7548
timestamp 1680363874
transform 1 0 748 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7420
timestamp 1680363874
transform 1 0 780 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7446
timestamp 1680363874
transform 1 0 804 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7466
timestamp 1680363874
transform 1 0 812 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8161
timestamp 1680363874
transform 1 0 796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8162
timestamp 1680363874
transform 1 0 812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8293
timestamp 1680363874
transform 1 0 820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8294
timestamp 1680363874
transform 1 0 828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8295
timestamp 1680363874
transform 1 0 836 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7447
timestamp 1680363874
transform 1 0 860 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8163
timestamp 1680363874
transform 1 0 852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8142
timestamp 1680363874
transform 1 0 868 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7421
timestamp 1680363874
transform 1 0 884 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7436
timestamp 1680363874
transform 1 0 892 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8138
timestamp 1680363874
transform 1 0 892 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_7467
timestamp 1680363874
transform 1 0 884 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7448
timestamp 1680363874
transform 1 0 908 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8143
timestamp 1680363874
transform 1 0 900 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8164
timestamp 1680363874
transform 1 0 884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8165
timestamp 1680363874
transform 1 0 908 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7526
timestamp 1680363874
transform 1 0 908 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7422
timestamp 1680363874
transform 1 0 940 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8166
timestamp 1680363874
transform 1 0 964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8296
timestamp 1680363874
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8297
timestamp 1680363874
transform 1 0 956 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8167
timestamp 1680363874
transform 1 0 980 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7449
timestamp 1680363874
transform 1 0 996 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8298
timestamp 1680363874
transform 1 0 988 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7549
timestamp 1680363874
transform 1 0 988 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7423
timestamp 1680363874
transform 1 0 1060 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7450
timestamp 1680363874
transform 1 0 1060 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8168
timestamp 1680363874
transform 1 0 1052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8169
timestamp 1680363874
transform 1 0 1060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8170
timestamp 1680363874
transform 1 0 1076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8171
timestamp 1680363874
transform 1 0 1092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8299
timestamp 1680363874
transform 1 0 1052 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8300
timestamp 1680363874
transform 1 0 1068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8301
timestamp 1680363874
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7550
timestamp 1680363874
transform 1 0 1084 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7424
timestamp 1680363874
transform 1 0 1100 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7527
timestamp 1680363874
transform 1 0 1108 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8172
timestamp 1680363874
transform 1 0 1148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8302
timestamp 1680363874
transform 1 0 1156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8303
timestamp 1680363874
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8173
timestamp 1680363874
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7425
timestamp 1680363874
transform 1 0 1252 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8174
timestamp 1680363874
transform 1 0 1260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8304
timestamp 1680363874
transform 1 0 1236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8175
timestamp 1680363874
transform 1 0 1324 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7509
timestamp 1680363874
transform 1 0 1348 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8176
timestamp 1680363874
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8305
timestamp 1680363874
transform 1 0 1348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7551
timestamp 1680363874
transform 1 0 1396 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8306
timestamp 1680363874
transform 1 0 1460 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7426
timestamp 1680363874
transform 1 0 1500 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7468
timestamp 1680363874
transform 1 0 1492 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7469
timestamp 1680363874
transform 1 0 1516 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8177
timestamp 1680363874
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8178
timestamp 1680363874
transform 1 0 1500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8179
timestamp 1680363874
transform 1 0 1516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8307
timestamp 1680363874
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8308
timestamp 1680363874
transform 1 0 1508 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7552
timestamp 1680363874
transform 1 0 1508 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8309
timestamp 1680363874
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7570
timestamp 1680363874
transform 1 0 1540 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7427
timestamp 1680363874
transform 1 0 1668 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7428
timestamp 1680363874
transform 1 0 1684 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7470
timestamp 1680363874
transform 1 0 1660 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8180
timestamp 1680363874
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8181
timestamp 1680363874
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8182
timestamp 1680363874
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8183
timestamp 1680363874
transform 1 0 1684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8310
timestamp 1680363874
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7528
timestamp 1680363874
transform 1 0 1620 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8311
timestamp 1680363874
transform 1 0 1660 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7553
timestamp 1680363874
transform 1 0 1572 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7554
timestamp 1680363874
transform 1 0 1596 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7529
timestamp 1680363874
transform 1 0 1668 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8184
timestamp 1680363874
transform 1 0 1700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8312
timestamp 1680363874
transform 1 0 1676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8313
timestamp 1680363874
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7571
timestamp 1680363874
transform 1 0 1692 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7471
timestamp 1680363874
transform 1 0 1732 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8185
timestamp 1680363874
transform 1 0 1740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8314
timestamp 1680363874
transform 1 0 1732 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7555
timestamp 1680363874
transform 1 0 1732 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7530
timestamp 1680363874
transform 1 0 1748 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7472
timestamp 1680363874
transform 1 0 1764 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7437
timestamp 1680363874
transform 1 0 1780 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8144
timestamp 1680363874
transform 1 0 1772 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7531
timestamp 1680363874
transform 1 0 1764 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7416
timestamp 1680363874
transform 1 0 1820 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7417
timestamp 1680363874
transform 1 0 1836 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7438
timestamp 1680363874
transform 1 0 1812 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8139
timestamp 1680363874
transform 1 0 1812 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_8145
timestamp 1680363874
transform 1 0 1820 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7473
timestamp 1680363874
transform 1 0 1860 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8186
timestamp 1680363874
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8187
timestamp 1680363874
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8188
timestamp 1680363874
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7556
timestamp 1680363874
transform 1 0 1804 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7572
timestamp 1680363874
transform 1 0 1812 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8315
timestamp 1680363874
transform 1 0 1908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8316
timestamp 1680363874
transform 1 0 1924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8189
timestamp 1680363874
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7510
timestamp 1680363874
transform 1 0 1980 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8317
timestamp 1680363874
transform 1 0 1980 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7557
timestamp 1680363874
transform 1 0 1996 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7418
timestamp 1680363874
transform 1 0 2028 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7474
timestamp 1680363874
transform 1 0 2020 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8190
timestamp 1680363874
transform 1 0 2012 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7475
timestamp 1680363874
transform 1 0 2052 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8191
timestamp 1680363874
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8318
timestamp 1680363874
transform 1 0 2020 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8319
timestamp 1680363874
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7532
timestamp 1680363874
transform 1 0 2044 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8192
timestamp 1680363874
transform 1 0 2060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8320
timestamp 1680363874
transform 1 0 2060 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7558
timestamp 1680363874
transform 1 0 2052 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7533
timestamp 1680363874
transform 1 0 2068 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8321
timestamp 1680363874
transform 1 0 2084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8322
timestamp 1680363874
transform 1 0 2092 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7559
timestamp 1680363874
transform 1 0 2116 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8390
timestamp 1680363874
transform 1 0 2132 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7419
timestamp 1680363874
transform 1 0 2236 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7439
timestamp 1680363874
transform 1 0 2236 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7476
timestamp 1680363874
transform 1 0 2212 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8193
timestamp 1680363874
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8194
timestamp 1680363874
transform 1 0 2156 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8195
timestamp 1680363874
transform 1 0 2212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8196
timestamp 1680363874
transform 1 0 2252 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7534
timestamp 1680363874
transform 1 0 2172 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7429
timestamp 1680363874
transform 1 0 2292 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8146
timestamp 1680363874
transform 1 0 2276 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8323
timestamp 1680363874
transform 1 0 2236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8324
timestamp 1680363874
transform 1 0 2252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8325
timestamp 1680363874
transform 1 0 2268 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7560
timestamp 1680363874
transform 1 0 2196 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8391
timestamp 1680363874
transform 1 0 2268 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7573
timestamp 1680363874
transform 1 0 2252 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7477
timestamp 1680363874
transform 1 0 2300 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8197
timestamp 1680363874
transform 1 0 2292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8198
timestamp 1680363874
transform 1 0 2300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8326
timestamp 1680363874
transform 1 0 2308 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7440
timestamp 1680363874
transform 1 0 2372 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7478
timestamp 1680363874
transform 1 0 2380 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8199
timestamp 1680363874
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8327
timestamp 1680363874
transform 1 0 2340 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7511
timestamp 1680363874
transform 1 0 2356 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8200
timestamp 1680363874
transform 1 0 2364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8328
timestamp 1680363874
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7535
timestamp 1680363874
transform 1 0 2364 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8329
timestamp 1680363874
transform 1 0 2372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7574
timestamp 1680363874
transform 1 0 2372 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7575
timestamp 1680363874
transform 1 0 2396 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7479
timestamp 1680363874
transform 1 0 2452 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8201
timestamp 1680363874
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8202
timestamp 1680363874
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8330
timestamp 1680363874
transform 1 0 2420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8331
timestamp 1680363874
transform 1 0 2452 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7451
timestamp 1680363874
transform 1 0 2468 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8332
timestamp 1680363874
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8203
timestamp 1680363874
transform 1 0 2492 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7536
timestamp 1680363874
transform 1 0 2500 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8392
timestamp 1680363874
transform 1 0 2500 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7430
timestamp 1680363874
transform 1 0 2540 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8147
timestamp 1680363874
transform 1 0 2524 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8204
timestamp 1680363874
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8148
timestamp 1680363874
transform 1 0 2564 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7480
timestamp 1680363874
transform 1 0 2572 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8333
timestamp 1680363874
transform 1 0 2572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8205
timestamp 1680363874
transform 1 0 2596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8334
timestamp 1680363874
transform 1 0 2580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8335
timestamp 1680363874
transform 1 0 2612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7576
timestamp 1680363874
transform 1 0 2612 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7481
timestamp 1680363874
transform 1 0 2708 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8206
timestamp 1680363874
transform 1 0 2660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8207
timestamp 1680363874
transform 1 0 2708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8336
timestamp 1680363874
transform 1 0 2628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7577
timestamp 1680363874
transform 1 0 2644 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7578
timestamp 1680363874
transform 1 0 2700 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7452
timestamp 1680363874
transform 1 0 2788 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7482
timestamp 1680363874
transform 1 0 2796 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7483
timestamp 1680363874
transform 1 0 2836 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8208
timestamp 1680363874
transform 1 0 2796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8209
timestamp 1680363874
transform 1 0 2828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8210
timestamp 1680363874
transform 1 0 2836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8337
timestamp 1680363874
transform 1 0 2748 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7512
timestamp 1680363874
transform 1 0 2844 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8211
timestamp 1680363874
transform 1 0 2852 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7579
timestamp 1680363874
transform 1 0 2828 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7484
timestamp 1680363874
transform 1 0 2892 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8212
timestamp 1680363874
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7513
timestamp 1680363874
transform 1 0 2900 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8213
timestamp 1680363874
transform 1 0 2916 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7514
timestamp 1680363874
transform 1 0 2924 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8338
timestamp 1680363874
transform 1 0 2900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8339
timestamp 1680363874
transform 1 0 2908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8340
timestamp 1680363874
transform 1 0 2924 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7580
timestamp 1680363874
transform 1 0 2924 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7485
timestamp 1680363874
transform 1 0 2956 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7453
timestamp 1680363874
transform 1 0 3012 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7454
timestamp 1680363874
transform 1 0 3092 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7455
timestamp 1680363874
transform 1 0 3132 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7486
timestamp 1680363874
transform 1 0 3124 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7487
timestamp 1680363874
transform 1 0 3156 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8214
timestamp 1680363874
transform 1 0 2948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8215
timestamp 1680363874
transform 1 0 2956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8216
timestamp 1680363874
transform 1 0 2972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8217
timestamp 1680363874
transform 1 0 2988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8218
timestamp 1680363874
transform 1 0 2996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8219
timestamp 1680363874
transform 1 0 3028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8220
timestamp 1680363874
transform 1 0 3092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8221
timestamp 1680363874
transform 1 0 3116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8222
timestamp 1680363874
transform 1 0 3132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8223
timestamp 1680363874
transform 1 0 3148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8224
timestamp 1680363874
transform 1 0 3164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8341
timestamp 1680363874
transform 1 0 2964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8342
timestamp 1680363874
transform 1 0 2980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8343
timestamp 1680363874
transform 1 0 3076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8344
timestamp 1680363874
transform 1 0 3092 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7537
timestamp 1680363874
transform 1 0 3100 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8345
timestamp 1680363874
transform 1 0 3108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8346
timestamp 1680363874
transform 1 0 3124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8347
timestamp 1680363874
transform 1 0 3132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8348
timestamp 1680363874
transform 1 0 3156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8349
timestamp 1680363874
transform 1 0 3164 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7581
timestamp 1680363874
transform 1 0 3092 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8225
timestamp 1680363874
transform 1 0 3196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8226
timestamp 1680363874
transform 1 0 3212 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7456
timestamp 1680363874
transform 1 0 3228 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8227
timestamp 1680363874
transform 1 0 3228 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7431
timestamp 1680363874
transform 1 0 3364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7457
timestamp 1680363874
transform 1 0 3300 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8228
timestamp 1680363874
transform 1 0 3260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8229
timestamp 1680363874
transform 1 0 3276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8230
timestamp 1680363874
transform 1 0 3284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8231
timestamp 1680363874
transform 1 0 3340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8232
timestamp 1680363874
transform 1 0 3380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8350
timestamp 1680363874
transform 1 0 3252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8351
timestamp 1680363874
transform 1 0 3268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8352
timestamp 1680363874
transform 1 0 3364 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7582
timestamp 1680363874
transform 1 0 3268 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7583
timestamp 1680363874
transform 1 0 3284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7432
timestamp 1680363874
transform 1 0 3428 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7441
timestamp 1680363874
transform 1 0 3500 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7442
timestamp 1680363874
transform 1 0 3524 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7458
timestamp 1680363874
transform 1 0 3524 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7488
timestamp 1680363874
transform 1 0 3532 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8233
timestamp 1680363874
transform 1 0 3404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8234
timestamp 1680363874
transform 1 0 3460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8235
timestamp 1680363874
transform 1 0 3500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8236
timestamp 1680363874
transform 1 0 3516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8237
timestamp 1680363874
transform 1 0 3532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8238
timestamp 1680363874
transform 1 0 3540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8353
timestamp 1680363874
transform 1 0 3396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8354
timestamp 1680363874
transform 1 0 3484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8355
timestamp 1680363874
transform 1 0 3500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8356
timestamp 1680363874
transform 1 0 3524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8357
timestamp 1680363874
transform 1 0 3532 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7584
timestamp 1680363874
transform 1 0 3404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7585
timestamp 1680363874
transform 1 0 3500 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7538
timestamp 1680363874
transform 1 0 3540 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7443
timestamp 1680363874
transform 1 0 3556 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7444
timestamp 1680363874
transform 1 0 3580 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8239
timestamp 1680363874
transform 1 0 3572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8358
timestamp 1680363874
transform 1 0 3580 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7586
timestamp 1680363874
transform 1 0 3564 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7489
timestamp 1680363874
transform 1 0 3604 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8240
timestamp 1680363874
transform 1 0 3596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8241
timestamp 1680363874
transform 1 0 3604 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7459
timestamp 1680363874
transform 1 0 3620 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8242
timestamp 1680363874
transform 1 0 3620 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7561
timestamp 1680363874
transform 1 0 3612 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7490
timestamp 1680363874
transform 1 0 3636 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8243
timestamp 1680363874
transform 1 0 3636 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7491
timestamp 1680363874
transform 1 0 3668 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8244
timestamp 1680363874
transform 1 0 3660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8245
timestamp 1680363874
transform 1 0 3676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8359
timestamp 1680363874
transform 1 0 3652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8360
timestamp 1680363874
transform 1 0 3668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8361
timestamp 1680363874
transform 1 0 3684 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8362
timestamp 1680363874
transform 1 0 3700 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7492
timestamp 1680363874
transform 1 0 3764 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8246
timestamp 1680363874
transform 1 0 3764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8247
timestamp 1680363874
transform 1 0 3780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8248
timestamp 1680363874
transform 1 0 3796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8363
timestamp 1680363874
transform 1 0 3764 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7539
timestamp 1680363874
transform 1 0 3796 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7493
timestamp 1680363874
transform 1 0 3828 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8249
timestamp 1680363874
transform 1 0 3828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8364
timestamp 1680363874
transform 1 0 3820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8365
timestamp 1680363874
transform 1 0 3828 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7587
timestamp 1680363874
transform 1 0 3828 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7494
timestamp 1680363874
transform 1 0 3852 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8250
timestamp 1680363874
transform 1 0 3852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8366
timestamp 1680363874
transform 1 0 3860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8367
timestamp 1680363874
transform 1 0 3868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8251
timestamp 1680363874
transform 1 0 3908 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7562
timestamp 1680363874
transform 1 0 3908 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8252
timestamp 1680363874
transform 1 0 3924 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7460
timestamp 1680363874
transform 1 0 4028 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7495
timestamp 1680363874
transform 1 0 3996 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7496
timestamp 1680363874
transform 1 0 4036 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8253
timestamp 1680363874
transform 1 0 3996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8254
timestamp 1680363874
transform 1 0 4028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8255
timestamp 1680363874
transform 1 0 4036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8368
timestamp 1680363874
transform 1 0 3948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8256
timestamp 1680363874
transform 1 0 4060 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7540
timestamp 1680363874
transform 1 0 4068 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7461
timestamp 1680363874
transform 1 0 4084 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8257
timestamp 1680363874
transform 1 0 4092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8369
timestamp 1680363874
transform 1 0 4076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8370
timestamp 1680363874
transform 1 0 4084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8371
timestamp 1680363874
transform 1 0 4100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8372
timestamp 1680363874
transform 1 0 4108 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7563
timestamp 1680363874
transform 1 0 4060 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8258
timestamp 1680363874
transform 1 0 4124 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7515
timestamp 1680363874
transform 1 0 4132 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7516
timestamp 1680363874
transform 1 0 4172 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8259
timestamp 1680363874
transform 1 0 4188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8373
timestamp 1680363874
transform 1 0 4212 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7433
timestamp 1680363874
transform 1 0 4228 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8260
timestamp 1680363874
transform 1 0 4228 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7588
timestamp 1680363874
transform 1 0 4220 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8374
timestamp 1680363874
transform 1 0 4252 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7497
timestamp 1680363874
transform 1 0 4284 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8261
timestamp 1680363874
transform 1 0 4268 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7517
timestamp 1680363874
transform 1 0 4276 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8262
timestamp 1680363874
transform 1 0 4284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8263
timestamp 1680363874
transform 1 0 4300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8375
timestamp 1680363874
transform 1 0 4292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7589
timestamp 1680363874
transform 1 0 4300 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8264
timestamp 1680363874
transform 1 0 4316 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7434
timestamp 1680363874
transform 1 0 4332 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7498
timestamp 1680363874
transform 1 0 4332 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8376
timestamp 1680363874
transform 1 0 4332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7499
timestamp 1680363874
transform 1 0 4420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7500
timestamp 1680363874
transform 1 0 4460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7435
timestamp 1680363874
transform 1 0 4476 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8265
timestamp 1680363874
transform 1 0 4420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8266
timestamp 1680363874
transform 1 0 4452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8267
timestamp 1680363874
transform 1 0 4460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8268
timestamp 1680363874
transform 1 0 4468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8269
timestamp 1680363874
transform 1 0 4476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8377
timestamp 1680363874
transform 1 0 4372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7564
timestamp 1680363874
transform 1 0 4388 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7565
timestamp 1680363874
transform 1 0 4412 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7566
timestamp 1680363874
transform 1 0 4452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7518
timestamp 1680363874
transform 1 0 4500 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8270
timestamp 1680363874
transform 1 0 4508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8271
timestamp 1680363874
transform 1 0 4524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8378
timestamp 1680363874
transform 1 0 4492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8379
timestamp 1680363874
transform 1 0 4500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8380
timestamp 1680363874
transform 1 0 4516 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7567
timestamp 1680363874
transform 1 0 4516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7519
timestamp 1680363874
transform 1 0 4532 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8272
timestamp 1680363874
transform 1 0 4564 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7520
timestamp 1680363874
transform 1 0 4572 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8273
timestamp 1680363874
transform 1 0 4588 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7521
timestamp 1680363874
transform 1 0 4604 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8381
timestamp 1680363874
transform 1 0 4580 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7541
timestamp 1680363874
transform 1 0 4596 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8382
timestamp 1680363874
transform 1 0 4604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8383
timestamp 1680363874
transform 1 0 4612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7568
timestamp 1680363874
transform 1 0 4612 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7501
timestamp 1680363874
transform 1 0 4628 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7462
timestamp 1680363874
transform 1 0 4668 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7502
timestamp 1680363874
transform 1 0 4668 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8274
timestamp 1680363874
transform 1 0 4628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8275
timestamp 1680363874
transform 1 0 4636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8276
timestamp 1680363874
transform 1 0 4652 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7522
timestamp 1680363874
transform 1 0 4660 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8277
timestamp 1680363874
transform 1 0 4668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8384
timestamp 1680363874
transform 1 0 4628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7542
timestamp 1680363874
transform 1 0 4636 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7463
timestamp 1680363874
transform 1 0 4692 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8385
timestamp 1680363874
transform 1 0 4644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8386
timestamp 1680363874
transform 1 0 4660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8387
timestamp 1680363874
transform 1 0 4668 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7569
timestamp 1680363874
transform 1 0 4628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7543
timestamp 1680363874
transform 1 0 4676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7503
timestamp 1680363874
transform 1 0 4700 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7504
timestamp 1680363874
transform 1 0 4740 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8278
timestamp 1680363874
transform 1 0 4700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8279
timestamp 1680363874
transform 1 0 4708 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7523
timestamp 1680363874
transform 1 0 4716 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8280
timestamp 1680363874
transform 1 0 4740 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7544
timestamp 1680363874
transform 1 0 4716 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8388
timestamp 1680363874
transform 1 0 4788 0 1 805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_78
timestamp 1680363874
transform 1 0 48 0 1 770
box -10 -3 10 3
use FILL  FILL_9402
timestamp 1680363874
transform 1 0 72 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_506
timestamp 1680363874
transform -1 0 176 0 1 770
box -8 -3 104 105
use FILL  FILL_9403
timestamp 1680363874
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_9406
timestamp 1680363874
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_9407
timestamp 1680363874
transform 1 0 192 0 1 770
box -8 -3 16 105
use FILL  FILL_9408
timestamp 1680363874
transform 1 0 200 0 1 770
box -8 -3 16 105
use FILL  FILL_9409
timestamp 1680363874
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_9410
timestamp 1680363874
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_9411
timestamp 1680363874
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_9412
timestamp 1680363874
transform 1 0 232 0 1 770
box -8 -3 16 105
use FILL  FILL_9413
timestamp 1680363874
transform 1 0 240 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_59
timestamp 1680363874
transform 1 0 248 0 1 770
box -8 -3 32 105
use FILL  FILL_9414
timestamp 1680363874
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_9415
timestamp 1680363874
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_9417
timestamp 1680363874
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_9418
timestamp 1680363874
transform 1 0 296 0 1 770
box -8 -3 16 105
use FILL  FILL_9419
timestamp 1680363874
transform 1 0 304 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7590
timestamp 1680363874
transform 1 0 340 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_60
timestamp 1680363874
transform 1 0 312 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_7591
timestamp 1680363874
transform 1 0 364 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_107
timestamp 1680363874
transform 1 0 336 0 1 770
box -8 -3 32 105
use FILL  FILL_9420
timestamp 1680363874
transform 1 0 360 0 1 770
box -8 -3 16 105
use FILL  FILL_9421
timestamp 1680363874
transform 1 0 368 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_108
timestamp 1680363874
transform 1 0 376 0 1 770
box -8 -3 32 105
use BUFX2  BUFX2_91
timestamp 1680363874
transform -1 0 424 0 1 770
box -5 -3 28 105
use FILL  FILL_9422
timestamp 1680363874
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_9423
timestamp 1680363874
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_9424
timestamp 1680363874
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_9425
timestamp 1680363874
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_9426
timestamp 1680363874
transform 1 0 456 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_509
timestamp 1680363874
transform -1 0 560 0 1 770
box -8 -3 104 105
use FILL  FILL_9427
timestamp 1680363874
transform 1 0 560 0 1 770
box -8 -3 16 105
use FILL  FILL_9428
timestamp 1680363874
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_9429
timestamp 1680363874
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_9430
timestamp 1680363874
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_9431
timestamp 1680363874
transform 1 0 592 0 1 770
box -8 -3 16 105
use FILL  FILL_9432
timestamp 1680363874
transform 1 0 600 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7592
timestamp 1680363874
transform 1 0 620 0 1 775
box -3 -3 3 3
use FILL  FILL_9433
timestamp 1680363874
transform 1 0 608 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7593
timestamp 1680363874
transform 1 0 684 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_510
timestamp 1680363874
transform -1 0 712 0 1 770
box -8 -3 104 105
use FILL  FILL_9434
timestamp 1680363874
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_9435
timestamp 1680363874
transform 1 0 720 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_360
timestamp 1680363874
transform 1 0 728 0 1 770
box -8 -3 46 105
use FILL  FILL_9436
timestamp 1680363874
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_9437
timestamp 1680363874
transform 1 0 776 0 1 770
box -8 -3 16 105
use FILL  FILL_9438
timestamp 1680363874
transform 1 0 784 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_319
timestamp 1680363874
transform 1 0 792 0 1 770
box -8 -3 46 105
use INVX2  INVX2_570
timestamp 1680363874
transform 1 0 832 0 1 770
box -9 -3 26 105
use FILL  FILL_9439
timestamp 1680363874
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_9440
timestamp 1680363874
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_9441
timestamp 1680363874
transform 1 0 864 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_68
timestamp 1680363874
transform 1 0 872 0 1 770
box -8 -3 40 105
use FILL  FILL_9460
timestamp 1680363874
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_9461
timestamp 1680363874
transform 1 0 912 0 1 770
box -8 -3 16 105
use FILL  FILL_9462
timestamp 1680363874
transform 1 0 920 0 1 770
box -8 -3 16 105
use FILL  FILL_9463
timestamp 1680363874
transform 1 0 928 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_362
timestamp 1680363874
transform 1 0 936 0 1 770
box -8 -3 46 105
use FILL  FILL_9464
timestamp 1680363874
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_9465
timestamp 1680363874
transform 1 0 984 0 1 770
box -8 -3 16 105
use INVX2  INVX2_573
timestamp 1680363874
transform -1 0 1008 0 1 770
box -9 -3 26 105
use FILL  FILL_9466
timestamp 1680363874
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_9475
timestamp 1680363874
transform 1 0 1016 0 1 770
box -8 -3 16 105
use FILL  FILL_9477
timestamp 1680363874
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_9479
timestamp 1680363874
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_9481
timestamp 1680363874
transform 1 0 1040 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_363
timestamp 1680363874
transform 1 0 1048 0 1 770
box -8 -3 46 105
use FILL  FILL_9482
timestamp 1680363874
transform 1 0 1088 0 1 770
box -8 -3 16 105
use FILL  FILL_9483
timestamp 1680363874
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_9484
timestamp 1680363874
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_9485
timestamp 1680363874
transform 1 0 1112 0 1 770
box -8 -3 16 105
use FILL  FILL_9486
timestamp 1680363874
transform 1 0 1120 0 1 770
box -8 -3 16 105
use FILL  FILL_9487
timestamp 1680363874
transform 1 0 1128 0 1 770
box -8 -3 16 105
use INVX2  INVX2_574
timestamp 1680363874
transform -1 0 1152 0 1 770
box -9 -3 26 105
use FILL  FILL_9488
timestamp 1680363874
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_9489
timestamp 1680363874
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_9490
timestamp 1680363874
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_9496
timestamp 1680363874
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_9498
timestamp 1680363874
transform 1 0 1184 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_92
timestamp 1680363874
transform -1 0 1216 0 1 770
box -5 -3 28 105
use FILL  FILL_9500
timestamp 1680363874
transform 1 0 1216 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7594
timestamp 1680363874
transform 1 0 1244 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_7595
timestamp 1680363874
transform 1 0 1268 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_514
timestamp 1680363874
transform 1 0 1224 0 1 770
box -8 -3 104 105
use FILL  FILL_9502
timestamp 1680363874
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_9503
timestamp 1680363874
transform 1 0 1328 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_515
timestamp 1680363874
transform 1 0 1336 0 1 770
box -8 -3 104 105
use INVX2  INVX2_577
timestamp 1680363874
transform 1 0 1432 0 1 770
box -9 -3 26 105
use FILL  FILL_9511
timestamp 1680363874
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_9515
timestamp 1680363874
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_9517
timestamp 1680363874
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_9519
timestamp 1680363874
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_9521
timestamp 1680363874
transform 1 0 1480 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_366
timestamp 1680363874
transform 1 0 1488 0 1 770
box -8 -3 46 105
use FILL  FILL_9523
timestamp 1680363874
transform 1 0 1528 0 1 770
box -8 -3 16 105
use FILL  FILL_9530
timestamp 1680363874
transform 1 0 1536 0 1 770
box -8 -3 16 105
use FILL  FILL_9532
timestamp 1680363874
transform 1 0 1544 0 1 770
box -8 -3 16 105
use FILL  FILL_9534
timestamp 1680363874
transform 1 0 1552 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7596
timestamp 1680363874
transform 1 0 1660 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_517
timestamp 1680363874
transform 1 0 1560 0 1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_367
timestamp 1680363874
transform 1 0 1656 0 1 770
box -8 -3 46 105
use FILL  FILL_9535
timestamp 1680363874
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_9546
timestamp 1680363874
transform 1 0 1704 0 1 770
box -8 -3 16 105
use FILL  FILL_9548
timestamp 1680363874
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_9549
timestamp 1680363874
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_9550
timestamp 1680363874
transform 1 0 1728 0 1 770
box -8 -3 16 105
use INVX2  INVX2_578
timestamp 1680363874
transform 1 0 1736 0 1 770
box -9 -3 26 105
use FILL  FILL_9551
timestamp 1680363874
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_9553
timestamp 1680363874
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_9555
timestamp 1680363874
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_9557
timestamp 1680363874
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_9558
timestamp 1680363874
transform 1 0 1784 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1680363874
transform 1 0 1792 0 1 770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_518
timestamp 1680363874
transform -1 0 1920 0 1 770
box -8 -3 104 105
use FILL  FILL_9559
timestamp 1680363874
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_9565
timestamp 1680363874
transform 1 0 1928 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_94
timestamp 1680363874
transform -1 0 1960 0 1 770
box -5 -3 28 105
use BUFX2  BUFX2_95
timestamp 1680363874
transform 1 0 1960 0 1 770
box -5 -3 28 105
use FILL  FILL_9566
timestamp 1680363874
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_9572
timestamp 1680363874
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_9573
timestamp 1680363874
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_9574
timestamp 1680363874
transform 1 0 2008 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_368
timestamp 1680363874
transform 1 0 2016 0 1 770
box -8 -3 46 105
use FILL  FILL_9575
timestamp 1680363874
transform 1 0 2056 0 1 770
box -8 -3 16 105
use FILL  FILL_9576
timestamp 1680363874
transform 1 0 2064 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7597
timestamp 1680363874
transform 1 0 2092 0 1 775
box -3 -3 3 3
use INVX2  INVX2_580
timestamp 1680363874
transform -1 0 2088 0 1 770
box -9 -3 26 105
use FILL  FILL_9577
timestamp 1680363874
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_9579
timestamp 1680363874
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_9580
timestamp 1680363874
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_9581
timestamp 1680363874
transform 1 0 2112 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7598
timestamp 1680363874
transform 1 0 2132 0 1 775
box -3 -3 3 3
use FILL  FILL_9582
timestamp 1680363874
transform 1 0 2120 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_109
timestamp 1680363874
transform 1 0 2128 0 1 770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_521
timestamp 1680363874
transform -1 0 2248 0 1 770
box -8 -3 104 105
use NOR2X1  NOR2X1_110
timestamp 1680363874
transform -1 0 2272 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_159
timestamp 1680363874
transform -1 0 2304 0 1 770
box -8 -3 34 105
use FILL  FILL_9584
timestamp 1680363874
transform 1 0 2304 0 1 770
box -8 -3 16 105
use INVX2  INVX2_581
timestamp 1680363874
transform -1 0 2328 0 1 770
box -9 -3 26 105
use FILL  FILL_9585
timestamp 1680363874
transform 1 0 2328 0 1 770
box -8 -3 16 105
use FILL  FILL_9586
timestamp 1680363874
transform 1 0 2336 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_327
timestamp 1680363874
transform 1 0 2344 0 1 770
box -8 -3 46 105
use FILL  FILL_9587
timestamp 1680363874
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_9588
timestamp 1680363874
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_9589
timestamp 1680363874
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_9590
timestamp 1680363874
transform 1 0 2408 0 1 770
box -8 -3 16 105
use FILL  FILL_9591
timestamp 1680363874
transform 1 0 2416 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_328
timestamp 1680363874
transform -1 0 2464 0 1 770
box -8 -3 46 105
use FILL  FILL_9592
timestamp 1680363874
transform 1 0 2464 0 1 770
box -8 -3 16 105
use FILL  FILL_9606
timestamp 1680363874
transform 1 0 2472 0 1 770
box -8 -3 16 105
use FILL  FILL_9607
timestamp 1680363874
transform 1 0 2480 0 1 770
box -8 -3 16 105
use FILL  FILL_9608
timestamp 1680363874
transform 1 0 2488 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_111
timestamp 1680363874
transform 1 0 2496 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_164
timestamp 1680363874
transform -1 0 2552 0 1 770
box -8 -3 34 105
use FILL  FILL_9609
timestamp 1680363874
transform 1 0 2552 0 1 770
box -8 -3 16 105
use FILL  FILL_9610
timestamp 1680363874
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_9616
timestamp 1680363874
transform 1 0 2568 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_165
timestamp 1680363874
transform -1 0 2608 0 1 770
box -8 -3 34 105
use FILL  FILL_9617
timestamp 1680363874
transform 1 0 2608 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_523
timestamp 1680363874
transform 1 0 2616 0 1 770
box -8 -3 104 105
use FILL  FILL_9618
timestamp 1680363874
transform 1 0 2712 0 1 770
box -8 -3 16 105
use FILL  FILL_9624
timestamp 1680363874
transform 1 0 2720 0 1 770
box -8 -3 16 105
use FILL  FILL_9626
timestamp 1680363874
transform 1 0 2728 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_525
timestamp 1680363874
transform 1 0 2736 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_7599
timestamp 1680363874
transform 1 0 2844 0 1 775
box -3 -3 3 3
use FILL  FILL_9628
timestamp 1680363874
transform 1 0 2832 0 1 770
box -8 -3 16 105
use INVX2  INVX2_586
timestamp 1680363874
transform -1 0 2856 0 1 770
box -9 -3 26 105
use FILL  FILL_9629
timestamp 1680363874
transform 1 0 2856 0 1 770
box -8 -3 16 105
use FILL  FILL_9630
timestamp 1680363874
transform 1 0 2864 0 1 770
box -8 -3 16 105
use FILL  FILL_9638
timestamp 1680363874
transform 1 0 2872 0 1 770
box -8 -3 16 105
use FILL  FILL_9640
timestamp 1680363874
transform 1 0 2880 0 1 770
box -8 -3 16 105
use FILL  FILL_9642
timestamp 1680363874
transform 1 0 2888 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_329
timestamp 1680363874
transform 1 0 2896 0 1 770
box -8 -3 46 105
use FILL  FILL_9644
timestamp 1680363874
transform 1 0 2936 0 1 770
box -8 -3 16 105
use FILL  FILL_9646
timestamp 1680363874
transform 1 0 2944 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7600
timestamp 1680363874
transform 1 0 2964 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_331
timestamp 1680363874
transform 1 0 2952 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_526
timestamp 1680363874
transform -1 0 3088 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_7601
timestamp 1680363874
transform 1 0 3132 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_371
timestamp 1680363874
transform 1 0 3088 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_332
timestamp 1680363874
transform 1 0 3128 0 1 770
box -8 -3 46 105
use FILL  FILL_9648
timestamp 1680363874
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_9649
timestamp 1680363874
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_9650
timestamp 1680363874
transform 1 0 3184 0 1 770
box -8 -3 16 105
use FILL  FILL_9651
timestamp 1680363874
transform 1 0 3192 0 1 770
box -8 -3 16 105
use FILL  FILL_9652
timestamp 1680363874
transform 1 0 3200 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7602
timestamp 1680363874
transform 1 0 3220 0 1 775
box -3 -3 3 3
use INVX2  INVX2_587
timestamp 1680363874
transform 1 0 3208 0 1 770
box -9 -3 26 105
use FILL  FILL_9653
timestamp 1680363874
transform 1 0 3224 0 1 770
box -8 -3 16 105
use FILL  FILL_9654
timestamp 1680363874
transform 1 0 3232 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_333
timestamp 1680363874
transform 1 0 3240 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_527
timestamp 1680363874
transform -1 0 3376 0 1 770
box -8 -3 104 105
use BUFX2  BUFX2_98
timestamp 1680363874
transform 1 0 3376 0 1 770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_528
timestamp 1680363874
transform -1 0 3496 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_7603
timestamp 1680363874
transform 1 0 3524 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_334
timestamp 1680363874
transform -1 0 3536 0 1 770
box -8 -3 46 105
use FILL  FILL_9655
timestamp 1680363874
transform 1 0 3536 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7604
timestamp 1680363874
transform 1 0 3556 0 1 775
box -3 -3 3 3
use FILL  FILL_9666
timestamp 1680363874
transform 1 0 3544 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_336
timestamp 1680363874
transform -1 0 3592 0 1 770
box -8 -3 46 105
use FILL  FILL_9667
timestamp 1680363874
transform 1 0 3592 0 1 770
box -8 -3 16 105
use FILL  FILL_9668
timestamp 1680363874
transform 1 0 3600 0 1 770
box -8 -3 16 105
use FILL  FILL_9672
timestamp 1680363874
transform 1 0 3608 0 1 770
box -8 -3 16 105
use FILL  FILL_9674
timestamp 1680363874
transform 1 0 3616 0 1 770
box -8 -3 16 105
use FILL  FILL_9676
timestamp 1680363874
transform 1 0 3624 0 1 770
box -8 -3 16 105
use FILL  FILL_9678
timestamp 1680363874
transform 1 0 3632 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_338
timestamp 1680363874
transform 1 0 3640 0 1 770
box -8 -3 46 105
use FILL  FILL_9680
timestamp 1680363874
transform 1 0 3680 0 1 770
box -8 -3 16 105
use FILL  FILL_9685
timestamp 1680363874
transform 1 0 3688 0 1 770
box -8 -3 16 105
use FILL  FILL_9687
timestamp 1680363874
transform 1 0 3696 0 1 770
box -8 -3 16 105
use FILL  FILL_9689
timestamp 1680363874
transform 1 0 3704 0 1 770
box -8 -3 16 105
use FILL  FILL_9691
timestamp 1680363874
transform 1 0 3712 0 1 770
box -8 -3 16 105
use FILL  FILL_9692
timestamp 1680363874
transform 1 0 3720 0 1 770
box -8 -3 16 105
use FILL  FILL_9693
timestamp 1680363874
transform 1 0 3728 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7605
timestamp 1680363874
transform 1 0 3748 0 1 775
box -3 -3 3 3
use FILL  FILL_9694
timestamp 1680363874
transform 1 0 3736 0 1 770
box -8 -3 16 105
use FILL  FILL_9695
timestamp 1680363874
transform 1 0 3744 0 1 770
box -8 -3 16 105
use FILL  FILL_9696
timestamp 1680363874
transform 1 0 3752 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_339
timestamp 1680363874
transform 1 0 3760 0 1 770
box -8 -3 46 105
use FILL  FILL_9697
timestamp 1680363874
transform 1 0 3800 0 1 770
box -8 -3 16 105
use FILL  FILL_9698
timestamp 1680363874
transform 1 0 3808 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7606
timestamp 1680363874
transform 1 0 3828 0 1 775
box -3 -3 3 3
use FILL  FILL_9699
timestamp 1680363874
transform 1 0 3816 0 1 770
box -8 -3 16 105
use FILL  FILL_9700
timestamp 1680363874
transform 1 0 3824 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_340
timestamp 1680363874
transform 1 0 3832 0 1 770
box -8 -3 46 105
use FILL  FILL_9702
timestamp 1680363874
transform 1 0 3872 0 1 770
box -8 -3 16 105
use FILL  FILL_9703
timestamp 1680363874
transform 1 0 3880 0 1 770
box -8 -3 16 105
use FILL  FILL_9704
timestamp 1680363874
transform 1 0 3888 0 1 770
box -8 -3 16 105
use FILL  FILL_9705
timestamp 1680363874
transform 1 0 3896 0 1 770
box -8 -3 16 105
use INVX2  INVX2_595
timestamp 1680363874
transform 1 0 3904 0 1 770
box -9 -3 26 105
use FILL  FILL_9706
timestamp 1680363874
transform 1 0 3920 0 1 770
box -8 -3 16 105
use FILL  FILL_9707
timestamp 1680363874
transform 1 0 3928 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_534
timestamp 1680363874
transform 1 0 3936 0 1 770
box -8 -3 104 105
use FILL  FILL_9709
timestamp 1680363874
transform 1 0 4032 0 1 770
box -8 -3 16 105
use FILL  FILL_9711
timestamp 1680363874
transform 1 0 4040 0 1 770
box -8 -3 16 105
use INVX2  INVX2_596
timestamp 1680363874
transform -1 0 4064 0 1 770
box -9 -3 26 105
use FILL  FILL_9713
timestamp 1680363874
transform 1 0 4064 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7607
timestamp 1680363874
transform 1 0 4100 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_341
timestamp 1680363874
transform -1 0 4112 0 1 770
box -8 -3 46 105
use FILL  FILL_9715
timestamp 1680363874
transform 1 0 4112 0 1 770
box -8 -3 16 105
use FILL  FILL_9717
timestamp 1680363874
transform 1 0 4120 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_536
timestamp 1680363874
transform -1 0 4224 0 1 770
box -8 -3 104 105
use FILL  FILL_9718
timestamp 1680363874
transform 1 0 4224 0 1 770
box -8 -3 16 105
use FILL  FILL_9719
timestamp 1680363874
transform 1 0 4232 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7608
timestamp 1680363874
transform 1 0 4252 0 1 775
box -3 -3 3 3
use FILL  FILL_9720
timestamp 1680363874
transform 1 0 4240 0 1 770
box -8 -3 16 105
use FILL  FILL_9721
timestamp 1680363874
transform 1 0 4248 0 1 770
box -8 -3 16 105
use FILL  FILL_9722
timestamp 1680363874
transform 1 0 4256 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_343
timestamp 1680363874
transform 1 0 4264 0 1 770
box -8 -3 46 105
use FILL  FILL_9723
timestamp 1680363874
transform 1 0 4304 0 1 770
box -8 -3 16 105
use FILL  FILL_9724
timestamp 1680363874
transform 1 0 4312 0 1 770
box -8 -3 16 105
use INVX2  INVX2_598
timestamp 1680363874
transform -1 0 4336 0 1 770
box -9 -3 26 105
use FILL  FILL_9725
timestamp 1680363874
transform 1 0 4336 0 1 770
box -8 -3 16 105
use FILL  FILL_9737
timestamp 1680363874
transform 1 0 4344 0 1 770
box -8 -3 16 105
use FILL  FILL_9739
timestamp 1680363874
transform 1 0 4352 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7609
timestamp 1680363874
transform 1 0 4380 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_537
timestamp 1680363874
transform 1 0 4360 0 1 770
box -8 -3 104 105
use INVX2  INVX2_600
timestamp 1680363874
transform -1 0 4472 0 1 770
box -9 -3 26 105
use FILL  FILL_9741
timestamp 1680363874
transform 1 0 4472 0 1 770
box -8 -3 16 105
use FILL  FILL_9742
timestamp 1680363874
transform 1 0 4480 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_347
timestamp 1680363874
transform 1 0 4488 0 1 770
box -8 -3 46 105
use FILL  FILL_9743
timestamp 1680363874
transform 1 0 4528 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7610
timestamp 1680363874
transform 1 0 4548 0 1 775
box -3 -3 3 3
use FILL  FILL_9754
timestamp 1680363874
transform 1 0 4536 0 1 770
box -8 -3 16 105
use FILL  FILL_9756
timestamp 1680363874
transform 1 0 4544 0 1 770
box -8 -3 16 105
use FILL  FILL_9758
timestamp 1680363874
transform 1 0 4552 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_375
timestamp 1680363874
transform 1 0 4560 0 1 770
box -8 -3 46 105
use FILL  FILL_9759
timestamp 1680363874
transform 1 0 4600 0 1 770
box -8 -3 16 105
use INVX2  INVX2_602
timestamp 1680363874
transform 1 0 4608 0 1 770
box -9 -3 26 105
use FILL  FILL_9760
timestamp 1680363874
transform 1 0 4624 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_349
timestamp 1680363874
transform 1 0 4632 0 1 770
box -8 -3 46 105
use FILL  FILL_9761
timestamp 1680363874
transform 1 0 4672 0 1 770
box -8 -3 16 105
use INVX2  INVX2_603
timestamp 1680363874
transform 1 0 4680 0 1 770
box -9 -3 26 105
use FILL  FILL_9762
timestamp 1680363874
transform 1 0 4696 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_538
timestamp 1680363874
transform -1 0 4800 0 1 770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_79
timestamp 1680363874
transform 1 0 4827 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_7666
timestamp 1680363874
transform 1 0 92 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7667
timestamp 1680363874
transform 1 0 164 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8393
timestamp 1680363874
transform 1 0 92 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7720
timestamp 1680363874
transform 1 0 92 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8510
timestamp 1680363874
transform 1 0 116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7721
timestamp 1680363874
transform 1 0 124 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8511
timestamp 1680363874
transform 1 0 172 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7668
timestamp 1680363874
transform 1 0 196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8394
timestamp 1680363874
transform 1 0 196 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7697
timestamp 1680363874
transform 1 0 236 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7698
timestamp 1680363874
transform 1 0 268 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8512
timestamp 1680363874
transform 1 0 236 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8513
timestamp 1680363874
transform 1 0 276 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7611
timestamp 1680363874
transform 1 0 340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7612
timestamp 1680363874
transform 1 0 356 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7669
timestamp 1680363874
transform 1 0 300 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8395
timestamp 1680363874
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8514
timestamp 1680363874
transform 1 0 340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7670
timestamp 1680363874
transform 1 0 476 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8396
timestamp 1680363874
transform 1 0 476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8515
timestamp 1680363874
transform 1 0 388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8516
timestamp 1680363874
transform 1 0 396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8517
timestamp 1680363874
transform 1 0 452 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7671
timestamp 1680363874
transform 1 0 556 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8397
timestamp 1680363874
transform 1 0 508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8518
timestamp 1680363874
transform 1 0 556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8398
timestamp 1680363874
transform 1 0 628 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7633
timestamp 1680363874
transform 1 0 676 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7672
timestamp 1680363874
transform 1 0 660 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8399
timestamp 1680363874
transform 1 0 660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8400
timestamp 1680363874
transform 1 0 676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8401
timestamp 1680363874
transform 1 0 684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8519
timestamp 1680363874
transform 1 0 636 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7722
timestamp 1680363874
transform 1 0 644 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8520
timestamp 1680363874
transform 1 0 652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8521
timestamp 1680363874
transform 1 0 668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8522
timestamp 1680363874
transform 1 0 684 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7634
timestamp 1680363874
transform 1 0 700 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7673
timestamp 1680363874
transform 1 0 748 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8402
timestamp 1680363874
transform 1 0 740 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7674
timestamp 1680363874
transform 1 0 780 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8403
timestamp 1680363874
transform 1 0 780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8404
timestamp 1680363874
transform 1 0 796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8523
timestamp 1680363874
transform 1 0 748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8524
timestamp 1680363874
transform 1 0 756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8525
timestamp 1680363874
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8526
timestamp 1680363874
transform 1 0 788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7748
timestamp 1680363874
transform 1 0 756 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7723
timestamp 1680363874
transform 1 0 796 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8527
timestamp 1680363874
transform 1 0 804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7780
timestamp 1680363874
transform 1 0 788 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7749
timestamp 1680363874
transform 1 0 804 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8405
timestamp 1680363874
transform 1 0 852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8528
timestamp 1680363874
transform 1 0 844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8529
timestamp 1680363874
transform 1 0 860 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7781
timestamp 1680363874
transform 1 0 828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7782
timestamp 1680363874
transform 1 0 860 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7635
timestamp 1680363874
transform 1 0 876 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8530
timestamp 1680363874
transform 1 0 876 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7750
timestamp 1680363874
transform 1 0 876 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8406
timestamp 1680363874
transform 1 0 892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8407
timestamp 1680363874
transform 1 0 924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8531
timestamp 1680363874
transform 1 0 916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7724
timestamp 1680363874
transform 1 0 924 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8532
timestamp 1680363874
transform 1 0 932 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7783
timestamp 1680363874
transform 1 0 916 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7675
timestamp 1680363874
transform 1 0 972 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8408
timestamp 1680363874
transform 1 0 972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8409
timestamp 1680363874
transform 1 0 980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8410
timestamp 1680363874
transform 1 0 996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8533
timestamp 1680363874
transform 1 0 988 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7751
timestamp 1680363874
transform 1 0 972 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7752
timestamp 1680363874
transform 1 0 996 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7784
timestamp 1680363874
transform 1 0 996 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8411
timestamp 1680363874
transform 1 0 1020 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7725
timestamp 1680363874
transform 1 0 1020 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8534
timestamp 1680363874
transform 1 0 1028 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7753
timestamp 1680363874
transform 1 0 1028 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8535
timestamp 1680363874
transform 1 0 1036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8412
timestamp 1680363874
transform 1 0 1060 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7699
timestamp 1680363874
transform 1 0 1084 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8413
timestamp 1680363874
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7700
timestamp 1680363874
transform 1 0 1100 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7676
timestamp 1680363874
transform 1 0 1164 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8414
timestamp 1680363874
transform 1 0 1108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8415
timestamp 1680363874
transform 1 0 1124 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8416
timestamp 1680363874
transform 1 0 1132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8417
timestamp 1680363874
transform 1 0 1156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8418
timestamp 1680363874
transform 1 0 1164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8536
timestamp 1680363874
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8537
timestamp 1680363874
transform 1 0 1116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7726
timestamp 1680363874
transform 1 0 1124 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8538
timestamp 1680363874
transform 1 0 1132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8539
timestamp 1680363874
transform 1 0 1148 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7754
timestamp 1680363874
transform 1 0 1132 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7785
timestamp 1680363874
transform 1 0 1100 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7829
timestamp 1680363874
transform 1 0 1132 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8419
timestamp 1680363874
transform 1 0 1196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8540
timestamp 1680363874
transform 1 0 1212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8541
timestamp 1680363874
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7755
timestamp 1680363874
transform 1 0 1212 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7786
timestamp 1680363874
transform 1 0 1204 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7787
timestamp 1680363874
transform 1 0 1220 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7815
timestamp 1680363874
transform 1 0 1212 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7636
timestamp 1680363874
transform 1 0 1236 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8420
timestamp 1680363874
transform 1 0 1244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8421
timestamp 1680363874
transform 1 0 1260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8422
timestamp 1680363874
transform 1 0 1276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8542
timestamp 1680363874
transform 1 0 1268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7830
timestamp 1680363874
transform 1 0 1252 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8543
timestamp 1680363874
transform 1 0 1284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8423
timestamp 1680363874
transform 1 0 1292 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7727
timestamp 1680363874
transform 1 0 1292 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7677
timestamp 1680363874
transform 1 0 1308 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8424
timestamp 1680363874
transform 1 0 1308 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7678
timestamp 1680363874
transform 1 0 1324 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7756
timestamp 1680363874
transform 1 0 1324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7816
timestamp 1680363874
transform 1 0 1316 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7637
timestamp 1680363874
transform 1 0 1364 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8425
timestamp 1680363874
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8544
timestamp 1680363874
transform 1 0 1412 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7757
timestamp 1680363874
transform 1 0 1412 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7788
timestamp 1680363874
transform 1 0 1388 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7758
timestamp 1680363874
transform 1 0 1452 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7789
timestamp 1680363874
transform 1 0 1468 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7728
timestamp 1680363874
transform 1 0 1484 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8545
timestamp 1680363874
transform 1 0 1492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8546
timestamp 1680363874
transform 1 0 1500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8426
timestamp 1680363874
transform 1 0 1516 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7679
timestamp 1680363874
transform 1 0 1564 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8427
timestamp 1680363874
transform 1 0 1588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8547
timestamp 1680363874
transform 1 0 1564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8548
timestamp 1680363874
transform 1 0 1580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7759
timestamp 1680363874
transform 1 0 1580 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8640
timestamp 1680363874
transform 1 0 1612 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7638
timestamp 1680363874
transform 1 0 1628 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7701
timestamp 1680363874
transform 1 0 1636 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8549
timestamp 1680363874
transform 1 0 1636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8550
timestamp 1680363874
transform 1 0 1652 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7760
timestamp 1680363874
transform 1 0 1652 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8647
timestamp 1680363874
transform 1 0 1660 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_7817
timestamp 1680363874
transform 1 0 1660 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7702
timestamp 1680363874
transform 1 0 1676 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8551
timestamp 1680363874
transform 1 0 1676 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7680
timestamp 1680363874
transform 1 0 1724 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7681
timestamp 1680363874
transform 1 0 1748 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8428
timestamp 1680363874
transform 1 0 1716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8429
timestamp 1680363874
transform 1 0 1724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8430
timestamp 1680363874
transform 1 0 1740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8431
timestamp 1680363874
transform 1 0 1748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8552
timestamp 1680363874
transform 1 0 1732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8641
timestamp 1680363874
transform 1 0 1708 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7790
timestamp 1680363874
transform 1 0 1700 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7761
timestamp 1680363874
transform 1 0 1716 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7639
timestamp 1680363874
transform 1 0 1884 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7682
timestamp 1680363874
transform 1 0 1796 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8432
timestamp 1680363874
transform 1 0 1796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8433
timestamp 1680363874
transform 1 0 1884 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8553
timestamp 1680363874
transform 1 0 1788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8554
timestamp 1680363874
transform 1 0 1796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8555
timestamp 1680363874
transform 1 0 1836 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7831
timestamp 1680363874
transform 1 0 1780 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7762
timestamp 1680363874
transform 1 0 1836 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7818
timestamp 1680363874
transform 1 0 1804 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7832
timestamp 1680363874
transform 1 0 1804 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7640
timestamp 1680363874
transform 1 0 1908 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8556
timestamp 1680363874
transform 1 0 1932 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8434
timestamp 1680363874
transform 1 0 1956 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7613
timestamp 1680363874
transform 1 0 1980 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7614
timestamp 1680363874
transform 1 0 2020 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7641
timestamp 1680363874
transform 1 0 2004 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7642
timestamp 1680363874
transform 1 0 2092 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8435
timestamp 1680363874
transform 1 0 2004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8557
timestamp 1680363874
transform 1 0 2036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8558
timestamp 1680363874
transform 1 0 2084 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7763
timestamp 1680363874
transform 1 0 2036 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7764
timestamp 1680363874
transform 1 0 2052 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8559
timestamp 1680363874
transform 1 0 2100 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7833
timestamp 1680363874
transform 1 0 2100 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8436
timestamp 1680363874
transform 1 0 2116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8437
timestamp 1680363874
transform 1 0 2148 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7703
timestamp 1680363874
transform 1 0 2164 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7643
timestamp 1680363874
transform 1 0 2188 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8438
timestamp 1680363874
transform 1 0 2172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8439
timestamp 1680363874
transform 1 0 2180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8560
timestamp 1680363874
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8642
timestamp 1680363874
transform 1 0 2148 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8440
timestamp 1680363874
transform 1 0 2204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8561
timestamp 1680363874
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8562
timestamp 1680363874
transform 1 0 2204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8643
timestamp 1680363874
transform 1 0 2204 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7791
timestamp 1680363874
transform 1 0 2204 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8441
timestamp 1680363874
transform 1 0 2220 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7644
timestamp 1680363874
transform 1 0 2268 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8644
timestamp 1680363874
transform 1 0 2260 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7792
timestamp 1680363874
transform 1 0 2260 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8442
timestamp 1680363874
transform 1 0 2284 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7704
timestamp 1680363874
transform 1 0 2292 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7729
timestamp 1680363874
transform 1 0 2292 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7615
timestamp 1680363874
transform 1 0 2308 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8563
timestamp 1680363874
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7819
timestamp 1680363874
transform 1 0 2308 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7616
timestamp 1680363874
transform 1 0 2420 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8443
timestamp 1680363874
transform 1 0 2404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8444
timestamp 1680363874
transform 1 0 2428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8445
timestamp 1680363874
transform 1 0 2436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8564
timestamp 1680363874
transform 1 0 2380 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7730
timestamp 1680363874
transform 1 0 2404 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8565
timestamp 1680363874
transform 1 0 2420 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7731
timestamp 1680363874
transform 1 0 2428 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8566
timestamp 1680363874
transform 1 0 2444 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8567
timestamp 1680363874
transform 1 0 2460 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7765
timestamp 1680363874
transform 1 0 2380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7766
timestamp 1680363874
transform 1 0 2420 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7820
timestamp 1680363874
transform 1 0 2372 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8645
timestamp 1680363874
transform 1 0 2460 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8446
timestamp 1680363874
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7617
timestamp 1680363874
transform 1 0 2492 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7732
timestamp 1680363874
transform 1 0 2484 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7793
timestamp 1680363874
transform 1 0 2508 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8447
timestamp 1680363874
transform 1 0 2524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8448
timestamp 1680363874
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8568
timestamp 1680363874
transform 1 0 2532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8569
timestamp 1680363874
transform 1 0 2540 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7767
timestamp 1680363874
transform 1 0 2532 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8646
timestamp 1680363874
transform 1 0 2540 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7794
timestamp 1680363874
transform 1 0 2540 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7768
timestamp 1680363874
transform 1 0 2564 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7834
timestamp 1680363874
transform 1 0 2564 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8449
timestamp 1680363874
transform 1 0 2588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8450
timestamp 1680363874
transform 1 0 2604 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7733
timestamp 1680363874
transform 1 0 2604 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8570
timestamp 1680363874
transform 1 0 2636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8571
timestamp 1680363874
transform 1 0 2700 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7769
timestamp 1680363874
transform 1 0 2604 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7770
timestamp 1680363874
transform 1 0 2692 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7734
timestamp 1680363874
transform 1 0 2708 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7645
timestamp 1680363874
transform 1 0 2764 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8451
timestamp 1680363874
transform 1 0 2748 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7705
timestamp 1680363874
transform 1 0 2756 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8452
timestamp 1680363874
transform 1 0 2764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8572
timestamp 1680363874
transform 1 0 2756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8573
timestamp 1680363874
transform 1 0 2772 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7795
timestamp 1680363874
transform 1 0 2748 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7821
timestamp 1680363874
transform 1 0 2772 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7706
timestamp 1680363874
transform 1 0 2788 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8574
timestamp 1680363874
transform 1 0 2788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8453
timestamp 1680363874
transform 1 0 2820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8454
timestamp 1680363874
transform 1 0 2828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8455
timestamp 1680363874
transform 1 0 2844 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7735
timestamp 1680363874
transform 1 0 2820 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7796
timestamp 1680363874
transform 1 0 2812 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7707
timestamp 1680363874
transform 1 0 2852 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8575
timestamp 1680363874
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7822
timestamp 1680363874
transform 1 0 2844 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7618
timestamp 1680363874
transform 1 0 2868 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8576
timestamp 1680363874
transform 1 0 2868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7646
timestamp 1680363874
transform 1 0 2900 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8456
timestamp 1680363874
transform 1 0 2900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8457
timestamp 1680363874
transform 1 0 2908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8458
timestamp 1680363874
transform 1 0 2924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8577
timestamp 1680363874
transform 1 0 2916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7797
timestamp 1680363874
transform 1 0 2924 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7619
timestamp 1680363874
transform 1 0 2940 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8459
timestamp 1680363874
transform 1 0 2940 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7647
timestamp 1680363874
transform 1 0 2980 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8460
timestamp 1680363874
transform 1 0 2964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8461
timestamp 1680363874
transform 1 0 2980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8462
timestamp 1680363874
transform 1 0 2988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8578
timestamp 1680363874
transform 1 0 2948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8579
timestamp 1680363874
transform 1 0 2956 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8580
timestamp 1680363874
transform 1 0 2972 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7736
timestamp 1680363874
transform 1 0 2980 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8581
timestamp 1680363874
transform 1 0 2996 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7620
timestamp 1680363874
transform 1 0 3012 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7708
timestamp 1680363874
transform 1 0 3004 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7709
timestamp 1680363874
transform 1 0 3020 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7621
timestamp 1680363874
transform 1 0 3116 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7622
timestamp 1680363874
transform 1 0 3156 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7623
timestamp 1680363874
transform 1 0 3204 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7648
timestamp 1680363874
transform 1 0 3036 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7649
timestamp 1680363874
transform 1 0 3108 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7710
timestamp 1680363874
transform 1 0 3060 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8463
timestamp 1680363874
transform 1 0 3108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8582
timestamp 1680363874
transform 1 0 3020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8583
timestamp 1680363874
transform 1 0 3028 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7737
timestamp 1680363874
transform 1 0 3036 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8584
timestamp 1680363874
transform 1 0 3060 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7650
timestamp 1680363874
transform 1 0 3196 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7624
timestamp 1680363874
transform 1 0 3252 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7625
timestamp 1680363874
transform 1 0 3308 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7626
timestamp 1680363874
transform 1 0 3332 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7651
timestamp 1680363874
transform 1 0 3228 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7652
timestamp 1680363874
transform 1 0 3244 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8464
timestamp 1680363874
transform 1 0 3132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8465
timestamp 1680363874
transform 1 0 3220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8466
timestamp 1680363874
transform 1 0 3244 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7711
timestamp 1680363874
transform 1 0 3268 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8467
timestamp 1680363874
transform 1 0 3332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8585
timestamp 1680363874
transform 1 0 3164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8586
timestamp 1680363874
transform 1 0 3220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8587
timestamp 1680363874
transform 1 0 3228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8588
timestamp 1680363874
transform 1 0 3268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8589
timestamp 1680363874
transform 1 0 3324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8590
timestamp 1680363874
transform 1 0 3332 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7835
timestamp 1680363874
transform 1 0 3140 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7836
timestamp 1680363874
transform 1 0 3180 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7798
timestamp 1680363874
transform 1 0 3276 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7799
timestamp 1680363874
transform 1 0 3332 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7837
timestamp 1680363874
transform 1 0 3300 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7838
timestamp 1680363874
transform 1 0 3324 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7712
timestamp 1680363874
transform 1 0 3340 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8468
timestamp 1680363874
transform 1 0 3348 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7653
timestamp 1680363874
transform 1 0 3364 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8591
timestamp 1680363874
transform 1 0 3356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8592
timestamp 1680363874
transform 1 0 3380 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7823
timestamp 1680363874
transform 1 0 3380 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7627
timestamp 1680363874
transform 1 0 3404 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7654
timestamp 1680363874
transform 1 0 3396 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7683
timestamp 1680363874
transform 1 0 3412 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8469
timestamp 1680363874
transform 1 0 3396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8470
timestamp 1680363874
transform 1 0 3404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8471
timestamp 1680363874
transform 1 0 3420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8593
timestamp 1680363874
transform 1 0 3412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8594
timestamp 1680363874
transform 1 0 3428 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7800
timestamp 1680363874
transform 1 0 3428 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8472
timestamp 1680363874
transform 1 0 3452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8595
timestamp 1680363874
transform 1 0 3444 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7738
timestamp 1680363874
transform 1 0 3452 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7655
timestamp 1680363874
transform 1 0 3468 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8596
timestamp 1680363874
transform 1 0 3468 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7801
timestamp 1680363874
transform 1 0 3460 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7684
timestamp 1680363874
transform 1 0 3484 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8473
timestamp 1680363874
transform 1 0 3484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8474
timestamp 1680363874
transform 1 0 3492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8475
timestamp 1680363874
transform 1 0 3508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8597
timestamp 1680363874
transform 1 0 3484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8598
timestamp 1680363874
transform 1 0 3516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7802
timestamp 1680363874
transform 1 0 3516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7628
timestamp 1680363874
transform 1 0 3532 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7656
timestamp 1680363874
transform 1 0 3532 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7657
timestamp 1680363874
transform 1 0 3580 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7685
timestamp 1680363874
transform 1 0 3572 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8476
timestamp 1680363874
transform 1 0 3556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8477
timestamp 1680363874
transform 1 0 3564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8478
timestamp 1680363874
transform 1 0 3572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8479
timestamp 1680363874
transform 1 0 3588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8480
timestamp 1680363874
transform 1 0 3596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8599
timestamp 1680363874
transform 1 0 3564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8600
timestamp 1680363874
transform 1 0 3580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7803
timestamp 1680363874
transform 1 0 3556 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7739
timestamp 1680363874
transform 1 0 3588 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7839
timestamp 1680363874
transform 1 0 3564 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8601
timestamp 1680363874
transform 1 0 3612 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7804
timestamp 1680363874
transform 1 0 3604 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7840
timestamp 1680363874
transform 1 0 3596 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7740
timestamp 1680363874
transform 1 0 3620 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7658
timestamp 1680363874
transform 1 0 3644 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7659
timestamp 1680363874
transform 1 0 3684 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8602
timestamp 1680363874
transform 1 0 3684 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7686
timestamp 1680363874
transform 1 0 3716 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7660
timestamp 1680363874
transform 1 0 3764 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7687
timestamp 1680363874
transform 1 0 3780 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8481
timestamp 1680363874
transform 1 0 3716 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7713
timestamp 1680363874
transform 1 0 3724 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8482
timestamp 1680363874
transform 1 0 3740 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7714
timestamp 1680363874
transform 1 0 3764 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7741
timestamp 1680363874
transform 1 0 3716 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8603
timestamp 1680363874
transform 1 0 3724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8604
timestamp 1680363874
transform 1 0 3764 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7742
timestamp 1680363874
transform 1 0 3812 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8605
timestamp 1680363874
transform 1 0 3820 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7805
timestamp 1680363874
transform 1 0 3740 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7824
timestamp 1680363874
transform 1 0 3732 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7629
timestamp 1680363874
transform 1 0 3844 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8483
timestamp 1680363874
transform 1 0 3844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8606
timestamp 1680363874
transform 1 0 3868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8607
timestamp 1680363874
transform 1 0 3924 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7688
timestamp 1680363874
transform 1 0 3988 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7689
timestamp 1680363874
transform 1 0 4028 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8484
timestamp 1680363874
transform 1 0 3948 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7715
timestamp 1680363874
transform 1 0 4028 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8608
timestamp 1680363874
transform 1 0 3996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8609
timestamp 1680363874
transform 1 0 4028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8610
timestamp 1680363874
transform 1 0 4036 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7771
timestamp 1680363874
transform 1 0 3972 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7772
timestamp 1680363874
transform 1 0 3996 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7806
timestamp 1680363874
transform 1 0 3948 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7773
timestamp 1680363874
transform 1 0 4036 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7807
timestamp 1680363874
transform 1 0 4044 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7661
timestamp 1680363874
transform 1 0 4100 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8485
timestamp 1680363874
transform 1 0 4076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8486
timestamp 1680363874
transform 1 0 4084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8487
timestamp 1680363874
transform 1 0 4100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8611
timestamp 1680363874
transform 1 0 4076 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7743
timestamp 1680363874
transform 1 0 4084 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8612
timestamp 1680363874
transform 1 0 4092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8613
timestamp 1680363874
transform 1 0 4108 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7774
timestamp 1680363874
transform 1 0 4076 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7808
timestamp 1680363874
transform 1 0 4068 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7841
timestamp 1680363874
transform 1 0 4108 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7744
timestamp 1680363874
transform 1 0 4124 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8614
timestamp 1680363874
transform 1 0 4132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7825
timestamp 1680363874
transform 1 0 4132 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7690
timestamp 1680363874
transform 1 0 4148 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8488
timestamp 1680363874
transform 1 0 4148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8489
timestamp 1680363874
transform 1 0 4164 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7716
timestamp 1680363874
transform 1 0 4172 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8615
timestamp 1680363874
transform 1 0 4156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8616
timestamp 1680363874
transform 1 0 4172 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7775
timestamp 1680363874
transform 1 0 4172 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8617
timestamp 1680363874
transform 1 0 4188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7809
timestamp 1680363874
transform 1 0 4180 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7691
timestamp 1680363874
transform 1 0 4260 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8490
timestamp 1680363874
transform 1 0 4228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8491
timestamp 1680363874
transform 1 0 4236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8492
timestamp 1680363874
transform 1 0 4252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8493
timestamp 1680363874
transform 1 0 4260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8618
timestamp 1680363874
transform 1 0 4220 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7745
timestamp 1680363874
transform 1 0 4236 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8619
timestamp 1680363874
transform 1 0 4244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8620
timestamp 1680363874
transform 1 0 4260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8621
timestamp 1680363874
transform 1 0 4268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7810
timestamp 1680363874
transform 1 0 4228 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7826
timestamp 1680363874
transform 1 0 4260 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7630
timestamp 1680363874
transform 1 0 4308 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7692
timestamp 1680363874
transform 1 0 4292 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7717
timestamp 1680363874
transform 1 0 4324 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8494
timestamp 1680363874
transform 1 0 4332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8622
timestamp 1680363874
transform 1 0 4308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8623
timestamp 1680363874
transform 1 0 4324 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7662
timestamp 1680363874
transform 1 0 4340 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8624
timestamp 1680363874
transform 1 0 4340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7631
timestamp 1680363874
transform 1 0 4372 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7663
timestamp 1680363874
transform 1 0 4372 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7693
timestamp 1680363874
transform 1 0 4404 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8495
timestamp 1680363874
transform 1 0 4388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8496
timestamp 1680363874
transform 1 0 4404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8625
timestamp 1680363874
transform 1 0 4380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8626
timestamp 1680363874
transform 1 0 4396 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7632
timestamp 1680363874
transform 1 0 4428 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7746
timestamp 1680363874
transform 1 0 4436 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8627
timestamp 1680363874
transform 1 0 4460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8497
timestamp 1680363874
transform 1 0 4484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8498
timestamp 1680363874
transform 1 0 4492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8499
timestamp 1680363874
transform 1 0 4508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8628
timestamp 1680363874
transform 1 0 4476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7747
timestamp 1680363874
transform 1 0 4492 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8629
timestamp 1680363874
transform 1 0 4500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8630
timestamp 1680363874
transform 1 0 4516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7827
timestamp 1680363874
transform 1 0 4492 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8500
timestamp 1680363874
transform 1 0 4572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8631
timestamp 1680363874
transform 1 0 4564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8632
timestamp 1680363874
transform 1 0 4580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7776
timestamp 1680363874
transform 1 0 4564 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7811
timestamp 1680363874
transform 1 0 4580 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7694
timestamp 1680363874
transform 1 0 4596 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7664
timestamp 1680363874
transform 1 0 4636 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8501
timestamp 1680363874
transform 1 0 4596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8502
timestamp 1680363874
transform 1 0 4604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8503
timestamp 1680363874
transform 1 0 4620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8633
timestamp 1680363874
transform 1 0 4596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8634
timestamp 1680363874
transform 1 0 4628 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7777
timestamp 1680363874
transform 1 0 4596 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7812
timestamp 1680363874
transform 1 0 4628 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7665
timestamp 1680363874
transform 1 0 4684 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7695
timestamp 1680363874
transform 1 0 4676 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8504
timestamp 1680363874
transform 1 0 4644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8505
timestamp 1680363874
transform 1 0 4652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8506
timestamp 1680363874
transform 1 0 4676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8507
timestamp 1680363874
transform 1 0 4684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8508
timestamp 1680363874
transform 1 0 4692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8635
timestamp 1680363874
transform 1 0 4652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8636
timestamp 1680363874
transform 1 0 4668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7696
timestamp 1680363874
transform 1 0 4708 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7718
timestamp 1680363874
transform 1 0 4700 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7719
timestamp 1680363874
transform 1 0 4740 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8509
timestamp 1680363874
transform 1 0 4788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8637
timestamp 1680363874
transform 1 0 4700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8638
timestamp 1680363874
transform 1 0 4708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8639
timestamp 1680363874
transform 1 0 4740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7778
timestamp 1680363874
transform 1 0 4668 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7779
timestamp 1680363874
transform 1 0 4692 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7813
timestamp 1680363874
transform 1 0 4644 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7814
timestamp 1680363874
transform 1 0 4668 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7828
timestamp 1680363874
transform 1 0 4652 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7842
timestamp 1680363874
transform 1 0 4644 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7843
timestamp 1680363874
transform 1 0 4724 0 1 685
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_80
timestamp 1680363874
transform 1 0 24 0 1 670
box -10 -3 10 3
use FILL  FILL_9404
timestamp 1680363874
transform 1 0 72 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_507
timestamp 1680363874
transform 1 0 80 0 -1 770
box -8 -3 104 105
use FILL  FILL_9405
timestamp 1680363874
transform 1 0 176 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_508
timestamp 1680363874
transform 1 0 184 0 -1 770
box -8 -3 104 105
use FILL  FILL_9416
timestamp 1680363874
transform 1 0 280 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_511
timestamp 1680363874
transform 1 0 288 0 -1 770
box -8 -3 104 105
use FILL  FILL_9442
timestamp 1680363874
transform 1 0 384 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_512
timestamp 1680363874
transform -1 0 488 0 -1 770
box -8 -3 104 105
use FILL  FILL_9443
timestamp 1680363874
transform 1 0 488 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_513
timestamp 1680363874
transform 1 0 496 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_571
timestamp 1680363874
transform 1 0 592 0 -1 770
box -9 -3 26 105
use FILL  FILL_9444
timestamp 1680363874
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9445
timestamp 1680363874
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_9446
timestamp 1680363874
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9447
timestamp 1680363874
transform 1 0 632 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_361
timestamp 1680363874
transform -1 0 680 0 -1 770
box -8 -3 46 105
use FILL  FILL_9448
timestamp 1680363874
transform 1 0 680 0 -1 770
box -8 -3 16 105
use FILL  FILL_9449
timestamp 1680363874
transform 1 0 688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9450
timestamp 1680363874
transform 1 0 696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9451
timestamp 1680363874
transform 1 0 704 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_572
timestamp 1680363874
transform 1 0 712 0 -1 770
box -9 -3 26 105
use FILL  FILL_9452
timestamp 1680363874
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_9453
timestamp 1680363874
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_9454
timestamp 1680363874
transform 1 0 744 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_320
timestamp 1680363874
transform 1 0 752 0 -1 770
box -8 -3 46 105
use FILL  FILL_9455
timestamp 1680363874
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_9456
timestamp 1680363874
transform 1 0 800 0 -1 770
box -8 -3 16 105
use FILL  FILL_9457
timestamp 1680363874
transform 1 0 808 0 -1 770
box -8 -3 16 105
use FILL  FILL_9458
timestamp 1680363874
transform 1 0 816 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_321
timestamp 1680363874
transform 1 0 824 0 -1 770
box -8 -3 46 105
use FILL  FILL_9459
timestamp 1680363874
transform 1 0 864 0 -1 770
box -8 -3 16 105
use FILL  FILL_9467
timestamp 1680363874
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_9468
timestamp 1680363874
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_9469
timestamp 1680363874
transform 1 0 888 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_322
timestamp 1680363874
transform 1 0 896 0 -1 770
box -8 -3 46 105
use FILL  FILL_9470
timestamp 1680363874
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_9471
timestamp 1680363874
transform 1 0 944 0 -1 770
box -8 -3 16 105
use FILL  FILL_9472
timestamp 1680363874
transform 1 0 952 0 -1 770
box -8 -3 16 105
use FILL  FILL_9473
timestamp 1680363874
transform 1 0 960 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_323
timestamp 1680363874
transform -1 0 1008 0 -1 770
box -8 -3 46 105
use FILL  FILL_9474
timestamp 1680363874
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_9476
timestamp 1680363874
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_9478
timestamp 1680363874
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_9480
timestamp 1680363874
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_575
timestamp 1680363874
transform 1 0 1040 0 -1 770
box -9 -3 26 105
use FILL  FILL_9491
timestamp 1680363874
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_9492
timestamp 1680363874
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_9493
timestamp 1680363874
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_9494
timestamp 1680363874
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7844
timestamp 1680363874
transform 1 0 1132 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_364
timestamp 1680363874
transform 1 0 1088 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_324
timestamp 1680363874
transform 1 0 1128 0 -1 770
box -8 -3 46 105
use FILL  FILL_9495
timestamp 1680363874
transform 1 0 1168 0 -1 770
box -8 -3 16 105
use FILL  FILL_9497
timestamp 1680363874
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_9499
timestamp 1680363874
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_93
timestamp 1680363874
transform -1 0 1216 0 -1 770
box -5 -3 28 105
use FILL  FILL_9501
timestamp 1680363874
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7845
timestamp 1680363874
transform 1 0 1236 0 1 675
box -3 -3 3 3
use FILL  FILL_9504
timestamp 1680363874
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_9505
timestamp 1680363874
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_365
timestamp 1680363874
transform 1 0 1240 0 -1 770
box -8 -3 46 105
use FILL  FILL_9506
timestamp 1680363874
transform 1 0 1280 0 -1 770
box -8 -3 16 105
use FILL  FILL_9507
timestamp 1680363874
transform 1 0 1288 0 -1 770
box -8 -3 16 105
use FILL  FILL_9508
timestamp 1680363874
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_9509
timestamp 1680363874
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_576
timestamp 1680363874
transform 1 0 1312 0 -1 770
box -9 -3 26 105
use FILL  FILL_9510
timestamp 1680363874
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_9512
timestamp 1680363874
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_9513
timestamp 1680363874
transform 1 0 1344 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_516
timestamp 1680363874
transform 1 0 1352 0 -1 770
box -8 -3 104 105
use FILL  FILL_9514
timestamp 1680363874
transform 1 0 1448 0 -1 770
box -8 -3 16 105
use FILL  FILL_9516
timestamp 1680363874
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use FILL  FILL_9518
timestamp 1680363874
transform 1 0 1464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9520
timestamp 1680363874
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_9522
timestamp 1680363874
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7846
timestamp 1680363874
transform 1 0 1500 0 1 675
box -3 -3 3 3
use FILL  FILL_9524
timestamp 1680363874
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_9525
timestamp 1680363874
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use FILL  FILL_9526
timestamp 1680363874
transform 1 0 1504 0 -1 770
box -8 -3 16 105
use FILL  FILL_9527
timestamp 1680363874
transform 1 0 1512 0 -1 770
box -8 -3 16 105
use FILL  FILL_9528
timestamp 1680363874
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_9529
timestamp 1680363874
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use FILL  FILL_9531
timestamp 1680363874
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_9533
timestamp 1680363874
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_9536
timestamp 1680363874
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_325
timestamp 1680363874
transform -1 0 1600 0 -1 770
box -8 -3 46 105
use FILL  FILL_9537
timestamp 1680363874
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_9538
timestamp 1680363874
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9539
timestamp 1680363874
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_9540
timestamp 1680363874
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9541
timestamp 1680363874
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1680363874
transform 1 0 1640 0 -1 770
box -8 -3 40 105
use FILL  FILL_9542
timestamp 1680363874
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_9543
timestamp 1680363874
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_9544
timestamp 1680363874
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9545
timestamp 1680363874
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9547
timestamp 1680363874
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_326
timestamp 1680363874
transform 1 0 1712 0 -1 770
box -8 -3 46 105
use M3_M2  M3_M2_7847
timestamp 1680363874
transform 1 0 1764 0 1 675
box -3 -3 3 3
use FILL  FILL_9552
timestamp 1680363874
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_9554
timestamp 1680363874
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7848
timestamp 1680363874
transform 1 0 1780 0 1 675
box -3 -3 3 3
use FILL  FILL_9556
timestamp 1680363874
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_9560
timestamp 1680363874
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_579
timestamp 1680363874
transform -1 0 1800 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_519
timestamp 1680363874
transform -1 0 1896 0 -1 770
box -8 -3 104 105
use FILL  FILL_9561
timestamp 1680363874
transform 1 0 1896 0 -1 770
box -8 -3 16 105
use FILL  FILL_9562
timestamp 1680363874
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use FILL  FILL_9563
timestamp 1680363874
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use FILL  FILL_9564
timestamp 1680363874
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_9567
timestamp 1680363874
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_96
timestamp 1680363874
transform 1 0 1936 0 -1 770
box -5 -3 28 105
use FILL  FILL_9568
timestamp 1680363874
transform 1 0 1960 0 -1 770
box -8 -3 16 105
use FILL  FILL_9569
timestamp 1680363874
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_9570
timestamp 1680363874
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_9571
timestamp 1680363874
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7849
timestamp 1680363874
transform 1 0 2060 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_520
timestamp 1680363874
transform 1 0 1992 0 -1 770
box -8 -3 104 105
use FILL  FILL_9578
timestamp 1680363874
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7850
timestamp 1680363874
transform 1 0 2116 0 1 675
box -3 -3 3 3
use BUFX2  BUFX2_97
timestamp 1680363874
transform 1 0 2096 0 -1 770
box -5 -3 28 105
use FILL  FILL_9583
timestamp 1680363874
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use FILL  FILL_9593
timestamp 1680363874
transform 1 0 2128 0 -1 770
box -8 -3 16 105
use FILL  FILL_9594
timestamp 1680363874
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_160
timestamp 1680363874
transform -1 0 2176 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1680363874
transform 1 0 2176 0 -1 770
box -8 -3 34 105
use FILL  FILL_9595
timestamp 1680363874
transform 1 0 2208 0 -1 770
box -8 -3 16 105
use FILL  FILL_9596
timestamp 1680363874
transform 1 0 2216 0 -1 770
box -8 -3 16 105
use FILL  FILL_9597
timestamp 1680363874
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_162
timestamp 1680363874
transform 1 0 2232 0 -1 770
box -8 -3 34 105
use FILL  FILL_9598
timestamp 1680363874
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_9599
timestamp 1680363874
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_9600
timestamp 1680363874
transform 1 0 2280 0 -1 770
box -8 -3 16 105
use FILL  FILL_9601
timestamp 1680363874
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_9602
timestamp 1680363874
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use FILL  FILL_9603
timestamp 1680363874
transform 1 0 2304 0 -1 770
box -8 -3 16 105
use FILL  FILL_9604
timestamp 1680363874
transform 1 0 2312 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_522
timestamp 1680363874
transform -1 0 2416 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_582
timestamp 1680363874
transform -1 0 2432 0 -1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_163
timestamp 1680363874
transform 1 0 2432 0 -1 770
box -8 -3 34 105
use FILL  FILL_9605
timestamp 1680363874
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9611
timestamp 1680363874
transform 1 0 2472 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_583
timestamp 1680363874
transform -1 0 2496 0 -1 770
box -9 -3 26 105
use FILL  FILL_9612
timestamp 1680363874
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_9613
timestamp 1680363874
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_9614
timestamp 1680363874
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_61
timestamp 1680363874
transform 1 0 2520 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_584
timestamp 1680363874
transform -1 0 2560 0 -1 770
box -9 -3 26 105
use FILL  FILL_9615
timestamp 1680363874
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_9619
timestamp 1680363874
transform 1 0 2568 0 -1 770
box -8 -3 16 105
use FILL  FILL_9620
timestamp 1680363874
transform 1 0 2576 0 -1 770
box -8 -3 16 105
use FILL  FILL_9621
timestamp 1680363874
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_524
timestamp 1680363874
transform 1 0 2592 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_585
timestamp 1680363874
transform 1 0 2688 0 -1 770
box -9 -3 26 105
use FILL  FILL_9622
timestamp 1680363874
transform 1 0 2704 0 -1 770
box -8 -3 16 105
use FILL  FILL_9623
timestamp 1680363874
transform 1 0 2712 0 -1 770
box -8 -3 16 105
use FILL  FILL_9625
timestamp 1680363874
transform 1 0 2720 0 -1 770
box -8 -3 16 105
use FILL  FILL_9627
timestamp 1680363874
transform 1 0 2728 0 -1 770
box -8 -3 16 105
use FILL  FILL_9631
timestamp 1680363874
transform 1 0 2736 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_369
timestamp 1680363874
transform 1 0 2744 0 -1 770
box -8 -3 46 105
use FILL  FILL_9632
timestamp 1680363874
transform 1 0 2784 0 -1 770
box -8 -3 16 105
use FILL  FILL_9633
timestamp 1680363874
transform 1 0 2792 0 -1 770
box -8 -3 16 105
use FILL  FILL_9634
timestamp 1680363874
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use FILL  FILL_9635
timestamp 1680363874
transform 1 0 2808 0 -1 770
box -8 -3 16 105
use FILL  FILL_9636
timestamp 1680363874
transform 1 0 2816 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_370
timestamp 1680363874
transform 1 0 2824 0 -1 770
box -8 -3 46 105
use FILL  FILL_9637
timestamp 1680363874
transform 1 0 2864 0 -1 770
box -8 -3 16 105
use FILL  FILL_9639
timestamp 1680363874
transform 1 0 2872 0 -1 770
box -8 -3 16 105
use FILL  FILL_9641
timestamp 1680363874
transform 1 0 2880 0 -1 770
box -8 -3 16 105
use FILL  FILL_9643
timestamp 1680363874
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_330
timestamp 1680363874
transform 1 0 2896 0 -1 770
box -8 -3 46 105
use FILL  FILL_9645
timestamp 1680363874
transform 1 0 2936 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7851
timestamp 1680363874
transform 1 0 2956 0 1 675
box -3 -3 3 3
use FILL  FILL_9647
timestamp 1680363874
transform 1 0 2944 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_335
timestamp 1680363874
transform 1 0 2952 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_588
timestamp 1680363874
transform 1 0 2992 0 -1 770
box -9 -3 26 105
use FILL  FILL_9656
timestamp 1680363874
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_9657
timestamp 1680363874
transform 1 0 3016 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_529
timestamp 1680363874
transform -1 0 3120 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_530
timestamp 1680363874
transform 1 0 3120 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_589
timestamp 1680363874
transform 1 0 3216 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_531
timestamp 1680363874
transform 1 0 3232 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_590
timestamp 1680363874
transform 1 0 3328 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_591
timestamp 1680363874
transform 1 0 3344 0 -1 770
box -9 -3 26 105
use FILL  FILL_9658
timestamp 1680363874
transform 1 0 3360 0 -1 770
box -8 -3 16 105
use FILL  FILL_9659
timestamp 1680363874
transform 1 0 3368 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_99
timestamp 1680363874
transform 1 0 3376 0 -1 770
box -5 -3 28 105
use OAI22X1  OAI22X1_372
timestamp 1680363874
transform 1 0 3400 0 -1 770
box -8 -3 46 105
use FILL  FILL_9660
timestamp 1680363874
transform 1 0 3440 0 -1 770
box -8 -3 16 105
use FILL  FILL_9661
timestamp 1680363874
transform 1 0 3448 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_592
timestamp 1680363874
transform -1 0 3472 0 -1 770
box -9 -3 26 105
use FILL  FILL_9662
timestamp 1680363874
transform 1 0 3472 0 -1 770
box -8 -3 16 105
use FILL  FILL_9663
timestamp 1680363874
transform 1 0 3480 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_373
timestamp 1680363874
transform 1 0 3488 0 -1 770
box -8 -3 46 105
use FILL  FILL_9664
timestamp 1680363874
transform 1 0 3528 0 -1 770
box -8 -3 16 105
use FILL  FILL_9665
timestamp 1680363874
transform 1 0 3536 0 -1 770
box -8 -3 16 105
use FILL  FILL_9669
timestamp 1680363874
transform 1 0 3544 0 -1 770
box -8 -3 16 105
use FILL  FILL_9670
timestamp 1680363874
transform 1 0 3552 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_337
timestamp 1680363874
transform 1 0 3560 0 -1 770
box -8 -3 46 105
use FILL  FILL_9671
timestamp 1680363874
transform 1 0 3600 0 -1 770
box -8 -3 16 105
use FILL  FILL_9673
timestamp 1680363874
transform 1 0 3608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9675
timestamp 1680363874
transform 1 0 3616 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7852
timestamp 1680363874
transform 1 0 3636 0 1 675
box -3 -3 3 3
use FILL  FILL_9677
timestamp 1680363874
transform 1 0 3624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9679
timestamp 1680363874
transform 1 0 3632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9681
timestamp 1680363874
transform 1 0 3640 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_593
timestamp 1680363874
transform 1 0 3648 0 -1 770
box -9 -3 26 105
use FILL  FILL_9682
timestamp 1680363874
transform 1 0 3664 0 -1 770
box -8 -3 16 105
use FILL  FILL_9683
timestamp 1680363874
transform 1 0 3672 0 -1 770
box -8 -3 16 105
use FILL  FILL_9684
timestamp 1680363874
transform 1 0 3680 0 -1 770
box -8 -3 16 105
use FILL  FILL_9686
timestamp 1680363874
transform 1 0 3688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9688
timestamp 1680363874
transform 1 0 3696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9690
timestamp 1680363874
transform 1 0 3704 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_594
timestamp 1680363874
transform 1 0 3712 0 -1 770
box -9 -3 26 105
use M3_M2  M3_M2_7853
timestamp 1680363874
transform 1 0 3788 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_532
timestamp 1680363874
transform 1 0 3728 0 -1 770
box -8 -3 104 105
use FILL  FILL_9701
timestamp 1680363874
transform 1 0 3824 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_533
timestamp 1680363874
transform 1 0 3832 0 -1 770
box -8 -3 104 105
use FILL  FILL_9708
timestamp 1680363874
transform 1 0 3928 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_535
timestamp 1680363874
transform 1 0 3936 0 -1 770
box -8 -3 104 105
use FILL  FILL_9710
timestamp 1680363874
transform 1 0 4032 0 -1 770
box -8 -3 16 105
use FILL  FILL_9712
timestamp 1680363874
transform 1 0 4040 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_597
timestamp 1680363874
transform -1 0 4064 0 -1 770
box -9 -3 26 105
use FILL  FILL_9714
timestamp 1680363874
transform 1 0 4064 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_342
timestamp 1680363874
transform -1 0 4112 0 -1 770
box -8 -3 46 105
use FILL  FILL_9716
timestamp 1680363874
transform 1 0 4112 0 -1 770
box -8 -3 16 105
use FILL  FILL_9726
timestamp 1680363874
transform 1 0 4120 0 -1 770
box -8 -3 16 105
use FILL  FILL_9727
timestamp 1680363874
transform 1 0 4128 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_344
timestamp 1680363874
transform 1 0 4136 0 -1 770
box -8 -3 46 105
use FILL  FILL_9728
timestamp 1680363874
transform 1 0 4176 0 -1 770
box -8 -3 16 105
use FILL  FILL_9729
timestamp 1680363874
transform 1 0 4184 0 -1 770
box -8 -3 16 105
use FILL  FILL_9730
timestamp 1680363874
transform 1 0 4192 0 -1 770
box -8 -3 16 105
use FILL  FILL_9731
timestamp 1680363874
transform 1 0 4200 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_599
timestamp 1680363874
transform -1 0 4224 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_345
timestamp 1680363874
transform -1 0 4264 0 -1 770
box -8 -3 46 105
use FILL  FILL_9732
timestamp 1680363874
transform 1 0 4264 0 -1 770
box -8 -3 16 105
use FILL  FILL_9733
timestamp 1680363874
transform 1 0 4272 0 -1 770
box -8 -3 16 105
use FILL  FILL_9734
timestamp 1680363874
transform 1 0 4280 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_346
timestamp 1680363874
transform 1 0 4288 0 -1 770
box -8 -3 46 105
use FILL  FILL_9735
timestamp 1680363874
transform 1 0 4328 0 -1 770
box -8 -3 16 105
use FILL  FILL_9736
timestamp 1680363874
transform 1 0 4336 0 -1 770
box -8 -3 16 105
use FILL  FILL_9738
timestamp 1680363874
transform 1 0 4344 0 -1 770
box -8 -3 16 105
use FILL  FILL_9740
timestamp 1680363874
transform 1 0 4352 0 -1 770
box -8 -3 16 105
use FILL  FILL_9744
timestamp 1680363874
transform 1 0 4360 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_374
timestamp 1680363874
transform 1 0 4368 0 -1 770
box -8 -3 46 105
use FILL  FILL_9745
timestamp 1680363874
transform 1 0 4408 0 -1 770
box -8 -3 16 105
use FILL  FILL_9746
timestamp 1680363874
transform 1 0 4416 0 -1 770
box -8 -3 16 105
use FILL  FILL_9747
timestamp 1680363874
transform 1 0 4424 0 -1 770
box -8 -3 16 105
use FILL  FILL_9748
timestamp 1680363874
transform 1 0 4432 0 -1 770
box -8 -3 16 105
use FILL  FILL_9749
timestamp 1680363874
transform 1 0 4440 0 -1 770
box -8 -3 16 105
use FILL  FILL_9750
timestamp 1680363874
transform 1 0 4448 0 -1 770
box -8 -3 16 105
use FILL  FILL_9751
timestamp 1680363874
transform 1 0 4456 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_601
timestamp 1680363874
transform -1 0 4480 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_348
timestamp 1680363874
transform 1 0 4480 0 -1 770
box -8 -3 46 105
use FILL  FILL_9752
timestamp 1680363874
transform 1 0 4520 0 -1 770
box -8 -3 16 105
use FILL  FILL_9753
timestamp 1680363874
transform 1 0 4528 0 -1 770
box -8 -3 16 105
use FILL  FILL_9755
timestamp 1680363874
transform 1 0 4536 0 -1 770
box -8 -3 16 105
use FILL  FILL_9757
timestamp 1680363874
transform 1 0 4544 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_376
timestamp 1680363874
transform 1 0 4552 0 -1 770
box -8 -3 46 105
use FILL  FILL_9763
timestamp 1680363874
transform 1 0 4592 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_377
timestamp 1680363874
transform 1 0 4600 0 -1 770
box -8 -3 46 105
use FILL  FILL_9764
timestamp 1680363874
transform 1 0 4640 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_350
timestamp 1680363874
transform 1 0 4648 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_604
timestamp 1680363874
transform 1 0 4688 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_539
timestamp 1680363874
transform -1 0 4800 0 -1 770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_81
timestamp 1680363874
transform 1 0 4851 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_8661
timestamp 1680363874
transform 1 0 84 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8662
timestamp 1680363874
transform 1 0 92 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8788
timestamp 1680363874
transform 1 0 76 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7942
timestamp 1680363874
transform 1 0 140 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8663
timestamp 1680363874
transform 1 0 148 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7943
timestamp 1680363874
transform 1 0 172 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8789
timestamp 1680363874
transform 1 0 172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8664
timestamp 1680363874
transform 1 0 228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8790
timestamp 1680363874
transform 1 0 196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8791
timestamp 1680363874
transform 1 0 300 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7981
timestamp 1680363874
transform 1 0 300 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8665
timestamp 1680363874
transform 1 0 316 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7878
timestamp 1680363874
transform 1 0 348 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7891
timestamp 1680363874
transform 1 0 340 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8792
timestamp 1680363874
transform 1 0 332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8652
timestamp 1680363874
transform 1 0 340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8666
timestamp 1680363874
transform 1 0 340 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7982
timestamp 1680363874
transform 1 0 340 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7908
timestamp 1680363874
transform 1 0 364 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8793
timestamp 1680363874
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8794
timestamp 1680363874
transform 1 0 364 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7879
timestamp 1680363874
transform 1 0 404 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7892
timestamp 1680363874
transform 1 0 404 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7909
timestamp 1680363874
transform 1 0 388 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8667
timestamp 1680363874
transform 1 0 380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8668
timestamp 1680363874
transform 1 0 388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8669
timestamp 1680363874
transform 1 0 404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8670
timestamp 1680363874
transform 1 0 420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8795
timestamp 1680363874
transform 1 0 388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8796
timestamp 1680363874
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8797
timestamp 1680363874
transform 1 0 412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8671
timestamp 1680363874
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8798
timestamp 1680363874
transform 1 0 436 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8799
timestamp 1680363874
transform 1 0 484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8672
timestamp 1680363874
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8673
timestamp 1680363874
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8800
timestamp 1680363874
transform 1 0 524 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7967
timestamp 1680363874
transform 1 0 596 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7983
timestamp 1680363874
transform 1 0 572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7944
timestamp 1680363874
transform 1 0 612 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8801
timestamp 1680363874
transform 1 0 628 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7945
timestamp 1680363874
transform 1 0 644 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8011
timestamp 1680363874
transform 1 0 644 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8674
timestamp 1680363874
transform 1 0 668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8675
timestamp 1680363874
transform 1 0 684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8802
timestamp 1680363874
transform 1 0 660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7968
timestamp 1680363874
transform 1 0 668 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8803
timestamp 1680363874
transform 1 0 676 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7984
timestamp 1680363874
transform 1 0 676 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8804
timestamp 1680363874
transform 1 0 716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8805
timestamp 1680363874
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8676
timestamp 1680363874
transform 1 0 748 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7969
timestamp 1680363874
transform 1 0 740 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8806
timestamp 1680363874
transform 1 0 748 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7946
timestamp 1680363874
transform 1 0 812 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8807
timestamp 1680363874
transform 1 0 812 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7861
timestamp 1680363874
transform 1 0 828 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7862
timestamp 1680363874
transform 1 0 868 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8677
timestamp 1680363874
transform 1 0 884 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7947
timestamp 1680363874
transform 1 0 892 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8678
timestamp 1680363874
transform 1 0 940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8808
timestamp 1680363874
transform 1 0 860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7880
timestamp 1680363874
transform 1 0 1100 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7881
timestamp 1680363874
transform 1 0 1116 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8679
timestamp 1680363874
transform 1 0 1052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8680
timestamp 1680363874
transform 1 0 1084 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8809
timestamp 1680363874
transform 1 0 1132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8649
timestamp 1680363874
transform 1 0 1148 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_8653
timestamp 1680363874
transform 1 0 1148 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7854
timestamp 1680363874
transform 1 0 1164 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_8650
timestamp 1680363874
transform 1 0 1188 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_7970
timestamp 1680363874
transform 1 0 1172 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7948
timestamp 1680363874
transform 1 0 1196 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7855
timestamp 1680363874
transform 1 0 1220 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_8654
timestamp 1680363874
transform 1 0 1212 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7910
timestamp 1680363874
transform 1 0 1236 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8655
timestamp 1680363874
transform 1 0 1260 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8681
timestamp 1680363874
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8682
timestamp 1680363874
transform 1 0 1236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8683
timestamp 1680363874
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8810
timestamp 1680363874
transform 1 0 1228 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7949
timestamp 1680363874
transform 1 0 1260 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8811
timestamp 1680363874
transform 1 0 1268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7882
timestamp 1680363874
transform 1 0 1300 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8651
timestamp 1680363874
transform 1 0 1300 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_7911
timestamp 1680363874
transform 1 0 1292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8656
timestamp 1680363874
transform 1 0 1308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8684
timestamp 1680363874
transform 1 0 1292 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7971
timestamp 1680363874
transform 1 0 1300 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7893
timestamp 1680363874
transform 1 0 1324 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8685
timestamp 1680363874
transform 1 0 1324 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7985
timestamp 1680363874
transform 1 0 1348 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8812
timestamp 1680363874
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7986
timestamp 1680363874
transform 1 0 1372 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8686
timestamp 1680363874
transform 1 0 1388 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7863
timestamp 1680363874
transform 1 0 1420 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7912
timestamp 1680363874
transform 1 0 1412 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8813
timestamp 1680363874
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7864
timestamp 1680363874
transform 1 0 1460 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8687
timestamp 1680363874
transform 1 0 1460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8814
timestamp 1680363874
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7913
timestamp 1680363874
transform 1 0 1476 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8688
timestamp 1680363874
transform 1 0 1476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8815
timestamp 1680363874
transform 1 0 1484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8816
timestamp 1680363874
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7914
timestamp 1680363874
transform 1 0 1516 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8689
timestamp 1680363874
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8817
timestamp 1680363874
transform 1 0 1516 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8690
timestamp 1680363874
transform 1 0 1524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8691
timestamp 1680363874
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7987
timestamp 1680363874
transform 1 0 1532 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8692
timestamp 1680363874
transform 1 0 1556 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7915
timestamp 1680363874
transform 1 0 1588 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8818
timestamp 1680363874
transform 1 0 1580 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7988
timestamp 1680363874
transform 1 0 1580 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7894
timestamp 1680363874
transform 1 0 1604 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7916
timestamp 1680363874
transform 1 0 1604 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8693
timestamp 1680363874
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8819
timestamp 1680363874
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8820
timestamp 1680363874
transform 1 0 1620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8821
timestamp 1680363874
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8822
timestamp 1680363874
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8694
timestamp 1680363874
transform 1 0 1692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8695
timestamp 1680363874
transform 1 0 1700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8696
timestamp 1680363874
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8697
timestamp 1680363874
transform 1 0 1740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8823
timestamp 1680363874
transform 1 0 1700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8824
timestamp 1680363874
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8825
timestamp 1680363874
transform 1 0 1732 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7865
timestamp 1680363874
transform 1 0 1756 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8826
timestamp 1680363874
transform 1 0 1756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8698
timestamp 1680363874
transform 1 0 1764 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7866
timestamp 1680363874
transform 1 0 1796 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8699
timestamp 1680363874
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8827
timestamp 1680363874
transform 1 0 1852 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7989
timestamp 1680363874
transform 1 0 1772 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7867
timestamp 1680363874
transform 1 0 1980 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7883
timestamp 1680363874
transform 1 0 1900 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8700
timestamp 1680363874
transform 1 0 1948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8828
timestamp 1680363874
transform 1 0 1900 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7990
timestamp 1680363874
transform 1 0 1932 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8701
timestamp 1680363874
transform 1 0 2004 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7917
timestamp 1680363874
transform 1 0 2068 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8702
timestamp 1680363874
transform 1 0 2028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8703
timestamp 1680363874
transform 1 0 2044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8704
timestamp 1680363874
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8705
timestamp 1680363874
transform 1 0 2068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8829
timestamp 1680363874
transform 1 0 2052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8706
timestamp 1680363874
transform 1 0 2100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8830
timestamp 1680363874
transform 1 0 2116 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7950
timestamp 1680363874
transform 1 0 2148 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8831
timestamp 1680363874
transform 1 0 2156 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7918
timestamp 1680363874
transform 1 0 2180 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8707
timestamp 1680363874
transform 1 0 2180 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7951
timestamp 1680363874
transform 1 0 2196 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8832
timestamp 1680363874
transform 1 0 2196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8648
timestamp 1680363874
transform 1 0 2204 0 1 645
box -2 -2 2 2
use M2_M1  M2_M1_8708
timestamp 1680363874
transform 1 0 2204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8833
timestamp 1680363874
transform 1 0 2204 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7884
timestamp 1680363874
transform 1 0 2236 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7919
timestamp 1680363874
transform 1 0 2228 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7856
timestamp 1680363874
transform 1 0 2260 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7920
timestamp 1680363874
transform 1 0 2244 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8657
timestamp 1680363874
transform 1 0 2260 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8709
timestamp 1680363874
transform 1 0 2244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8710
timestamp 1680363874
transform 1 0 2260 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7952
timestamp 1680363874
transform 1 0 2268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7991
timestamp 1680363874
transform 1 0 2260 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8834
timestamp 1680363874
transform 1 0 2276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8711
timestamp 1680363874
transform 1 0 2300 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7857
timestamp 1680363874
transform 1 0 2348 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7885
timestamp 1680363874
transform 1 0 2324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7921
timestamp 1680363874
transform 1 0 2316 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7992
timestamp 1680363874
transform 1 0 2308 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8712
timestamp 1680363874
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8835
timestamp 1680363874
transform 1 0 2324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8836
timestamp 1680363874
transform 1 0 2332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7868
timestamp 1680363874
transform 1 0 2364 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8658
timestamp 1680363874
transform 1 0 2356 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8713
timestamp 1680363874
transform 1 0 2372 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7953
timestamp 1680363874
transform 1 0 2380 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8714
timestamp 1680363874
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8837
timestamp 1680363874
transform 1 0 2356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8838
timestamp 1680363874
transform 1 0 2364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8839
timestamp 1680363874
transform 1 0 2380 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7993
timestamp 1680363874
transform 1 0 2356 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7858
timestamp 1680363874
transform 1 0 2412 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7869
timestamp 1680363874
transform 1 0 2404 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7922
timestamp 1680363874
transform 1 0 2404 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8659
timestamp 1680363874
transform 1 0 2412 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8840
timestamp 1680363874
transform 1 0 2412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7886
timestamp 1680363874
transform 1 0 2444 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7923
timestamp 1680363874
transform 1 0 2436 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8841
timestamp 1680363874
transform 1 0 2420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7994
timestamp 1680363874
transform 1 0 2412 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7859
timestamp 1680363874
transform 1 0 2460 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7924
timestamp 1680363874
transform 1 0 2452 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8715
timestamp 1680363874
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8716
timestamp 1680363874
transform 1 0 2452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8842
timestamp 1680363874
transform 1 0 2444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8843
timestamp 1680363874
transform 1 0 2452 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8012
timestamp 1680363874
transform 1 0 2452 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8717
timestamp 1680363874
transform 1 0 2500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8844
timestamp 1680363874
transform 1 0 2492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8845
timestamp 1680363874
transform 1 0 2508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8846
timestamp 1680363874
transform 1 0 2516 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7995
timestamp 1680363874
transform 1 0 2508 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7860
timestamp 1680363874
transform 1 0 2532 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_8660
timestamp 1680363874
transform 1 0 2532 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8718
timestamp 1680363874
transform 1 0 2556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8719
timestamp 1680363874
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8847
timestamp 1680363874
transform 1 0 2564 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7954
timestamp 1680363874
transform 1 0 2612 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8720
timestamp 1680363874
transform 1 0 2620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8721
timestamp 1680363874
transform 1 0 2644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8848
timestamp 1680363874
transform 1 0 2604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8849
timestamp 1680363874
transform 1 0 2612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8850
timestamp 1680363874
transform 1 0 2636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8851
timestamp 1680363874
transform 1 0 2660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8722
timestamp 1680363874
transform 1 0 2684 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7972
timestamp 1680363874
transform 1 0 2684 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8852
timestamp 1680363874
transform 1 0 2708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7996
timestamp 1680363874
transform 1 0 2708 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7925
timestamp 1680363874
transform 1 0 2780 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8723
timestamp 1680363874
transform 1 0 2780 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7955
timestamp 1680363874
transform 1 0 2796 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8724
timestamp 1680363874
transform 1 0 2812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8725
timestamp 1680363874
transform 1 0 2820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8853
timestamp 1680363874
transform 1 0 2732 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7997
timestamp 1680363874
transform 1 0 2732 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7956
timestamp 1680363874
transform 1 0 2828 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8726
timestamp 1680363874
transform 1 0 2844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8854
timestamp 1680363874
transform 1 0 2828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8907
timestamp 1680363874
transform 1 0 2836 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7895
timestamp 1680363874
transform 1 0 2860 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8727
timestamp 1680363874
transform 1 0 2868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8855
timestamp 1680363874
transform 1 0 2860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7973
timestamp 1680363874
transform 1 0 2868 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8908
timestamp 1680363874
transform 1 0 2868 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_8013
timestamp 1680363874
transform 1 0 2868 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7896
timestamp 1680363874
transform 1 0 2892 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7926
timestamp 1680363874
transform 1 0 2900 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8728
timestamp 1680363874
transform 1 0 2900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8856
timestamp 1680363874
transform 1 0 2892 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7957
timestamp 1680363874
transform 1 0 2916 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8857
timestamp 1680363874
transform 1 0 2908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8858
timestamp 1680363874
transform 1 0 2916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8729
timestamp 1680363874
transform 1 0 2924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8730
timestamp 1680363874
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8859
timestamp 1680363874
transform 1 0 2932 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7998
timestamp 1680363874
transform 1 0 2932 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8731
timestamp 1680363874
transform 1 0 2956 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7958
timestamp 1680363874
transform 1 0 2964 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8860
timestamp 1680363874
transform 1 0 2964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8732
timestamp 1680363874
transform 1 0 2996 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7974
timestamp 1680363874
transform 1 0 2996 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7870
timestamp 1680363874
transform 1 0 3012 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8733
timestamp 1680363874
transform 1 0 3036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8734
timestamp 1680363874
transform 1 0 3092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8861
timestamp 1680363874
transform 1 0 3012 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7999
timestamp 1680363874
transform 1 0 3092 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8735
timestamp 1680363874
transform 1 0 3140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8736
timestamp 1680363874
transform 1 0 3156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8737
timestamp 1680363874
transform 1 0 3164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8862
timestamp 1680363874
transform 1 0 3132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8863
timestamp 1680363874
transform 1 0 3148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8000
timestamp 1680363874
transform 1 0 3132 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8001
timestamp 1680363874
transform 1 0 3164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8014
timestamp 1680363874
transform 1 0 3148 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8864
timestamp 1680363874
transform 1 0 3180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8015
timestamp 1680363874
transform 1 0 3180 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8909
timestamp 1680363874
transform 1 0 3204 0 1 585
box -2 -2 2 2
use M2_M1  M2_M1_8865
timestamp 1680363874
transform 1 0 3212 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7975
timestamp 1680363874
transform 1 0 3228 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8002
timestamp 1680363874
transform 1 0 3220 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8910
timestamp 1680363874
transform 1 0 3220 0 1 585
box -2 -2 2 2
use M3_M2  M3_M2_7897
timestamp 1680363874
transform 1 0 3244 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8738
timestamp 1680363874
transform 1 0 3268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8739
timestamp 1680363874
transform 1 0 3276 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7927
timestamp 1680363874
transform 1 0 3292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8866
timestamp 1680363874
transform 1 0 3292 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7928
timestamp 1680363874
transform 1 0 3324 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7959
timestamp 1680363874
transform 1 0 3308 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8740
timestamp 1680363874
transform 1 0 3324 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7960
timestamp 1680363874
transform 1 0 3332 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8867
timestamp 1680363874
transform 1 0 3300 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8016
timestamp 1680363874
transform 1 0 3300 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8741
timestamp 1680363874
transform 1 0 3348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8868
timestamp 1680363874
transform 1 0 3332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8869
timestamp 1680363874
transform 1 0 3340 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7976
timestamp 1680363874
transform 1 0 3348 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7929
timestamp 1680363874
transform 1 0 3372 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7930
timestamp 1680363874
transform 1 0 3428 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8742
timestamp 1680363874
transform 1 0 3372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8743
timestamp 1680363874
transform 1 0 3380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8744
timestamp 1680363874
transform 1 0 3436 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7961
timestamp 1680363874
transform 1 0 3460 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8745
timestamp 1680363874
transform 1 0 3476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8870
timestamp 1680363874
transform 1 0 3460 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8003
timestamp 1680363874
transform 1 0 3500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7898
timestamp 1680363874
transform 1 0 3540 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7899
timestamp 1680363874
transform 1 0 3556 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7931
timestamp 1680363874
transform 1 0 3524 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8746
timestamp 1680363874
transform 1 0 3524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8747
timestamp 1680363874
transform 1 0 3540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8748
timestamp 1680363874
transform 1 0 3556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8871
timestamp 1680363874
transform 1 0 3524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8872
timestamp 1680363874
transform 1 0 3532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8873
timestamp 1680363874
transform 1 0 3556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8004
timestamp 1680363874
transform 1 0 3556 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7932
timestamp 1680363874
transform 1 0 3580 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8749
timestamp 1680363874
transform 1 0 3580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8750
timestamp 1680363874
transform 1 0 3596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8751
timestamp 1680363874
transform 1 0 3612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8752
timestamp 1680363874
transform 1 0 3620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8874
timestamp 1680363874
transform 1 0 3572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8875
timestamp 1680363874
transform 1 0 3580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8876
timestamp 1680363874
transform 1 0 3604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8877
timestamp 1680363874
transform 1 0 3628 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7871
timestamp 1680363874
transform 1 0 3668 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7872
timestamp 1680363874
transform 1 0 3708 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8753
timestamp 1680363874
transform 1 0 3684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8754
timestamp 1680363874
transform 1 0 3732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8878
timestamp 1680363874
transform 1 0 3716 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7962
timestamp 1680363874
transform 1 0 3740 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8017
timestamp 1680363874
transform 1 0 3732 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8879
timestamp 1680363874
transform 1 0 3764 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7963
timestamp 1680363874
transform 1 0 3780 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8755
timestamp 1680363874
transform 1 0 3804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8880
timestamp 1680363874
transform 1 0 3780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8881
timestamp 1680363874
transform 1 0 3796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8882
timestamp 1680363874
transform 1 0 3820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8756
timestamp 1680363874
transform 1 0 3868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8883
timestamp 1680363874
transform 1 0 3860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8005
timestamp 1680363874
transform 1 0 3860 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7933
timestamp 1680363874
transform 1 0 3892 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8757
timestamp 1680363874
transform 1 0 3892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8758
timestamp 1680363874
transform 1 0 3908 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7964
timestamp 1680363874
transform 1 0 3916 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8884
timestamp 1680363874
transform 1 0 3892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8885
timestamp 1680363874
transform 1 0 3916 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8006
timestamp 1680363874
transform 1 0 3908 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8759
timestamp 1680363874
transform 1 0 3948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8886
timestamp 1680363874
transform 1 0 3940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7977
timestamp 1680363874
transform 1 0 3948 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8760
timestamp 1680363874
transform 1 0 3972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8761
timestamp 1680363874
transform 1 0 3988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8762
timestamp 1680363874
transform 1 0 3996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8887
timestamp 1680363874
transform 1 0 3980 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7978
timestamp 1680363874
transform 1 0 3996 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8007
timestamp 1680363874
transform 1 0 3972 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8008
timestamp 1680363874
transform 1 0 4020 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8018
timestamp 1680363874
transform 1 0 4028 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7887
timestamp 1680363874
transform 1 0 4044 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7900
timestamp 1680363874
transform 1 0 4140 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7901
timestamp 1680363874
transform 1 0 4180 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7934
timestamp 1680363874
transform 1 0 4076 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7935
timestamp 1680363874
transform 1 0 4116 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8763
timestamp 1680363874
transform 1 0 4044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8764
timestamp 1680363874
transform 1 0 4060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8765
timestamp 1680363874
transform 1 0 4076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8888
timestamp 1680363874
transform 1 0 4036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8889
timestamp 1680363874
transform 1 0 4068 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8019
timestamp 1680363874
transform 1 0 4052 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7965
timestamp 1680363874
transform 1 0 4092 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8766
timestamp 1680363874
transform 1 0 4140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8767
timestamp 1680363874
transform 1 0 4172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8768
timestamp 1680363874
transform 1 0 4180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8890
timestamp 1680363874
transform 1 0 4092 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8891
timestamp 1680363874
transform 1 0 4180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8009
timestamp 1680363874
transform 1 0 4156 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7873
timestamp 1680363874
transform 1 0 4252 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7874
timestamp 1680363874
transform 1 0 4276 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7936
timestamp 1680363874
transform 1 0 4292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7937
timestamp 1680363874
transform 1 0 4332 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7966
timestamp 1680363874
transform 1 0 4244 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8769
timestamp 1680363874
transform 1 0 4292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8770
timestamp 1680363874
transform 1 0 4324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8771
timestamp 1680363874
transform 1 0 4332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8892
timestamp 1680363874
transform 1 0 4244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8893
timestamp 1680363874
transform 1 0 4332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7902
timestamp 1680363874
transform 1 0 4348 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8772
timestamp 1680363874
transform 1 0 4348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8773
timestamp 1680363874
transform 1 0 4380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8894
timestamp 1680363874
transform 1 0 4372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8895
timestamp 1680363874
transform 1 0 4388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8896
timestamp 1680363874
transform 1 0 4396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7875
timestamp 1680363874
transform 1 0 4412 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7888
timestamp 1680363874
transform 1 0 4412 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8774
timestamp 1680363874
transform 1 0 4412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8897
timestamp 1680363874
transform 1 0 4412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7889
timestamp 1680363874
transform 1 0 4476 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7903
timestamp 1680363874
transform 1 0 4476 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7876
timestamp 1680363874
transform 1 0 4516 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8775
timestamp 1680363874
transform 1 0 4460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8776
timestamp 1680363874
transform 1 0 4508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8898
timestamp 1680363874
transform 1 0 4428 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8020
timestamp 1680363874
transform 1 0 4428 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8021
timestamp 1680363874
transform 1 0 4532 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7904
timestamp 1680363874
transform 1 0 4556 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7938
timestamp 1680363874
transform 1 0 4548 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8777
timestamp 1680363874
transform 1 0 4556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8899
timestamp 1680363874
transform 1 0 4548 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7890
timestamp 1680363874
transform 1 0 4572 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8778
timestamp 1680363874
transform 1 0 4572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8900
timestamp 1680363874
transform 1 0 4572 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7905
timestamp 1680363874
transform 1 0 4588 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7877
timestamp 1680363874
transform 1 0 4620 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7939
timestamp 1680363874
transform 1 0 4604 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8779
timestamp 1680363874
transform 1 0 4604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8780
timestamp 1680363874
transform 1 0 4620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8781
timestamp 1680363874
transform 1 0 4628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8901
timestamp 1680363874
transform 1 0 4596 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7979
timestamp 1680363874
transform 1 0 4604 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8902
timestamp 1680363874
transform 1 0 4612 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7980
timestamp 1680363874
transform 1 0 4628 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7906
timestamp 1680363874
transform 1 0 4668 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8782
timestamp 1680363874
transform 1 0 4644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8783
timestamp 1680363874
transform 1 0 4660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8784
timestamp 1680363874
transform 1 0 4684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8903
timestamp 1680363874
transform 1 0 4652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8904
timestamp 1680363874
transform 1 0 4668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8905
timestamp 1680363874
transform 1 0 4676 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7907
timestamp 1680363874
transform 1 0 4700 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7940
timestamp 1680363874
transform 1 0 4692 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7941
timestamp 1680363874
transform 1 0 4732 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8785
timestamp 1680363874
transform 1 0 4692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8786
timestamp 1680363874
transform 1 0 4700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8787
timestamp 1680363874
transform 1 0 4732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8906
timestamp 1680363874
transform 1 0 4780 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8010
timestamp 1680363874
transform 1 0 4868 0 1 595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_82
timestamp 1680363874
transform 1 0 48 0 1 570
box -10 -3 10 3
use INVX2  INVX2_605
timestamp 1680363874
transform 1 0 72 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_8022
timestamp 1680363874
transform 1 0 172 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_540
timestamp 1680363874
transform -1 0 184 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_541
timestamp 1680363874
transform 1 0 184 0 1 570
box -8 -3 104 105
use INVX2  INVX2_606
timestamp 1680363874
transform 1 0 280 0 1 570
box -9 -3 26 105
use FILL  FILL_9765
timestamp 1680363874
transform 1 0 296 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_166
timestamp 1680363874
transform 1 0 304 0 1 570
box -8 -3 34 105
use FILL  FILL_9766
timestamp 1680363874
transform 1 0 336 0 1 570
box -8 -3 16 105
use INVX2  INVX2_607
timestamp 1680363874
transform -1 0 360 0 1 570
box -9 -3 26 105
use INVX2  INVX2_608
timestamp 1680363874
transform 1 0 360 0 1 570
box -9 -3 26 105
use FILL  FILL_9767
timestamp 1680363874
transform 1 0 376 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_351
timestamp 1680363874
transform 1 0 384 0 1 570
box -8 -3 46 105
use FILL  FILL_9768
timestamp 1680363874
transform 1 0 424 0 1 570
box -8 -3 16 105
use FILL  FILL_9769
timestamp 1680363874
transform 1 0 432 0 1 570
box -8 -3 16 105
use FILL  FILL_9770
timestamp 1680363874
transform 1 0 440 0 1 570
box -8 -3 16 105
use FILL  FILL_9771
timestamp 1680363874
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_9772
timestamp 1680363874
transform 1 0 456 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8023
timestamp 1680363874
transform 1 0 484 0 1 575
box -3 -3 3 3
use BUFX2  BUFX2_100
timestamp 1680363874
transform 1 0 464 0 1 570
box -5 -3 28 105
use FILL  FILL_9773
timestamp 1680363874
transform 1 0 488 0 1 570
box -8 -3 16 105
use FILL  FILL_9774
timestamp 1680363874
transform 1 0 496 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8024
timestamp 1680363874
transform 1 0 516 0 1 575
box -3 -3 3 3
use FILL  FILL_9775
timestamp 1680363874
transform 1 0 504 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_542
timestamp 1680363874
transform 1 0 512 0 1 570
box -8 -3 104 105
use FILL  FILL_9776
timestamp 1680363874
transform 1 0 608 0 1 570
box -8 -3 16 105
use FILL  FILL_9777
timestamp 1680363874
transform 1 0 616 0 1 570
box -8 -3 16 105
use FILL  FILL_9778
timestamp 1680363874
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_9779
timestamp 1680363874
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_9780
timestamp 1680363874
transform 1 0 640 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8025
timestamp 1680363874
transform 1 0 660 0 1 575
box -3 -3 3 3
use FILL  FILL_9804
timestamp 1680363874
transform 1 0 648 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_380
timestamp 1680363874
transform -1 0 696 0 1 570
box -8 -3 46 105
use FILL  FILL_9805
timestamp 1680363874
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_9806
timestamp 1680363874
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_9807
timestamp 1680363874
transform 1 0 712 0 1 570
box -8 -3 16 105
use FILL  FILL_9808
timestamp 1680363874
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_9809
timestamp 1680363874
transform 1 0 728 0 1 570
box -8 -3 16 105
use FILL  FILL_9810
timestamp 1680363874
transform 1 0 736 0 1 570
box -8 -3 16 105
use INVX2  INVX2_613
timestamp 1680363874
transform 1 0 744 0 1 570
box -9 -3 26 105
use FILL  FILL_9811
timestamp 1680363874
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_9815
timestamp 1680363874
transform 1 0 768 0 1 570
box -8 -3 16 105
use FILL  FILL_9817
timestamp 1680363874
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_9819
timestamp 1680363874
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_9820
timestamp 1680363874
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_9821
timestamp 1680363874
transform 1 0 800 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8026
timestamp 1680363874
transform 1 0 820 0 1 575
box -3 -3 3 3
use FILL  FILL_9822
timestamp 1680363874
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_9823
timestamp 1680363874
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_9824
timestamp 1680363874
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_9826
timestamp 1680363874
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_9828
timestamp 1680363874
transform 1 0 840 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_545
timestamp 1680363874
transform 1 0 848 0 1 570
box -8 -3 104 105
use FILL  FILL_9830
timestamp 1680363874
transform 1 0 944 0 1 570
box -8 -3 16 105
use FILL  FILL_9837
timestamp 1680363874
transform 1 0 952 0 1 570
box -8 -3 16 105
use FILL  FILL_9839
timestamp 1680363874
transform 1 0 960 0 1 570
box -8 -3 16 105
use FILL  FILL_9841
timestamp 1680363874
transform 1 0 968 0 1 570
box -8 -3 16 105
use FILL  FILL_9843
timestamp 1680363874
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_9845
timestamp 1680363874
transform 1 0 984 0 1 570
box -8 -3 16 105
use FILL  FILL_9846
timestamp 1680363874
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_9847
timestamp 1680363874
transform 1 0 1000 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8027
timestamp 1680363874
transform 1 0 1020 0 1 575
box -3 -3 3 3
use FILL  FILL_9848
timestamp 1680363874
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_9849
timestamp 1680363874
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_9851
timestamp 1680363874
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_9853
timestamp 1680363874
transform 1 0 1032 0 1 570
box -8 -3 16 105
use FILL  FILL_9855
timestamp 1680363874
transform 1 0 1040 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_546
timestamp 1680363874
transform -1 0 1144 0 1 570
box -8 -3 104 105
use FILL  FILL_9856
timestamp 1680363874
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_9857
timestamp 1680363874
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_9858
timestamp 1680363874
transform 1 0 1160 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1680363874
transform 1 0 1168 0 1 570
box -8 -3 40 105
use FILL  FILL_9859
timestamp 1680363874
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_9860
timestamp 1680363874
transform 1 0 1208 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_353
timestamp 1680363874
transform -1 0 1256 0 1 570
box -8 -3 46 105
use FILL  FILL_9861
timestamp 1680363874
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_9862
timestamp 1680363874
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_9863
timestamp 1680363874
transform 1 0 1272 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_74
timestamp 1680363874
transform 1 0 1280 0 1 570
box -8 -3 40 105
use FILL  FILL_9864
timestamp 1680363874
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_9865
timestamp 1680363874
transform 1 0 1320 0 1 570
box -8 -3 16 105
use FILL  FILL_9866
timestamp 1680363874
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_9867
timestamp 1680363874
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_9868
timestamp 1680363874
transform 1 0 1344 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_101
timestamp 1680363874
transform 1 0 1352 0 1 570
box -5 -3 28 105
use FILL  FILL_9869
timestamp 1680363874
transform 1 0 1376 0 1 570
box -8 -3 16 105
use FILL  FILL_9870
timestamp 1680363874
transform 1 0 1384 0 1 570
box -8 -3 16 105
use FILL  FILL_9871
timestamp 1680363874
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_9872
timestamp 1680363874
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_9873
timestamp 1680363874
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_9888
timestamp 1680363874
transform 1 0 1416 0 1 570
box -8 -3 16 105
use FILL  FILL_9890
timestamp 1680363874
transform 1 0 1424 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_385
timestamp 1680363874
transform 1 0 1432 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_8028
timestamp 1680363874
transform 1 0 1484 0 1 575
box -3 -3 3 3
use FILL  FILL_9891
timestamp 1680363874
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_9892
timestamp 1680363874
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_9893
timestamp 1680363874
transform 1 0 1488 0 1 570
box -8 -3 16 105
use INVX2  INVX2_618
timestamp 1680363874
transform 1 0 1496 0 1 570
box -9 -3 26 105
use INVX2  INVX2_619
timestamp 1680363874
transform 1 0 1512 0 1 570
box -9 -3 26 105
use FILL  FILL_9894
timestamp 1680363874
transform 1 0 1528 0 1 570
box -8 -3 16 105
use FILL  FILL_9897
timestamp 1680363874
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_9899
timestamp 1680363874
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_9901
timestamp 1680363874
transform 1 0 1552 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_102
timestamp 1680363874
transform 1 0 1560 0 1 570
box -5 -3 28 105
use FILL  FILL_9903
timestamp 1680363874
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_9904
timestamp 1680363874
transform 1 0 1592 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_103
timestamp 1680363874
transform 1 0 1600 0 1 570
box -5 -3 28 105
use FILL  FILL_9905
timestamp 1680363874
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_9910
timestamp 1680363874
transform 1 0 1632 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_104
timestamp 1680363874
transform -1 0 1664 0 1 570
box -5 -3 28 105
use FILL  FILL_9911
timestamp 1680363874
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_9912
timestamp 1680363874
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_9913
timestamp 1680363874
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_9916
timestamp 1680363874
transform 1 0 1688 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8029
timestamp 1680363874
transform 1 0 1732 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_386
timestamp 1680363874
transform 1 0 1696 0 1 570
box -8 -3 46 105
use INVX2  INVX2_620
timestamp 1680363874
transform -1 0 1752 0 1 570
box -9 -3 26 105
use FILL  FILL_9918
timestamp 1680363874
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_9925
timestamp 1680363874
transform 1 0 1760 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8030
timestamp 1680363874
transform 1 0 1868 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_549
timestamp 1680363874
transform -1 0 1864 0 1 570
box -8 -3 104 105
use FILL  FILL_9926
timestamp 1680363874
transform 1 0 1864 0 1 570
box -8 -3 16 105
use FILL  FILL_9927
timestamp 1680363874
transform 1 0 1872 0 1 570
box -8 -3 16 105
use FILL  FILL_9928
timestamp 1680363874
transform 1 0 1880 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_550
timestamp 1680363874
transform 1 0 1888 0 1 570
box -8 -3 104 105
use FILL  FILL_9929
timestamp 1680363874
transform 1 0 1984 0 1 570
box -8 -3 16 105
use INVX2  INVX2_622
timestamp 1680363874
transform 1 0 1992 0 1 570
box -9 -3 26 105
use FILL  FILL_9943
timestamp 1680363874
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_9947
timestamp 1680363874
transform 1 0 2016 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8031
timestamp 1680363874
transform 1 0 2060 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_358
timestamp 1680363874
transform -1 0 2064 0 1 570
box -8 -3 46 105
use FILL  FILL_9948
timestamp 1680363874
transform 1 0 2064 0 1 570
box -8 -3 16 105
use FILL  FILL_9949
timestamp 1680363874
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_9950
timestamp 1680363874
transform 1 0 2080 0 1 570
box -8 -3 16 105
use FILL  FILL_9953
timestamp 1680363874
transform 1 0 2088 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8032
timestamp 1680363874
transform 1 0 2108 0 1 575
box -3 -3 3 3
use BUFX2  BUFX2_107
timestamp 1680363874
transform 1 0 2096 0 1 570
box -5 -3 28 105
use FILL  FILL_9955
timestamp 1680363874
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_9956
timestamp 1680363874
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_9957
timestamp 1680363874
transform 1 0 2136 0 1 570
box -8 -3 16 105
use FILL  FILL_9958
timestamp 1680363874
transform 1 0 2144 0 1 570
box -8 -3 16 105
use FILL  FILL_9959
timestamp 1680363874
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_9960
timestamp 1680363874
transform 1 0 2160 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_168
timestamp 1680363874
transform 1 0 2168 0 1 570
box -8 -3 34 105
use FILL  FILL_9961
timestamp 1680363874
transform 1 0 2200 0 1 570
box -8 -3 16 105
use FILL  FILL_9964
timestamp 1680363874
transform 1 0 2208 0 1 570
box -8 -3 16 105
use FILL  FILL_9966
timestamp 1680363874
transform 1 0 2216 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8033
timestamp 1680363874
transform 1 0 2236 0 1 575
box -3 -3 3 3
use FILL  FILL_9967
timestamp 1680363874
transform 1 0 2224 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_169
timestamp 1680363874
transform 1 0 2232 0 1 570
box -8 -3 34 105
use FILL  FILL_9968
timestamp 1680363874
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_9969
timestamp 1680363874
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_9971
timestamp 1680363874
transform 1 0 2280 0 1 570
box -8 -3 16 105
use FILL  FILL_9973
timestamp 1680363874
transform 1 0 2288 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_108
timestamp 1680363874
transform 1 0 2296 0 1 570
box -5 -3 28 105
use FILL  FILL_9975
timestamp 1680363874
transform 1 0 2320 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_170
timestamp 1680363874
transform 1 0 2328 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_8034
timestamp 1680363874
transform 1 0 2388 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_390
timestamp 1680363874
transform 1 0 2360 0 1 570
box -8 -3 46 105
use FILL  FILL_9976
timestamp 1680363874
transform 1 0 2400 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8035
timestamp 1680363874
transform 1 0 2420 0 1 575
box -3 -3 3 3
use FILL  FILL_9977
timestamp 1680363874
transform 1 0 2408 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8036
timestamp 1680363874
transform 1 0 2444 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_171
timestamp 1680363874
transform -1 0 2448 0 1 570
box -8 -3 34 105
use FILL  FILL_9978
timestamp 1680363874
transform 1 0 2448 0 1 570
box -8 -3 16 105
use FILL  FILL_9993
timestamp 1680363874
transform 1 0 2456 0 1 570
box -8 -3 16 105
use FILL  FILL_9995
timestamp 1680363874
transform 1 0 2464 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_391
timestamp 1680363874
transform 1 0 2472 0 1 570
box -8 -3 46 105
use FILL  FILL_9997
timestamp 1680363874
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_10004
timestamp 1680363874
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_10006
timestamp 1680363874
transform 1 0 2528 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_173
timestamp 1680363874
transform -1 0 2568 0 1 570
box -8 -3 34 105
use FILL  FILL_10007
timestamp 1680363874
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_10008
timestamp 1680363874
transform 1 0 2576 0 1 570
box -8 -3 16 105
use FILL  FILL_10009
timestamp 1680363874
transform 1 0 2584 0 1 570
box -8 -3 16 105
use INVX2  INVX2_626
timestamp 1680363874
transform -1 0 2608 0 1 570
box -9 -3 26 105
use FILL  FILL_10010
timestamp 1680363874
transform 1 0 2608 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_392
timestamp 1680363874
transform 1 0 2616 0 1 570
box -8 -3 46 105
use FILL  FILL_10011
timestamp 1680363874
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_10019
timestamp 1680363874
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_10020
timestamp 1680363874
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_10021
timestamp 1680363874
transform 1 0 2680 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_110
timestamp 1680363874
transform 1 0 2688 0 1 570
box -5 -3 28 105
use FILL  FILL_10022
timestamp 1680363874
transform 1 0 2712 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_552
timestamp 1680363874
transform 1 0 2720 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_8037
timestamp 1680363874
transform 1 0 2828 0 1 575
box -3 -3 3 3
use NOR2X1  NOR2X1_113
timestamp 1680363874
transform -1 0 2840 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1680363874
transform -1 0 2864 0 1 570
box -8 -3 32 105
use FILL  FILL_10023
timestamp 1680363874
transform 1 0 2864 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_111
timestamp 1680363874
transform 1 0 2872 0 1 570
box -5 -3 28 105
use INVX2  INVX2_629
timestamp 1680363874
transform -1 0 2912 0 1 570
box -9 -3 26 105
use INVX2  INVX2_630
timestamp 1680363874
transform 1 0 2912 0 1 570
box -9 -3 26 105
use FILL  FILL_10029
timestamp 1680363874
transform 1 0 2928 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_359
timestamp 1680363874
transform -1 0 2976 0 1 570
box -8 -3 46 105
use FILL  FILL_10030
timestamp 1680363874
transform 1 0 2976 0 1 570
box -8 -3 16 105
use FILL  FILL_10045
timestamp 1680363874
transform 1 0 2984 0 1 570
box -8 -3 16 105
use FILL  FILL_10046
timestamp 1680363874
transform 1 0 2992 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_554
timestamp 1680363874
transform 1 0 3000 0 1 570
box -8 -3 104 105
use FILL  FILL_10047
timestamp 1680363874
transform 1 0 3096 0 1 570
box -8 -3 16 105
use FILL  FILL_10056
timestamp 1680363874
transform 1 0 3104 0 1 570
box -8 -3 16 105
use FILL  FILL_10058
timestamp 1680363874
transform 1 0 3112 0 1 570
box -8 -3 16 105
use FILL  FILL_10059
timestamp 1680363874
transform 1 0 3120 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8038
timestamp 1680363874
transform 1 0 3140 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_8039
timestamp 1680363874
transform 1 0 3172 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_395
timestamp 1680363874
transform -1 0 3168 0 1 570
box -8 -3 46 105
use FILL  FILL_10060
timestamp 1680363874
transform 1 0 3168 0 1 570
box -8 -3 16 105
use FILL  FILL_10064
timestamp 1680363874
transform 1 0 3176 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8040
timestamp 1680363874
transform 1 0 3204 0 1 575
box -3 -3 3 3
use INVX2  INVX2_632
timestamp 1680363874
transform -1 0 3200 0 1 570
box -9 -3 26 105
use FILL  FILL_10065
timestamp 1680363874
transform 1 0 3200 0 1 570
box -8 -3 16 105
use FILL  FILL_10066
timestamp 1680363874
transform 1 0 3208 0 1 570
box -8 -3 16 105
use FILL  FILL_10067
timestamp 1680363874
transform 1 0 3216 0 1 570
box -8 -3 16 105
use FILL  FILL_10068
timestamp 1680363874
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_10069
timestamp 1680363874
transform 1 0 3232 0 1 570
box -8 -3 16 105
use FILL  FILL_10073
timestamp 1680363874
transform 1 0 3240 0 1 570
box -8 -3 16 105
use FILL  FILL_10075
timestamp 1680363874
transform 1 0 3248 0 1 570
box -8 -3 16 105
use FILL  FILL_10077
timestamp 1680363874
transform 1 0 3256 0 1 570
box -8 -3 16 105
use INVX2  INVX2_633
timestamp 1680363874
transform -1 0 3280 0 1 570
box -9 -3 26 105
use FILL  FILL_10078
timestamp 1680363874
transform 1 0 3280 0 1 570
box -8 -3 16 105
use FILL  FILL_10081
timestamp 1680363874
transform 1 0 3288 0 1 570
box -8 -3 16 105
use FILL  FILL_10082
timestamp 1680363874
transform 1 0 3296 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_361
timestamp 1680363874
transform -1 0 3344 0 1 570
box -8 -3 46 105
use FILL  FILL_10083
timestamp 1680363874
transform 1 0 3344 0 1 570
box -8 -3 16 105
use FILL  FILL_10084
timestamp 1680363874
transform 1 0 3352 0 1 570
box -8 -3 16 105
use INVX2  INVX2_635
timestamp 1680363874
transform 1 0 3360 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_555
timestamp 1680363874
transform -1 0 3472 0 1 570
box -8 -3 104 105
use INVX2  INVX2_636
timestamp 1680363874
transform -1 0 3488 0 1 570
box -9 -3 26 105
use FILL  FILL_10085
timestamp 1680363874
transform 1 0 3488 0 1 570
box -8 -3 16 105
use FILL  FILL_10086
timestamp 1680363874
transform 1 0 3496 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8041
timestamp 1680363874
transform 1 0 3516 0 1 575
box -3 -3 3 3
use FILL  FILL_10087
timestamp 1680363874
transform 1 0 3504 0 1 570
box -8 -3 16 105
use FILL  FILL_10092
timestamp 1680363874
transform 1 0 3512 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8042
timestamp 1680363874
transform 1 0 3548 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_362
timestamp 1680363874
transform 1 0 3520 0 1 570
box -8 -3 46 105
use FILL  FILL_10094
timestamp 1680363874
transform 1 0 3560 0 1 570
box -8 -3 16 105
use FILL  FILL_10096
timestamp 1680363874
transform 1 0 3568 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_363
timestamp 1680363874
transform 1 0 3576 0 1 570
box -8 -3 46 105
use FILL  FILL_10097
timestamp 1680363874
transform 1 0 3616 0 1 570
box -8 -3 16 105
use FILL  FILL_10098
timestamp 1680363874
transform 1 0 3624 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_558
timestamp 1680363874
transform -1 0 3728 0 1 570
box -8 -3 104 105
use BUFX2  BUFX2_112
timestamp 1680363874
transform 1 0 3728 0 1 570
box -5 -3 28 105
use FILL  FILL_10099
timestamp 1680363874
transform 1 0 3752 0 1 570
box -8 -3 16 105
use FILL  FILL_10105
timestamp 1680363874
transform 1 0 3760 0 1 570
box -8 -3 16 105
use FILL  FILL_10107
timestamp 1680363874
transform 1 0 3768 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_398
timestamp 1680363874
transform 1 0 3776 0 1 570
box -8 -3 46 105
use FILL  FILL_10109
timestamp 1680363874
transform 1 0 3816 0 1 570
box -8 -3 16 105
use FILL  FILL_10114
timestamp 1680363874
transform 1 0 3824 0 1 570
box -8 -3 16 105
use FILL  FILL_10116
timestamp 1680363874
transform 1 0 3832 0 1 570
box -8 -3 16 105
use FILL  FILL_10118
timestamp 1680363874
transform 1 0 3840 0 1 570
box -8 -3 16 105
use FILL  FILL_10120
timestamp 1680363874
transform 1 0 3848 0 1 570
box -8 -3 16 105
use INVX2  INVX2_639
timestamp 1680363874
transform 1 0 3856 0 1 570
box -9 -3 26 105
use FILL  FILL_10121
timestamp 1680363874
transform 1 0 3872 0 1 570
box -8 -3 16 105
use FILL  FILL_10122
timestamp 1680363874
transform 1 0 3880 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_365
timestamp 1680363874
transform 1 0 3888 0 1 570
box -8 -3 46 105
use FILL  FILL_10123
timestamp 1680363874
transform 1 0 3928 0 1 570
box -8 -3 16 105
use FILL  FILL_10124
timestamp 1680363874
transform 1 0 3936 0 1 570
box -8 -3 16 105
use FILL  FILL_10125
timestamp 1680363874
transform 1 0 3944 0 1 570
box -8 -3 16 105
use FILL  FILL_10126
timestamp 1680363874
transform 1 0 3952 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8043
timestamp 1680363874
transform 1 0 3980 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_399
timestamp 1680363874
transform -1 0 4000 0 1 570
box -8 -3 46 105
use FILL  FILL_10127
timestamp 1680363874
transform 1 0 4000 0 1 570
box -8 -3 16 105
use FILL  FILL_10128
timestamp 1680363874
transform 1 0 4008 0 1 570
box -8 -3 16 105
use FILL  FILL_10129
timestamp 1680363874
transform 1 0 4016 0 1 570
box -8 -3 16 105
use FILL  FILL_10130
timestamp 1680363874
transform 1 0 4024 0 1 570
box -8 -3 16 105
use FILL  FILL_10131
timestamp 1680363874
transform 1 0 4032 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8044
timestamp 1680363874
transform 1 0 4068 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_366
timestamp 1680363874
transform -1 0 4080 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_560
timestamp 1680363874
transform 1 0 4080 0 1 570
box -8 -3 104 105
use INVX2  INVX2_640
timestamp 1680363874
transform 1 0 4176 0 1 570
box -9 -3 26 105
use FILL  FILL_10132
timestamp 1680363874
transform 1 0 4192 0 1 570
box -8 -3 16 105
use FILL  FILL_10133
timestamp 1680363874
transform 1 0 4200 0 1 570
box -8 -3 16 105
use FILL  FILL_10156
timestamp 1680363874
transform 1 0 4208 0 1 570
box -8 -3 16 105
use FILL  FILL_10158
timestamp 1680363874
transform 1 0 4216 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8045
timestamp 1680363874
transform 1 0 4236 0 1 575
box -3 -3 3 3
use FILL  FILL_10160
timestamp 1680363874
transform 1 0 4224 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_561
timestamp 1680363874
transform 1 0 4232 0 1 570
box -8 -3 104 105
use INVX2  INVX2_642
timestamp 1680363874
transform 1 0 4328 0 1 570
box -9 -3 26 105
use FILL  FILL_10162
timestamp 1680363874
transform 1 0 4344 0 1 570
box -8 -3 16 105
use FILL  FILL_10173
timestamp 1680363874
transform 1 0 4352 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_369
timestamp 1680363874
transform 1 0 4360 0 1 570
box -8 -3 46 105
use FILL  FILL_10175
timestamp 1680363874
transform 1 0 4400 0 1 570
box -8 -3 16 105
use FILL  FILL_10176
timestamp 1680363874
transform 1 0 4408 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_562
timestamp 1680363874
transform 1 0 4416 0 1 570
box -8 -3 104 105
use FILL  FILL_10177
timestamp 1680363874
transform 1 0 4512 0 1 570
box -8 -3 16 105
use FILL  FILL_10191
timestamp 1680363874
transform 1 0 4520 0 1 570
box -8 -3 16 105
use FILL  FILL_10192
timestamp 1680363874
transform 1 0 4528 0 1 570
box -8 -3 16 105
use FILL  FILL_10193
timestamp 1680363874
transform 1 0 4536 0 1 570
box -8 -3 16 105
use INVX2  INVX2_645
timestamp 1680363874
transform 1 0 4544 0 1 570
box -9 -3 26 105
use FILL  FILL_10194
timestamp 1680363874
transform 1 0 4560 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8046
timestamp 1680363874
transform 1 0 4580 0 1 575
box -3 -3 3 3
use FILL  FILL_10195
timestamp 1680363874
transform 1 0 4568 0 1 570
box -8 -3 16 105
use FILL  FILL_10196
timestamp 1680363874
transform 1 0 4576 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_370
timestamp 1680363874
transform 1 0 4584 0 1 570
box -8 -3 46 105
use FILL  FILL_10197
timestamp 1680363874
transform 1 0 4624 0 1 570
box -8 -3 16 105
use FILL  FILL_10200
timestamp 1680363874
transform 1 0 4632 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_371
timestamp 1680363874
transform 1 0 4640 0 1 570
box -8 -3 46 105
use INVX2  INVX2_646
timestamp 1680363874
transform 1 0 4680 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_564
timestamp 1680363874
transform -1 0 4792 0 1 570
box -8 -3 104 105
use FILL  FILL_10202
timestamp 1680363874
transform 1 0 4792 0 1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_83
timestamp 1680363874
transform 1 0 4827 0 1 570
box -10 -3 10 3
use M2_M1  M2_M1_9134
timestamp 1680363874
transform 1 0 68 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9018
timestamp 1680363874
transform 1 0 108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8197
timestamp 1680363874
transform 1 0 108 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9142
timestamp 1680363874
transform 1 0 116 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_8911
timestamp 1680363874
transform 1 0 140 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8914
timestamp 1680363874
transform 1 0 132 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8217
timestamp 1680363874
transform 1 0 124 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9135
timestamp 1680363874
transform 1 0 140 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8218
timestamp 1680363874
transform 1 0 148 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8912
timestamp 1680363874
transform 1 0 164 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_8047
timestamp 1680363874
transform 1 0 204 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8915
timestamp 1680363874
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9019
timestamp 1680363874
transform 1 0 180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9020
timestamp 1680363874
transform 1 0 196 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8159
timestamp 1680363874
transform 1 0 180 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9136
timestamp 1680363874
transform 1 0 188 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8198
timestamp 1680363874
transform 1 0 196 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8048
timestamp 1680363874
transform 1 0 244 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8078
timestamp 1680363874
transform 1 0 244 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8916
timestamp 1680363874
transform 1 0 228 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8113
timestamp 1680363874
transform 1 0 236 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8917
timestamp 1680363874
transform 1 0 252 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8114
timestamp 1680363874
transform 1 0 276 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9021
timestamp 1680363874
transform 1 0 236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9022
timestamp 1680363874
transform 1 0 244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9023
timestamp 1680363874
transform 1 0 260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9024
timestamp 1680363874
transform 1 0 276 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8160
timestamp 1680363874
transform 1 0 260 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8060
timestamp 1680363874
transform 1 0 292 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8918
timestamp 1680363874
transform 1 0 292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8919
timestamp 1680363874
transform 1 0 300 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8061
timestamp 1680363874
transform 1 0 332 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8079
timestamp 1680363874
transform 1 0 324 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8920
timestamp 1680363874
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8921
timestamp 1680363874
transform 1 0 332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9025
timestamp 1680363874
transform 1 0 308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9137
timestamp 1680363874
transform 1 0 324 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8161
timestamp 1680363874
transform 1 0 332 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8080
timestamp 1680363874
transform 1 0 364 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8922
timestamp 1680363874
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8923
timestamp 1680363874
transform 1 0 380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9026
timestamp 1680363874
transform 1 0 356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9027
timestamp 1680363874
transform 1 0 372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9028
timestamp 1680363874
transform 1 0 396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8162
timestamp 1680363874
transform 1 0 396 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8049
timestamp 1680363874
transform 1 0 524 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8081
timestamp 1680363874
transform 1 0 468 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8924
timestamp 1680363874
transform 1 0 516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9029
timestamp 1680363874
transform 1 0 468 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8138
timestamp 1680363874
transform 1 0 476 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8925
timestamp 1680363874
transform 1 0 532 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8139
timestamp 1680363874
transform 1 0 532 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8926
timestamp 1680363874
transform 1 0 588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9030
timestamp 1680363874
transform 1 0 588 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8163
timestamp 1680363874
transform 1 0 588 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8927
timestamp 1680363874
transform 1 0 604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8928
timestamp 1680363874
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9031
timestamp 1680363874
transform 1 0 596 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8140
timestamp 1680363874
transform 1 0 604 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9032
timestamp 1680363874
transform 1 0 612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8164
timestamp 1680363874
transform 1 0 612 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8929
timestamp 1680363874
transform 1 0 644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9033
timestamp 1680363874
transform 1 0 652 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8199
timestamp 1680363874
transform 1 0 652 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8229
timestamp 1680363874
transform 1 0 644 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8050
timestamp 1680363874
transform 1 0 668 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8082
timestamp 1680363874
transform 1 0 716 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8930
timestamp 1680363874
transform 1 0 668 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8141
timestamp 1680363874
transform 1 0 708 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8115
timestamp 1680363874
transform 1 0 756 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8931
timestamp 1680363874
transform 1 0 764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9034
timestamp 1680363874
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9035
timestamp 1680363874
transform 1 0 748 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9036
timestamp 1680363874
transform 1 0 756 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8200
timestamp 1680363874
transform 1 0 692 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8219
timestamp 1680363874
transform 1 0 684 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8220
timestamp 1680363874
transform 1 0 700 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8230
timestamp 1680363874
transform 1 0 676 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8083
timestamp 1680363874
transform 1 0 804 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8932
timestamp 1680363874
transform 1 0 804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8933
timestamp 1680363874
transform 1 0 820 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8142
timestamp 1680363874
transform 1 0 804 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9037
timestamp 1680363874
transform 1 0 812 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8165
timestamp 1680363874
transform 1 0 812 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8143
timestamp 1680363874
transform 1 0 828 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8201
timestamp 1680363874
transform 1 0 820 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8051
timestamp 1680363874
transform 1 0 860 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8934
timestamp 1680363874
transform 1 0 884 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8116
timestamp 1680363874
transform 1 0 892 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9038
timestamp 1680363874
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9039
timestamp 1680363874
transform 1 0 892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9040
timestamp 1680363874
transform 1 0 900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8166
timestamp 1680363874
transform 1 0 876 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8167
timestamp 1680363874
transform 1 0 900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8221
timestamp 1680363874
transform 1 0 892 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8935
timestamp 1680363874
transform 1 0 916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8936
timestamp 1680363874
transform 1 0 940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9138
timestamp 1680363874
transform 1 0 948 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9041
timestamp 1680363874
transform 1 0 972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9042
timestamp 1680363874
transform 1 0 996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9139
timestamp 1680363874
transform 1 0 1012 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9143
timestamp 1680363874
transform 1 0 1004 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_8117
timestamp 1680363874
transform 1 0 1036 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8222
timestamp 1680363874
transform 1 0 1044 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8937
timestamp 1680363874
transform 1 0 1052 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8231
timestamp 1680363874
transform 1 0 1060 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8118
timestamp 1680363874
transform 1 0 1076 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8084
timestamp 1680363874
transform 1 0 1092 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9043
timestamp 1680363874
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8052
timestamp 1680363874
transform 1 0 1132 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8085
timestamp 1680363874
transform 1 0 1124 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8086
timestamp 1680363874
transform 1 0 1172 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8938
timestamp 1680363874
transform 1 0 1124 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8144
timestamp 1680363874
transform 1 0 1124 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8145
timestamp 1680363874
transform 1 0 1148 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9044
timestamp 1680363874
transform 1 0 1172 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8202
timestamp 1680363874
transform 1 0 1204 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8232
timestamp 1680363874
transform 1 0 1180 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8062
timestamp 1680363874
transform 1 0 1244 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8087
timestamp 1680363874
transform 1 0 1260 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8119
timestamp 1680363874
transform 1 0 1236 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8939
timestamp 1680363874
transform 1 0 1244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8940
timestamp 1680363874
transform 1 0 1260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9045
timestamp 1680363874
transform 1 0 1236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9046
timestamp 1680363874
transform 1 0 1252 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8146
timestamp 1680363874
transform 1 0 1260 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9047
timestamp 1680363874
transform 1 0 1276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9048
timestamp 1680363874
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8941
timestamp 1680363874
transform 1 0 1300 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8063
timestamp 1680363874
transform 1 0 1316 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8942
timestamp 1680363874
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8943
timestamp 1680363874
transform 1 0 1340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8944
timestamp 1680363874
transform 1 0 1356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9049
timestamp 1680363874
transform 1 0 1332 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8147
timestamp 1680363874
transform 1 0 1340 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9050
timestamp 1680363874
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8168
timestamp 1680363874
transform 1 0 1324 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8088
timestamp 1680363874
transform 1 0 1388 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8945
timestamp 1680363874
transform 1 0 1372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8946
timestamp 1680363874
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9051
timestamp 1680363874
transform 1 0 1364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9052
timestamp 1680363874
transform 1 0 1380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9053
timestamp 1680363874
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8169
timestamp 1680363874
transform 1 0 1364 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8170
timestamp 1680363874
transform 1 0 1380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8203
timestamp 1680363874
transform 1 0 1348 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8204
timestamp 1680363874
transform 1 0 1372 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8947
timestamp 1680363874
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8223
timestamp 1680363874
transform 1 0 1412 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8064
timestamp 1680363874
transform 1 0 1436 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8065
timestamp 1680363874
transform 1 0 1500 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8089
timestamp 1680363874
transform 1 0 1460 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8948
timestamp 1680363874
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8148
timestamp 1680363874
transform 1 0 1436 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8949
timestamp 1680363874
transform 1 0 1524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9054
timestamp 1680363874
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9055
timestamp 1680363874
transform 1 0 1516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8171
timestamp 1680363874
transform 1 0 1524 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8053
timestamp 1680363874
transform 1 0 1596 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8120
timestamp 1680363874
transform 1 0 1620 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9056
timestamp 1680363874
transform 1 0 1572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9057
timestamp 1680363874
transform 1 0 1588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9058
timestamp 1680363874
transform 1 0 1604 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8172
timestamp 1680363874
transform 1 0 1572 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8149
timestamp 1680363874
transform 1 0 1612 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8090
timestamp 1680363874
transform 1 0 1644 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8950
timestamp 1680363874
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8951
timestamp 1680363874
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8952
timestamp 1680363874
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8066
timestamp 1680363874
transform 1 0 1692 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8091
timestamp 1680363874
transform 1 0 1684 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9059
timestamp 1680363874
transform 1 0 1660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9060
timestamp 1680363874
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9061
timestamp 1680363874
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8173
timestamp 1680363874
transform 1 0 1676 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8121
timestamp 1680363874
transform 1 0 1748 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8953
timestamp 1680363874
transform 1 0 1764 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8054
timestamp 1680363874
transform 1 0 1788 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8122
timestamp 1680363874
transform 1 0 1788 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8954
timestamp 1680363874
transform 1 0 1796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8955
timestamp 1680363874
transform 1 0 1812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9062
timestamp 1680363874
transform 1 0 1780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9063
timestamp 1680363874
transform 1 0 1788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9064
timestamp 1680363874
transform 1 0 1804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9065
timestamp 1680363874
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8174
timestamp 1680363874
transform 1 0 1780 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8175
timestamp 1680363874
transform 1 0 1828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8205
timestamp 1680363874
transform 1 0 1820 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8956
timestamp 1680363874
transform 1 0 1852 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8176
timestamp 1680363874
transform 1 0 1852 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8224
timestamp 1680363874
transform 1 0 1852 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8067
timestamp 1680363874
transform 1 0 1884 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9066
timestamp 1680363874
transform 1 0 1884 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8206
timestamp 1680363874
transform 1 0 1908 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9067
timestamp 1680363874
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8055
timestamp 1680363874
transform 1 0 1956 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8957
timestamp 1680363874
transform 1 0 1948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8958
timestamp 1680363874
transform 1 0 1964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8959
timestamp 1680363874
transform 1 0 1980 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8150
timestamp 1680363874
transform 1 0 1948 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9068
timestamp 1680363874
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8207
timestamp 1680363874
transform 1 0 1948 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8056
timestamp 1680363874
transform 1 0 2004 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8092
timestamp 1680363874
transform 1 0 2020 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9069
timestamp 1680363874
transform 1 0 1996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9070
timestamp 1680363874
transform 1 0 2004 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8151
timestamp 1680363874
transform 1 0 2012 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8208
timestamp 1680363874
transform 1 0 2004 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8093
timestamp 1680363874
transform 1 0 2068 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8960
timestamp 1680363874
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8961
timestamp 1680363874
transform 1 0 2060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8962
timestamp 1680363874
transform 1 0 2068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9071
timestamp 1680363874
transform 1 0 2052 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9072
timestamp 1680363874
transform 1 0 2068 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8152
timestamp 1680363874
transform 1 0 2092 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8068
timestamp 1680363874
transform 1 0 2116 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8094
timestamp 1680363874
transform 1 0 2164 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8963
timestamp 1680363874
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9073
timestamp 1680363874
transform 1 0 2164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8123
timestamp 1680363874
transform 1 0 2212 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8095
timestamp 1680363874
transform 1 0 2252 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8964
timestamp 1680363874
transform 1 0 2236 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8124
timestamp 1680363874
transform 1 0 2244 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8965
timestamp 1680363874
transform 1 0 2252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9074
timestamp 1680363874
transform 1 0 2228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9075
timestamp 1680363874
transform 1 0 2244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9076
timestamp 1680363874
transform 1 0 2260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8966
timestamp 1680363874
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9077
timestamp 1680363874
transform 1 0 2284 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8177
timestamp 1680363874
transform 1 0 2292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8225
timestamp 1680363874
transform 1 0 2284 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8057
timestamp 1680363874
transform 1 0 2324 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_9078
timestamp 1680363874
transform 1 0 2316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8967
timestamp 1680363874
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9140
timestamp 1680363874
transform 1 0 2348 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8968
timestamp 1680363874
transform 1 0 2364 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8125
timestamp 1680363874
transform 1 0 2412 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9079
timestamp 1680363874
transform 1 0 2404 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8069
timestamp 1680363874
transform 1 0 2444 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9080
timestamp 1680363874
transform 1 0 2500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8969
timestamp 1680363874
transform 1 0 2548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8970
timestamp 1680363874
transform 1 0 2572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9081
timestamp 1680363874
transform 1 0 2564 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8058
timestamp 1680363874
transform 1 0 2588 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_9082
timestamp 1680363874
transform 1 0 2588 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8096
timestamp 1680363874
transform 1 0 2628 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8971
timestamp 1680363874
transform 1 0 2612 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8972
timestamp 1680363874
transform 1 0 2628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9083
timestamp 1680363874
transform 1 0 2620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9084
timestamp 1680363874
transform 1 0 2636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8178
timestamp 1680363874
transform 1 0 2636 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8973
timestamp 1680363874
transform 1 0 2660 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8059
timestamp 1680363874
transform 1 0 2684 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8070
timestamp 1680363874
transform 1 0 2676 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8071
timestamp 1680363874
transform 1 0 2708 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8097
timestamp 1680363874
transform 1 0 2700 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8974
timestamp 1680363874
transform 1 0 2676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9085
timestamp 1680363874
transform 1 0 2700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8209
timestamp 1680363874
transform 1 0 2772 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8072
timestamp 1680363874
transform 1 0 2812 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8098
timestamp 1680363874
transform 1 0 2804 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8913
timestamp 1680363874
transform 1 0 2812 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_9086
timestamp 1680363874
transform 1 0 2796 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8179
timestamp 1680363874
transform 1 0 2796 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8099
timestamp 1680363874
transform 1 0 2820 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8975
timestamp 1680363874
transform 1 0 2812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8976
timestamp 1680363874
transform 1 0 2836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9087
timestamp 1680363874
transform 1 0 2828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9088
timestamp 1680363874
transform 1 0 2860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9141
timestamp 1680363874
transform 1 0 2836 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8180
timestamp 1680363874
transform 1 0 2844 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8181
timestamp 1680363874
transform 1 0 2860 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9144
timestamp 1680363874
transform 1 0 2892 0 1 485
box -2 -2 2 2
use M2_M1  M2_M1_8977
timestamp 1680363874
transform 1 0 2932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9145
timestamp 1680363874
transform 1 0 2924 0 1 485
box -2 -2 2 2
use M2_M1  M2_M1_8978
timestamp 1680363874
transform 1 0 2956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9089
timestamp 1680363874
transform 1 0 3036 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8073
timestamp 1680363874
transform 1 0 3068 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8979
timestamp 1680363874
transform 1 0 3052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8980
timestamp 1680363874
transform 1 0 3068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9090
timestamp 1680363874
transform 1 0 3060 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8182
timestamp 1680363874
transform 1 0 3060 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8126
timestamp 1680363874
transform 1 0 3108 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8100
timestamp 1680363874
transform 1 0 3156 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8981
timestamp 1680363874
transform 1 0 3116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8982
timestamp 1680363874
transform 1 0 3124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8983
timestamp 1680363874
transform 1 0 3140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9091
timestamp 1680363874
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8153
timestamp 1680363874
transform 1 0 3116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8127
timestamp 1680363874
transform 1 0 3148 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8984
timestamp 1680363874
transform 1 0 3156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8985
timestamp 1680363874
transform 1 0 3164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9092
timestamp 1680363874
transform 1 0 3132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9093
timestamp 1680363874
transform 1 0 3148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9094
timestamp 1680363874
transform 1 0 3156 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8183
timestamp 1680363874
transform 1 0 3132 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8986
timestamp 1680363874
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8987
timestamp 1680363874
transform 1 0 3228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9095
timestamp 1680363874
transform 1 0 3196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9096
timestamp 1680363874
transform 1 0 3212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8988
timestamp 1680363874
transform 1 0 3268 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8128
timestamp 1680363874
transform 1 0 3300 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8989
timestamp 1680363874
transform 1 0 3380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9097
timestamp 1680363874
transform 1 0 3292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9098
timestamp 1680363874
transform 1 0 3300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9099
timestamp 1680363874
transform 1 0 3332 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8184
timestamp 1680363874
transform 1 0 3292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8185
timestamp 1680363874
transform 1 0 3332 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8233
timestamp 1680363874
transform 1 0 3380 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8154
timestamp 1680363874
transform 1 0 3404 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8101
timestamp 1680363874
transform 1 0 3420 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8102
timestamp 1680363874
transform 1 0 3460 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8990
timestamp 1680363874
transform 1 0 3420 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8129
timestamp 1680363874
transform 1 0 3484 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8991
timestamp 1680363874
transform 1 0 3508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9100
timestamp 1680363874
transform 1 0 3468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9101
timestamp 1680363874
transform 1 0 3500 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8130
timestamp 1680363874
transform 1 0 3516 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9102
timestamp 1680363874
transform 1 0 3516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8992
timestamp 1680363874
transform 1 0 3540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9103
timestamp 1680363874
transform 1 0 3548 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8210
timestamp 1680363874
transform 1 0 3548 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8234
timestamp 1680363874
transform 1 0 3532 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8103
timestamp 1680363874
transform 1 0 3572 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8104
timestamp 1680363874
transform 1 0 3596 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8993
timestamp 1680363874
transform 1 0 3572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8994
timestamp 1680363874
transform 1 0 3580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8995
timestamp 1680363874
transform 1 0 3596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8996
timestamp 1680363874
transform 1 0 3604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9104
timestamp 1680363874
transform 1 0 3572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9105
timestamp 1680363874
transform 1 0 3588 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8226
timestamp 1680363874
transform 1 0 3572 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9106
timestamp 1680363874
transform 1 0 3612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8105
timestamp 1680363874
transform 1 0 3652 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8131
timestamp 1680363874
transform 1 0 3652 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8132
timestamp 1680363874
transform 1 0 3668 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8997
timestamp 1680363874
transform 1 0 3716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9107
timestamp 1680363874
transform 1 0 3628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9108
timestamp 1680363874
transform 1 0 3636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9109
timestamp 1680363874
transform 1 0 3668 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8155
timestamp 1680363874
transform 1 0 3676 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8186
timestamp 1680363874
transform 1 0 3628 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8187
timestamp 1680363874
transform 1 0 3668 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8211
timestamp 1680363874
transform 1 0 3684 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8227
timestamp 1680363874
transform 1 0 3628 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8228
timestamp 1680363874
transform 1 0 3652 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9110
timestamp 1680363874
transform 1 0 3788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8212
timestamp 1680363874
transform 1 0 3804 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8188
timestamp 1680363874
transform 1 0 3820 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8998
timestamp 1680363874
transform 1 0 3860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8999
timestamp 1680363874
transform 1 0 3868 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8156
timestamp 1680363874
transform 1 0 3852 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9111
timestamp 1680363874
transform 1 0 3860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9112
timestamp 1680363874
transform 1 0 3876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9113
timestamp 1680363874
transform 1 0 3892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9114
timestamp 1680363874
transform 1 0 3900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8189
timestamp 1680363874
transform 1 0 3868 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8213
timestamp 1680363874
transform 1 0 3860 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8214
timestamp 1680363874
transform 1 0 3900 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8106
timestamp 1680363874
transform 1 0 3916 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9000
timestamp 1680363874
transform 1 0 3916 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8107
timestamp 1680363874
transform 1 0 3956 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9001
timestamp 1680363874
transform 1 0 3940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9002
timestamp 1680363874
transform 1 0 3956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9115
timestamp 1680363874
transform 1 0 3948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9003
timestamp 1680363874
transform 1 0 3988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9116
timestamp 1680363874
transform 1 0 3980 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8133
timestamp 1680363874
transform 1 0 4020 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9117
timestamp 1680363874
transform 1 0 4028 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8190
timestamp 1680363874
transform 1 0 4028 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9004
timestamp 1680363874
transform 1 0 4060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9118
timestamp 1680363874
transform 1 0 4092 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8108
timestamp 1680363874
transform 1 0 4148 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9005
timestamp 1680363874
transform 1 0 4140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9006
timestamp 1680363874
transform 1 0 4156 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8134
timestamp 1680363874
transform 1 0 4164 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9007
timestamp 1680363874
transform 1 0 4172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9119
timestamp 1680363874
transform 1 0 4148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9120
timestamp 1680363874
transform 1 0 4164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9121
timestamp 1680363874
transform 1 0 4180 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8109
timestamp 1680363874
transform 1 0 4196 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9008
timestamp 1680363874
transform 1 0 4196 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8191
timestamp 1680363874
transform 1 0 4180 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9122
timestamp 1680363874
transform 1 0 4204 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8192
timestamp 1680363874
transform 1 0 4204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8135
timestamp 1680363874
transform 1 0 4236 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8074
timestamp 1680363874
transform 1 0 4284 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9009
timestamp 1680363874
transform 1 0 4284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9123
timestamp 1680363874
transform 1 0 4292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8110
timestamp 1680363874
transform 1 0 4324 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8075
timestamp 1680363874
transform 1 0 4340 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8076
timestamp 1680363874
transform 1 0 4388 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8111
timestamp 1680363874
transform 1 0 4380 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8215
timestamp 1680363874
transform 1 0 4372 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9010
timestamp 1680363874
transform 1 0 4388 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8136
timestamp 1680363874
transform 1 0 4396 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8112
timestamp 1680363874
transform 1 0 4428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9011
timestamp 1680363874
transform 1 0 4404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9012
timestamp 1680363874
transform 1 0 4420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9013
timestamp 1680363874
transform 1 0 4428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9124
timestamp 1680363874
transform 1 0 4388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9125
timestamp 1680363874
transform 1 0 4396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9126
timestamp 1680363874
transform 1 0 4412 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8157
timestamp 1680363874
transform 1 0 4420 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8077
timestamp 1680363874
transform 1 0 4468 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9127
timestamp 1680363874
transform 1 0 4508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9014
timestamp 1680363874
transform 1 0 4532 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8137
timestamp 1680363874
transform 1 0 4564 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9128
timestamp 1680363874
transform 1 0 4556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9129
timestamp 1680363874
transform 1 0 4612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9130
timestamp 1680363874
transform 1 0 4620 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8193
timestamp 1680363874
transform 1 0 4612 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8216
timestamp 1680363874
transform 1 0 4620 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8194
timestamp 1680363874
transform 1 0 4636 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9015
timestamp 1680363874
transform 1 0 4652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9016
timestamp 1680363874
transform 1 0 4668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9017
timestamp 1680363874
transform 1 0 4676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9131
timestamp 1680363874
transform 1 0 4660 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8158
timestamp 1680363874
transform 1 0 4668 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9132
timestamp 1680363874
transform 1 0 4684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8195
timestamp 1680363874
transform 1 0 4676 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8196
timestamp 1680363874
transform 1 0 4716 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9133
timestamp 1680363874
transform 1 0 4748 0 1 525
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_84
timestamp 1680363874
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_9781
timestamp 1680363874
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_9782
timestamp 1680363874
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_9783
timestamp 1680363874
transform 1 0 88 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_71
timestamp 1680363874
transform 1 0 96 0 -1 570
box -8 -3 40 105
use FILL  FILL_9784
timestamp 1680363874
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_9785
timestamp 1680363874
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_9786
timestamp 1680363874
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_9787
timestamp 1680363874
transform 1 0 152 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_112
timestamp 1680363874
transform 1 0 160 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1680363874
transform -1 0 208 0 -1 570
box -8 -3 32 105
use FILL  FILL_9788
timestamp 1680363874
transform 1 0 208 0 -1 570
box -8 -3 16 105
use FILL  FILL_9789
timestamp 1680363874
transform 1 0 216 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_609
timestamp 1680363874
transform 1 0 224 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_352
timestamp 1680363874
transform 1 0 240 0 -1 570
box -8 -3 46 105
use FILL  FILL_9790
timestamp 1680363874
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_9791
timestamp 1680363874
transform 1 0 288 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_167
timestamp 1680363874
transform 1 0 296 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_610
timestamp 1680363874
transform 1 0 328 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_378
timestamp 1680363874
transform 1 0 344 0 -1 570
box -8 -3 46 105
use FILL  FILL_9792
timestamp 1680363874
transform 1 0 384 0 -1 570
box -8 -3 16 105
use FILL  FILL_9793
timestamp 1680363874
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_9794
timestamp 1680363874
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_9795
timestamp 1680363874
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_9796
timestamp 1680363874
transform 1 0 416 0 -1 570
box -8 -3 16 105
use FILL  FILL_9797
timestamp 1680363874
transform 1 0 424 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_543
timestamp 1680363874
transform -1 0 528 0 -1 570
box -8 -3 104 105
use FILL  FILL_9798
timestamp 1680363874
transform 1 0 528 0 -1 570
box -8 -3 16 105
use FILL  FILL_9799
timestamp 1680363874
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_9800
timestamp 1680363874
transform 1 0 544 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_611
timestamp 1680363874
transform 1 0 552 0 -1 570
box -9 -3 26 105
use FILL  FILL_9801
timestamp 1680363874
transform 1 0 568 0 -1 570
box -8 -3 16 105
use FILL  FILL_9802
timestamp 1680363874
transform 1 0 576 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_612
timestamp 1680363874
transform 1 0 584 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_379
timestamp 1680363874
transform -1 0 640 0 -1 570
box -8 -3 46 105
use FILL  FILL_9803
timestamp 1680363874
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_9812
timestamp 1680363874
transform 1 0 648 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_544
timestamp 1680363874
transform 1 0 656 0 -1 570
box -8 -3 104 105
use FILL  FILL_9813
timestamp 1680363874
transform 1 0 752 0 -1 570
box -8 -3 16 105
use FILL  FILL_9814
timestamp 1680363874
transform 1 0 760 0 -1 570
box -8 -3 16 105
use FILL  FILL_9816
timestamp 1680363874
transform 1 0 768 0 -1 570
box -8 -3 16 105
use FILL  FILL_9818
timestamp 1680363874
transform 1 0 776 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_381
timestamp 1680363874
transform 1 0 784 0 -1 570
box -8 -3 46 105
use FILL  FILL_9825
timestamp 1680363874
transform 1 0 824 0 -1 570
box -8 -3 16 105
use FILL  FILL_9827
timestamp 1680363874
transform 1 0 832 0 -1 570
box -8 -3 16 105
use FILL  FILL_9829
timestamp 1680363874
transform 1 0 840 0 -1 570
box -8 -3 16 105
use FILL  FILL_9831
timestamp 1680363874
transform 1 0 848 0 -1 570
box -8 -3 16 105
use FILL  FILL_9832
timestamp 1680363874
transform 1 0 856 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_382
timestamp 1680363874
transform -1 0 904 0 -1 570
box -8 -3 46 105
use FILL  FILL_9833
timestamp 1680363874
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_9834
timestamp 1680363874
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_9835
timestamp 1680363874
transform 1 0 920 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_614
timestamp 1680363874
transform -1 0 944 0 -1 570
box -9 -3 26 105
use FILL  FILL_9836
timestamp 1680363874
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_9838
timestamp 1680363874
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_9840
timestamp 1680363874
transform 1 0 960 0 -1 570
box -8 -3 16 105
use FILL  FILL_9842
timestamp 1680363874
transform 1 0 968 0 -1 570
box -8 -3 16 105
use FILL  FILL_9844
timestamp 1680363874
transform 1 0 976 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_72
timestamp 1680363874
transform 1 0 984 0 -1 570
box -8 -3 40 105
use FILL  FILL_9850
timestamp 1680363874
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_9852
timestamp 1680363874
transform 1 0 1024 0 -1 570
box -8 -3 16 105
use FILL  FILL_9854
timestamp 1680363874
transform 1 0 1032 0 -1 570
box -8 -3 16 105
use FILL  FILL_9874
timestamp 1680363874
transform 1 0 1040 0 -1 570
box -8 -3 16 105
use FILL  FILL_9875
timestamp 1680363874
transform 1 0 1048 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_615
timestamp 1680363874
transform 1 0 1056 0 -1 570
box -9 -3 26 105
use FILL  FILL_9876
timestamp 1680363874
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_9877
timestamp 1680363874
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_9878
timestamp 1680363874
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_9879
timestamp 1680363874
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_9880
timestamp 1680363874
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_547
timestamp 1680363874
transform 1 0 1112 0 -1 570
box -8 -3 104 105
use FILL  FILL_9881
timestamp 1680363874
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_9882
timestamp 1680363874
transform 1 0 1216 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_616
timestamp 1680363874
transform 1 0 1224 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_383
timestamp 1680363874
transform -1 0 1280 0 -1 570
box -8 -3 46 105
use FILL  FILL_9883
timestamp 1680363874
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_9884
timestamp 1680363874
transform 1 0 1288 0 -1 570
box -8 -3 16 105
use FILL  FILL_9885
timestamp 1680363874
transform 1 0 1296 0 -1 570
box -8 -3 16 105
use FILL  FILL_9886
timestamp 1680363874
transform 1 0 1304 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_354
timestamp 1680363874
transform -1 0 1352 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_617
timestamp 1680363874
transform 1 0 1352 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_384
timestamp 1680363874
transform -1 0 1408 0 -1 570
box -8 -3 46 105
use FILL  FILL_9887
timestamp 1680363874
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_9889
timestamp 1680363874
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_548
timestamp 1680363874
transform 1 0 1424 0 -1 570
box -8 -3 104 105
use FILL  FILL_9895
timestamp 1680363874
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_9896
timestamp 1680363874
transform 1 0 1528 0 -1 570
box -8 -3 16 105
use FILL  FILL_9898
timestamp 1680363874
transform 1 0 1536 0 -1 570
box -8 -3 16 105
use FILL  FILL_9900
timestamp 1680363874
transform 1 0 1544 0 -1 570
box -8 -3 16 105
use FILL  FILL_9902
timestamp 1680363874
transform 1 0 1552 0 -1 570
box -8 -3 16 105
use FILL  FILL_9906
timestamp 1680363874
transform 1 0 1560 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_355
timestamp 1680363874
transform -1 0 1608 0 -1 570
box -8 -3 46 105
use FILL  FILL_9907
timestamp 1680363874
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_9908
timestamp 1680363874
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_9909
timestamp 1680363874
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_9914
timestamp 1680363874
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_356
timestamp 1680363874
transform 1 0 1640 0 -1 570
box -8 -3 46 105
use FILL  FILL_9915
timestamp 1680363874
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_9917
timestamp 1680363874
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_9919
timestamp 1680363874
transform 1 0 1696 0 -1 570
box -8 -3 16 105
use FILL  FILL_9920
timestamp 1680363874
transform 1 0 1704 0 -1 570
box -8 -3 16 105
use FILL  FILL_9921
timestamp 1680363874
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_9922
timestamp 1680363874
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_621
timestamp 1680363874
transform -1 0 1744 0 -1 570
box -9 -3 26 105
use FILL  FILL_9923
timestamp 1680363874
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_9924
timestamp 1680363874
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_9930
timestamp 1680363874
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_9931
timestamp 1680363874
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_9932
timestamp 1680363874
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_357
timestamp 1680363874
transform 1 0 1784 0 -1 570
box -8 -3 46 105
use FILL  FILL_9933
timestamp 1680363874
transform 1 0 1824 0 -1 570
box -8 -3 16 105
use FILL  FILL_9934
timestamp 1680363874
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_9935
timestamp 1680363874
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use FILL  FILL_9936
timestamp 1680363874
transform 1 0 1848 0 -1 570
box -8 -3 16 105
use FILL  FILL_9937
timestamp 1680363874
transform 1 0 1856 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_105
timestamp 1680363874
transform -1 0 1888 0 -1 570
box -5 -3 28 105
use FILL  FILL_9938
timestamp 1680363874
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_9939
timestamp 1680363874
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_106
timestamp 1680363874
transform -1 0 1928 0 -1 570
box -5 -3 28 105
use FILL  FILL_9940
timestamp 1680363874
transform 1 0 1928 0 -1 570
box -8 -3 16 105
use FILL  FILL_9941
timestamp 1680363874
transform 1 0 1936 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_387
timestamp 1680363874
transform -1 0 1984 0 -1 570
box -8 -3 46 105
use FILL  FILL_9942
timestamp 1680363874
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_9944
timestamp 1680363874
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_9945
timestamp 1680363874
transform 1 0 2000 0 -1 570
box -8 -3 16 105
use FILL  FILL_9946
timestamp 1680363874
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_9951
timestamp 1680363874
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_388
timestamp 1680363874
transform 1 0 2024 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_623
timestamp 1680363874
transform 1 0 2064 0 -1 570
box -9 -3 26 105
use FILL  FILL_9952
timestamp 1680363874
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_9954
timestamp 1680363874
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use FILL  FILL_9962
timestamp 1680363874
transform 1 0 2096 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_551
timestamp 1680363874
transform 1 0 2104 0 -1 570
box -8 -3 104 105
use FILL  FILL_9963
timestamp 1680363874
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_9965
timestamp 1680363874
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_624
timestamp 1680363874
transform 1 0 2216 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_389
timestamp 1680363874
transform -1 0 2272 0 -1 570
box -8 -3 46 105
use FILL  FILL_9970
timestamp 1680363874
transform 1 0 2272 0 -1 570
box -8 -3 16 105
use FILL  FILL_9972
timestamp 1680363874
transform 1 0 2280 0 -1 570
box -8 -3 16 105
use FILL  FILL_9974
timestamp 1680363874
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_9979
timestamp 1680363874
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_9980
timestamp 1680363874
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_172
timestamp 1680363874
transform 1 0 2312 0 -1 570
box -8 -3 34 105
use FILL  FILL_9981
timestamp 1680363874
transform 1 0 2344 0 -1 570
box -8 -3 16 105
use FILL  FILL_9982
timestamp 1680363874
transform 1 0 2352 0 -1 570
box -8 -3 16 105
use FILL  FILL_9983
timestamp 1680363874
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_9984
timestamp 1680363874
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9985
timestamp 1680363874
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use FILL  FILL_9986
timestamp 1680363874
transform 1 0 2384 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_625
timestamp 1680363874
transform 1 0 2392 0 -1 570
box -9 -3 26 105
use FILL  FILL_9987
timestamp 1680363874
transform 1 0 2408 0 -1 570
box -8 -3 16 105
use FILL  FILL_9988
timestamp 1680363874
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_9989
timestamp 1680363874
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_9990
timestamp 1680363874
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_9991
timestamp 1680363874
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use FILL  FILL_9992
timestamp 1680363874
transform 1 0 2448 0 -1 570
box -8 -3 16 105
use FILL  FILL_9994
timestamp 1680363874
transform 1 0 2456 0 -1 570
box -8 -3 16 105
use FILL  FILL_9996
timestamp 1680363874
transform 1 0 2464 0 -1 570
box -8 -3 16 105
use FILL  FILL_9998
timestamp 1680363874
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_9999
timestamp 1680363874
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_10000
timestamp 1680363874
transform 1 0 2488 0 -1 570
box -8 -3 16 105
use FILL  FILL_10001
timestamp 1680363874
transform 1 0 2496 0 -1 570
box -8 -3 16 105
use FILL  FILL_10002
timestamp 1680363874
transform 1 0 2504 0 -1 570
box -8 -3 16 105
use FILL  FILL_10003
timestamp 1680363874
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_10005
timestamp 1680363874
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_10012
timestamp 1680363874
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_10013
timestamp 1680363874
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_627
timestamp 1680363874
transform 1 0 2544 0 -1 570
box -9 -3 26 105
use FILL  FILL_10014
timestamp 1680363874
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_109
timestamp 1680363874
transform -1 0 2592 0 -1 570
box -5 -3 28 105
use FILL  FILL_10015
timestamp 1680363874
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_10016
timestamp 1680363874
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_393
timestamp 1680363874
transform 1 0 2608 0 -1 570
box -8 -3 46 105
use FILL  FILL_10017
timestamp 1680363874
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_10018
timestamp 1680363874
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_553
timestamp 1680363874
transform 1 0 2664 0 -1 570
box -8 -3 104 105
use FILL  FILL_10024
timestamp 1680363874
transform 1 0 2760 0 -1 570
box -8 -3 16 105
use FILL  FILL_10025
timestamp 1680363874
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use FILL  FILL_10026
timestamp 1680363874
transform 1 0 2776 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_628
timestamp 1680363874
transform 1 0 2784 0 -1 570
box -9 -3 26 105
use FILL  FILL_10027
timestamp 1680363874
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_115
timestamp 1680363874
transform 1 0 2808 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_174
timestamp 1680363874
transform -1 0 2864 0 -1 570
box -8 -3 34 105
use FILL  FILL_10028
timestamp 1680363874
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_10031
timestamp 1680363874
transform 1 0 2872 0 -1 570
box -8 -3 16 105
use FILL  FILL_10032
timestamp 1680363874
transform 1 0 2880 0 -1 570
box -8 -3 16 105
use FILL  FILL_10033
timestamp 1680363874
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use FILL  FILL_10034
timestamp 1680363874
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_10035
timestamp 1680363874
transform 1 0 2904 0 -1 570
box -8 -3 16 105
use FILL  FILL_10036
timestamp 1680363874
transform 1 0 2912 0 -1 570
box -8 -3 16 105
use FILL  FILL_10037
timestamp 1680363874
transform 1 0 2920 0 -1 570
box -8 -3 16 105
use FILL  FILL_10038
timestamp 1680363874
transform 1 0 2928 0 -1 570
box -8 -3 16 105
use FILL  FILL_10039
timestamp 1680363874
transform 1 0 2936 0 -1 570
box -8 -3 16 105
use FILL  FILL_10040
timestamp 1680363874
transform 1 0 2944 0 -1 570
box -8 -3 16 105
use FILL  FILL_10041
timestamp 1680363874
transform 1 0 2952 0 -1 570
box -8 -3 16 105
use FILL  FILL_10042
timestamp 1680363874
transform 1 0 2960 0 -1 570
box -8 -3 16 105
use FILL  FILL_10043
timestamp 1680363874
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_10044
timestamp 1680363874
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_631
timestamp 1680363874
transform 1 0 2984 0 -1 570
box -9 -3 26 105
use FILL  FILL_10048
timestamp 1680363874
transform 1 0 3000 0 -1 570
box -8 -3 16 105
use FILL  FILL_10049
timestamp 1680363874
transform 1 0 3008 0 -1 570
box -8 -3 16 105
use FILL  FILL_10050
timestamp 1680363874
transform 1 0 3016 0 -1 570
box -8 -3 16 105
use FILL  FILL_10051
timestamp 1680363874
transform 1 0 3024 0 -1 570
box -8 -3 16 105
use FILL  FILL_10052
timestamp 1680363874
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_10053
timestamp 1680363874
transform 1 0 3040 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_394
timestamp 1680363874
transform -1 0 3088 0 -1 570
box -8 -3 46 105
use FILL  FILL_10054
timestamp 1680363874
transform 1 0 3088 0 -1 570
box -8 -3 16 105
use FILL  FILL_10055
timestamp 1680363874
transform 1 0 3096 0 -1 570
box -8 -3 16 105
use FILL  FILL_10057
timestamp 1680363874
transform 1 0 3104 0 -1 570
box -8 -3 16 105
use FILL  FILL_10061
timestamp 1680363874
transform 1 0 3112 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_396
timestamp 1680363874
transform -1 0 3160 0 -1 570
box -8 -3 46 105
use FILL  FILL_10062
timestamp 1680363874
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use FILL  FILL_10063
timestamp 1680363874
transform 1 0 3168 0 -1 570
box -8 -3 16 105
use FILL  FILL_10070
timestamp 1680363874
transform 1 0 3176 0 -1 570
box -8 -3 16 105
use FILL  FILL_10071
timestamp 1680363874
transform 1 0 3184 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_360
timestamp 1680363874
transform -1 0 3232 0 -1 570
box -8 -3 46 105
use FILL  FILL_10072
timestamp 1680363874
transform 1 0 3232 0 -1 570
box -8 -3 16 105
use FILL  FILL_10074
timestamp 1680363874
transform 1 0 3240 0 -1 570
box -8 -3 16 105
use FILL  FILL_10076
timestamp 1680363874
transform 1 0 3248 0 -1 570
box -8 -3 16 105
use FILL  FILL_10079
timestamp 1680363874
transform 1 0 3256 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_634
timestamp 1680363874
transform 1 0 3264 0 -1 570
box -9 -3 26 105
use FILL  FILL_10080
timestamp 1680363874
transform 1 0 3280 0 -1 570
box -8 -3 16 105
use FILL  FILL_10088
timestamp 1680363874
transform 1 0 3288 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_556
timestamp 1680363874
transform -1 0 3392 0 -1 570
box -8 -3 104 105
use FILL  FILL_10089
timestamp 1680363874
transform 1 0 3392 0 -1 570
box -8 -3 16 105
use FILL  FILL_10090
timestamp 1680363874
transform 1 0 3400 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_557
timestamp 1680363874
transform 1 0 3408 0 -1 570
box -8 -3 104 105
use FILL  FILL_10091
timestamp 1680363874
transform 1 0 3504 0 -1 570
box -8 -3 16 105
use FILL  FILL_10093
timestamp 1680363874
transform 1 0 3512 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_397
timestamp 1680363874
transform 1 0 3520 0 -1 570
box -8 -3 46 105
use FILL  FILL_10095
timestamp 1680363874
transform 1 0 3560 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_364
timestamp 1680363874
transform 1 0 3568 0 -1 570
box -8 -3 46 105
use FILL  FILL_10100
timestamp 1680363874
transform 1 0 3608 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_637
timestamp 1680363874
transform 1 0 3616 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_559
timestamp 1680363874
transform -1 0 3728 0 -1 570
box -8 -3 104 105
use FILL  FILL_10101
timestamp 1680363874
transform 1 0 3728 0 -1 570
box -8 -3 16 105
use FILL  FILL_10102
timestamp 1680363874
transform 1 0 3736 0 -1 570
box -8 -3 16 105
use FILL  FILL_10103
timestamp 1680363874
transform 1 0 3744 0 -1 570
box -8 -3 16 105
use FILL  FILL_10104
timestamp 1680363874
transform 1 0 3752 0 -1 570
box -8 -3 16 105
use FILL  FILL_10106
timestamp 1680363874
transform 1 0 3760 0 -1 570
box -8 -3 16 105
use FILL  FILL_10108
timestamp 1680363874
transform 1 0 3768 0 -1 570
box -8 -3 16 105
use FILL  FILL_10110
timestamp 1680363874
transform 1 0 3776 0 -1 570
box -8 -3 16 105
use FILL  FILL_10111
timestamp 1680363874
transform 1 0 3784 0 -1 570
box -8 -3 16 105
use FILL  FILL_10112
timestamp 1680363874
transform 1 0 3792 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_638
timestamp 1680363874
transform -1 0 3816 0 -1 570
box -9 -3 26 105
use FILL  FILL_10113
timestamp 1680363874
transform 1 0 3816 0 -1 570
box -8 -3 16 105
use FILL  FILL_10115
timestamp 1680363874
transform 1 0 3824 0 -1 570
box -8 -3 16 105
use FILL  FILL_10117
timestamp 1680363874
transform 1 0 3832 0 -1 570
box -8 -3 16 105
use FILL  FILL_10119
timestamp 1680363874
transform 1 0 3840 0 -1 570
box -8 -3 16 105
use FILL  FILL_10134
timestamp 1680363874
transform 1 0 3848 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_367
timestamp 1680363874
transform -1 0 3896 0 -1 570
box -8 -3 46 105
use FILL  FILL_10135
timestamp 1680363874
transform 1 0 3896 0 -1 570
box -8 -3 16 105
use FILL  FILL_10136
timestamp 1680363874
transform 1 0 3904 0 -1 570
box -8 -3 16 105
use FILL  FILL_10137
timestamp 1680363874
transform 1 0 3912 0 -1 570
box -8 -3 16 105
use FILL  FILL_10138
timestamp 1680363874
transform 1 0 3920 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_368
timestamp 1680363874
transform -1 0 3968 0 -1 570
box -8 -3 46 105
use FILL  FILL_10139
timestamp 1680363874
transform 1 0 3968 0 -1 570
box -8 -3 16 105
use FILL  FILL_10140
timestamp 1680363874
transform 1 0 3976 0 -1 570
box -8 -3 16 105
use FILL  FILL_10141
timestamp 1680363874
transform 1 0 3984 0 -1 570
box -8 -3 16 105
use FILL  FILL_10142
timestamp 1680363874
transform 1 0 3992 0 -1 570
box -8 -3 16 105
use FILL  FILL_10143
timestamp 1680363874
transform 1 0 4000 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_113
timestamp 1680363874
transform -1 0 4032 0 -1 570
box -5 -3 28 105
use FILL  FILL_10144
timestamp 1680363874
transform 1 0 4032 0 -1 570
box -8 -3 16 105
use FILL  FILL_10145
timestamp 1680363874
transform 1 0 4040 0 -1 570
box -8 -3 16 105
use FILL  FILL_10146
timestamp 1680363874
transform 1 0 4048 0 -1 570
box -8 -3 16 105
use FILL  FILL_10147
timestamp 1680363874
transform 1 0 4056 0 -1 570
box -8 -3 16 105
use FILL  FILL_10148
timestamp 1680363874
transform 1 0 4064 0 -1 570
box -8 -3 16 105
use FILL  FILL_10149
timestamp 1680363874
transform 1 0 4072 0 -1 570
box -8 -3 16 105
use FILL  FILL_10150
timestamp 1680363874
transform 1 0 4080 0 -1 570
box -8 -3 16 105
use FILL  FILL_10151
timestamp 1680363874
transform 1 0 4088 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_641
timestamp 1680363874
transform 1 0 4096 0 -1 570
box -9 -3 26 105
use FILL  FILL_10152
timestamp 1680363874
transform 1 0 4112 0 -1 570
box -8 -3 16 105
use FILL  FILL_10153
timestamp 1680363874
transform 1 0 4120 0 -1 570
box -8 -3 16 105
use FILL  FILL_10154
timestamp 1680363874
transform 1 0 4128 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_400
timestamp 1680363874
transform 1 0 4136 0 -1 570
box -8 -3 46 105
use BUFX2  BUFX2_114
timestamp 1680363874
transform 1 0 4176 0 -1 570
box -5 -3 28 105
use FILL  FILL_10155
timestamp 1680363874
transform 1 0 4200 0 -1 570
box -8 -3 16 105
use FILL  FILL_10157
timestamp 1680363874
transform 1 0 4208 0 -1 570
box -8 -3 16 105
use FILL  FILL_10159
timestamp 1680363874
transform 1 0 4216 0 -1 570
box -8 -3 16 105
use FILL  FILL_10161
timestamp 1680363874
transform 1 0 4224 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_115
timestamp 1680363874
transform 1 0 4232 0 -1 570
box -5 -3 28 105
use FILL  FILL_10163
timestamp 1680363874
transform 1 0 4256 0 -1 570
box -8 -3 16 105
use FILL  FILL_10164
timestamp 1680363874
transform 1 0 4264 0 -1 570
box -8 -3 16 105
use FILL  FILL_10165
timestamp 1680363874
transform 1 0 4272 0 -1 570
box -8 -3 16 105
use FILL  FILL_10166
timestamp 1680363874
transform 1 0 4280 0 -1 570
box -8 -3 16 105
use FILL  FILL_10167
timestamp 1680363874
transform 1 0 4288 0 -1 570
box -8 -3 16 105
use FILL  FILL_10168
timestamp 1680363874
transform 1 0 4296 0 -1 570
box -8 -3 16 105
use FILL  FILL_10169
timestamp 1680363874
transform 1 0 4304 0 -1 570
box -8 -3 16 105
use FILL  FILL_10170
timestamp 1680363874
transform 1 0 4312 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_643
timestamp 1680363874
transform 1 0 4320 0 -1 570
box -9 -3 26 105
use FILL  FILL_10171
timestamp 1680363874
transform 1 0 4336 0 -1 570
box -8 -3 16 105
use FILL  FILL_10172
timestamp 1680363874
transform 1 0 4344 0 -1 570
box -8 -3 16 105
use FILL  FILL_10174
timestamp 1680363874
transform 1 0 4352 0 -1 570
box -8 -3 16 105
use FILL  FILL_10178
timestamp 1680363874
transform 1 0 4360 0 -1 570
box -8 -3 16 105
use FILL  FILL_10179
timestamp 1680363874
transform 1 0 4368 0 -1 570
box -8 -3 16 105
use FILL  FILL_10180
timestamp 1680363874
transform 1 0 4376 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_401
timestamp 1680363874
transform 1 0 4384 0 -1 570
box -8 -3 46 105
use FILL  FILL_10181
timestamp 1680363874
transform 1 0 4424 0 -1 570
box -8 -3 16 105
use FILL  FILL_10182
timestamp 1680363874
transform 1 0 4432 0 -1 570
box -8 -3 16 105
use FILL  FILL_10183
timestamp 1680363874
transform 1 0 4440 0 -1 570
box -8 -3 16 105
use FILL  FILL_10184
timestamp 1680363874
transform 1 0 4448 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_644
timestamp 1680363874
transform 1 0 4456 0 -1 570
box -9 -3 26 105
use FILL  FILL_10185
timestamp 1680363874
transform 1 0 4472 0 -1 570
box -8 -3 16 105
use FILL  FILL_10186
timestamp 1680363874
transform 1 0 4480 0 -1 570
box -8 -3 16 105
use FILL  FILL_10187
timestamp 1680363874
transform 1 0 4488 0 -1 570
box -8 -3 16 105
use FILL  FILL_10188
timestamp 1680363874
transform 1 0 4496 0 -1 570
box -8 -3 16 105
use FILL  FILL_10189
timestamp 1680363874
transform 1 0 4504 0 -1 570
box -8 -3 16 105
use FILL  FILL_10190
timestamp 1680363874
transform 1 0 4512 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_563
timestamp 1680363874
transform 1 0 4520 0 -1 570
box -8 -3 104 105
use FILL  FILL_10198
timestamp 1680363874
transform 1 0 4616 0 -1 570
box -8 -3 16 105
use FILL  FILL_10199
timestamp 1680363874
transform 1 0 4624 0 -1 570
box -8 -3 16 105
use FILL  FILL_10201
timestamp 1680363874
transform 1 0 4632 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_372
timestamp 1680363874
transform 1 0 4640 0 -1 570
box -8 -3 46 105
use FILL  FILL_10203
timestamp 1680363874
transform 1 0 4680 0 -1 570
box -8 -3 16 105
use FILL  FILL_10204
timestamp 1680363874
transform 1 0 4688 0 -1 570
box -8 -3 16 105
use FILL  FILL_10205
timestamp 1680363874
transform 1 0 4696 0 -1 570
box -8 -3 16 105
use FILL  FILL_10206
timestamp 1680363874
transform 1 0 4704 0 -1 570
box -8 -3 16 105
use FILL  FILL_10207
timestamp 1680363874
transform 1 0 4712 0 -1 570
box -8 -3 16 105
use FILL  FILL_10208
timestamp 1680363874
transform 1 0 4720 0 -1 570
box -8 -3 16 105
use FILL  FILL_10209
timestamp 1680363874
transform 1 0 4728 0 -1 570
box -8 -3 16 105
use FILL  FILL_10210
timestamp 1680363874
transform 1 0 4736 0 -1 570
box -8 -3 16 105
use FILL  FILL_10211
timestamp 1680363874
transform 1 0 4744 0 -1 570
box -8 -3 16 105
use FILL  FILL_10212
timestamp 1680363874
transform 1 0 4752 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_647
timestamp 1680363874
transform 1 0 4760 0 -1 570
box -9 -3 26 105
use FILL  FILL_10213
timestamp 1680363874
transform 1 0 4776 0 -1 570
box -8 -3 16 105
use FILL  FILL_10214
timestamp 1680363874
transform 1 0 4784 0 -1 570
box -8 -3 16 105
use FILL  FILL_10215
timestamp 1680363874
transform 1 0 4792 0 -1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_85
timestamp 1680363874
transform 1 0 4851 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_9156
timestamp 1680363874
transform 1 0 84 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9278
timestamp 1680363874
transform 1 0 100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9279
timestamp 1680363874
transform 1 0 124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9148
timestamp 1680363874
transform 1 0 140 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9157
timestamp 1680363874
transform 1 0 132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9280
timestamp 1680363874
transform 1 0 140 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8357
timestamp 1680363874
transform 1 0 140 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9281
timestamp 1680363874
transform 1 0 164 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8253
timestamp 1680363874
transform 1 0 188 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9282
timestamp 1680363874
transform 1 0 180 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8358
timestamp 1680363874
transform 1 0 180 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9158
timestamp 1680363874
transform 1 0 188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9159
timestamp 1680363874
transform 1 0 204 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8254
timestamp 1680363874
transform 1 0 252 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9149
timestamp 1680363874
transform 1 0 252 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9160
timestamp 1680363874
transform 1 0 236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9283
timestamp 1680363874
transform 1 0 252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9161
timestamp 1680363874
transform 1 0 284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9284
timestamp 1680363874
transform 1 0 276 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8241
timestamp 1680363874
transform 1 0 324 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9162
timestamp 1680363874
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9285
timestamp 1680363874
transform 1 0 356 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8242
timestamp 1680363874
transform 1 0 388 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9163
timestamp 1680363874
transform 1 0 388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9164
timestamp 1680363874
transform 1 0 404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9165
timestamp 1680363874
transform 1 0 412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9286
timestamp 1680363874
transform 1 0 380 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8342
timestamp 1680363874
transform 1 0 388 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9287
timestamp 1680363874
transform 1 0 396 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8343
timestamp 1680363874
transform 1 0 412 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9288
timestamp 1680363874
transform 1 0 420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8282
timestamp 1680363874
transform 1 0 532 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9166
timestamp 1680363874
transform 1 0 476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9167
timestamp 1680363874
transform 1 0 532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9289
timestamp 1680363874
transform 1 0 556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9290
timestamp 1680363874
transform 1 0 572 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8283
timestamp 1680363874
transform 1 0 620 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9168
timestamp 1680363874
transform 1 0 628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9291
timestamp 1680363874
transform 1 0 628 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8255
timestamp 1680363874
transform 1 0 668 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8284
timestamp 1680363874
transform 1 0 652 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9169
timestamp 1680363874
transform 1 0 636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9170
timestamp 1680363874
transform 1 0 652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9171
timestamp 1680363874
transform 1 0 668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9292
timestamp 1680363874
transform 1 0 644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9293
timestamp 1680363874
transform 1 0 660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9294
timestamp 1680363874
transform 1 0 676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9172
timestamp 1680363874
transform 1 0 692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9173
timestamp 1680363874
transform 1 0 700 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8344
timestamp 1680363874
transform 1 0 692 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9295
timestamp 1680363874
transform 1 0 708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9296
timestamp 1680363874
transform 1 0 724 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8345
timestamp 1680363874
transform 1 0 732 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8243
timestamp 1680363874
transform 1 0 780 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8313
timestamp 1680363874
transform 1 0 772 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8359
timestamp 1680363874
transform 1 0 772 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8285
timestamp 1680363874
transform 1 0 796 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9146
timestamp 1680363874
transform 1 0 836 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_9150
timestamp 1680363874
transform 1 0 828 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9174
timestamp 1680363874
transform 1 0 780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9175
timestamp 1680363874
transform 1 0 804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9176
timestamp 1680363874
transform 1 0 820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9297
timestamp 1680363874
transform 1 0 788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9298
timestamp 1680363874
transform 1 0 796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9299
timestamp 1680363874
transform 1 0 812 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8393
timestamp 1680363874
transform 1 0 804 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8360
timestamp 1680363874
transform 1 0 828 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9177
timestamp 1680363874
transform 1 0 844 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8346
timestamp 1680363874
transform 1 0 844 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8256
timestamp 1680363874
transform 1 0 868 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9178
timestamp 1680363874
transform 1 0 868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9151
timestamp 1680363874
transform 1 0 900 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9179
timestamp 1680363874
transform 1 0 916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9180
timestamp 1680363874
transform 1 0 932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9300
timestamp 1680363874
transform 1 0 908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9301
timestamp 1680363874
transform 1 0 924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9302
timestamp 1680363874
transform 1 0 940 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8361
timestamp 1680363874
transform 1 0 908 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8394
timestamp 1680363874
transform 1 0 948 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9147
timestamp 1680363874
transform 1 0 972 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_9152
timestamp 1680363874
transform 1 0 964 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8244
timestamp 1680363874
transform 1 0 1012 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8257
timestamp 1680363874
transform 1 0 1004 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9153
timestamp 1680363874
transform 1 0 1004 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9181
timestamp 1680363874
transform 1 0 988 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8314
timestamp 1680363874
transform 1 0 1004 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9182
timestamp 1680363874
transform 1 0 1012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9183
timestamp 1680363874
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9184
timestamp 1680363874
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9303
timestamp 1680363874
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9304
timestamp 1680363874
transform 1 0 1028 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8362
timestamp 1680363874
transform 1 0 1012 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9185
timestamp 1680363874
transform 1 0 1052 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8258
timestamp 1680363874
transform 1 0 1068 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9305
timestamp 1680363874
transform 1 0 1076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9306
timestamp 1680363874
transform 1 0 1084 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8315
timestamp 1680363874
transform 1 0 1092 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9186
timestamp 1680363874
transform 1 0 1116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9187
timestamp 1680363874
transform 1 0 1164 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8286
timestamp 1680363874
transform 1 0 1212 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8316
timestamp 1680363874
transform 1 0 1188 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9188
timestamp 1680363874
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9189
timestamp 1680363874
transform 1 0 1212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9307
timestamp 1680363874
transform 1 0 1188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9308
timestamp 1680363874
transform 1 0 1228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8245
timestamp 1680363874
transform 1 0 1276 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8287
timestamp 1680363874
transform 1 0 1284 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8317
timestamp 1680363874
transform 1 0 1284 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9190
timestamp 1680363874
transform 1 0 1308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9309
timestamp 1680363874
transform 1 0 1260 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8363
timestamp 1680363874
transform 1 0 1308 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9310
timestamp 1680363874
transform 1 0 1348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9191
timestamp 1680363874
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9192
timestamp 1680363874
transform 1 0 1372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9193
timestamp 1680363874
transform 1 0 1388 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8259
timestamp 1680363874
transform 1 0 1404 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8288
timestamp 1680363874
transform 1 0 1404 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9194
timestamp 1680363874
transform 1 0 1404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9311
timestamp 1680363874
transform 1 0 1380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9312
timestamp 1680363874
transform 1 0 1396 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8364
timestamp 1680363874
transform 1 0 1380 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8395
timestamp 1680363874
transform 1 0 1404 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8318
timestamp 1680363874
transform 1 0 1420 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9195
timestamp 1680363874
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9313
timestamp 1680363874
transform 1 0 1412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9314
timestamp 1680363874
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9196
timestamp 1680363874
transform 1 0 1532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9315
timestamp 1680363874
transform 1 0 1524 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8235
timestamp 1680363874
transform 1 0 1548 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8236
timestamp 1680363874
transform 1 0 1588 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8246
timestamp 1680363874
transform 1 0 1564 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8260
timestamp 1680363874
transform 1 0 1596 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8289
timestamp 1680363874
transform 1 0 1572 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9197
timestamp 1680363874
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9198
timestamp 1680363874
transform 1 0 1580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9199
timestamp 1680363874
transform 1 0 1596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9316
timestamp 1680363874
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8365
timestamp 1680363874
transform 1 0 1572 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9317
timestamp 1680363874
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8247
timestamp 1680363874
transform 1 0 1620 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8261
timestamp 1680363874
transform 1 0 1612 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8262
timestamp 1680363874
transform 1 0 1652 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8290
timestamp 1680363874
transform 1 0 1636 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8291
timestamp 1680363874
transform 1 0 1652 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9200
timestamp 1680363874
transform 1 0 1636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9201
timestamp 1680363874
transform 1 0 1652 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8319
timestamp 1680363874
transform 1 0 1660 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9318
timestamp 1680363874
transform 1 0 1628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9319
timestamp 1680363874
transform 1 0 1644 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8366
timestamp 1680363874
transform 1 0 1628 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8396
timestamp 1680363874
transform 1 0 1628 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9320
timestamp 1680363874
transform 1 0 1676 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8237
timestamp 1680363874
transform 1 0 1700 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9321
timestamp 1680363874
transform 1 0 1700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9322
timestamp 1680363874
transform 1 0 1708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8367
timestamp 1680363874
transform 1 0 1708 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8397
timestamp 1680363874
transform 1 0 1708 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8292
timestamp 1680363874
transform 1 0 1740 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9202
timestamp 1680363874
transform 1 0 1724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9203
timestamp 1680363874
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9323
timestamp 1680363874
transform 1 0 1732 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9324
timestamp 1680363874
transform 1 0 1748 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8368
timestamp 1680363874
transform 1 0 1724 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9325
timestamp 1680363874
transform 1 0 1772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9326
timestamp 1680363874
transform 1 0 1780 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8369
timestamp 1680363874
transform 1 0 1788 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8398
timestamp 1680363874
transform 1 0 1780 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8293
timestamp 1680363874
transform 1 0 1844 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9204
timestamp 1680363874
transform 1 0 1828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9205
timestamp 1680363874
transform 1 0 1844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9327
timestamp 1680363874
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9328
timestamp 1680363874
transform 1 0 1852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9206
timestamp 1680363874
transform 1 0 1876 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8399
timestamp 1680363874
transform 1 0 1868 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8248
timestamp 1680363874
transform 1 0 1908 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8320
timestamp 1680363874
transform 1 0 1900 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9329
timestamp 1680363874
transform 1 0 1900 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8263
timestamp 1680363874
transform 1 0 1964 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8294
timestamp 1680363874
transform 1 0 1948 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8295
timestamp 1680363874
transform 1 0 1972 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8321
timestamp 1680363874
transform 1 0 1924 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9207
timestamp 1680363874
transform 1 0 1972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9330
timestamp 1680363874
transform 1 0 1924 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8370
timestamp 1680363874
transform 1 0 1924 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8371
timestamp 1680363874
transform 1 0 1988 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8372
timestamp 1680363874
transform 1 0 2004 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8249
timestamp 1680363874
transform 1 0 2028 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8264
timestamp 1680363874
transform 1 0 2028 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8250
timestamp 1680363874
transform 1 0 2060 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8296
timestamp 1680363874
transform 1 0 2044 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9208
timestamp 1680363874
transform 1 0 2020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9209
timestamp 1680363874
transform 1 0 2028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9210
timestamp 1680363874
transform 1 0 2044 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8322
timestamp 1680363874
transform 1 0 2052 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9211
timestamp 1680363874
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9331
timestamp 1680363874
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9332
timestamp 1680363874
transform 1 0 2052 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8373
timestamp 1680363874
transform 1 0 2052 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8400
timestamp 1680363874
transform 1 0 2052 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8251
timestamp 1680363874
transform 1 0 2100 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8265
timestamp 1680363874
transform 1 0 2100 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9333
timestamp 1680363874
transform 1 0 2100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9334
timestamp 1680363874
transform 1 0 2108 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8401
timestamp 1680363874
transform 1 0 2100 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8266
timestamp 1680363874
transform 1 0 2132 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8297
timestamp 1680363874
transform 1 0 2148 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9212
timestamp 1680363874
transform 1 0 2132 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8323
timestamp 1680363874
transform 1 0 2140 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9213
timestamp 1680363874
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9335
timestamp 1680363874
transform 1 0 2140 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8238
timestamp 1680363874
transform 1 0 2180 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8267
timestamp 1680363874
transform 1 0 2172 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9214
timestamp 1680363874
transform 1 0 2172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9215
timestamp 1680363874
transform 1 0 2204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9336
timestamp 1680363874
transform 1 0 2172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9337
timestamp 1680363874
transform 1 0 2180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9338
timestamp 1680363874
transform 1 0 2196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9339
timestamp 1680363874
transform 1 0 2212 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8374
timestamp 1680363874
transform 1 0 2196 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8402
timestamp 1680363874
transform 1 0 2204 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8268
timestamp 1680363874
transform 1 0 2228 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8403
timestamp 1680363874
transform 1 0 2236 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8269
timestamp 1680363874
transform 1 0 2260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8298
timestamp 1680363874
transform 1 0 2332 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8299
timestamp 1680363874
transform 1 0 2348 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9216
timestamp 1680363874
transform 1 0 2252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9217
timestamp 1680363874
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8324
timestamp 1680363874
transform 1 0 2332 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8239
timestamp 1680363874
transform 1 0 2380 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8240
timestamp 1680363874
transform 1 0 2404 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9218
timestamp 1680363874
transform 1 0 2348 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9219
timestamp 1680363874
transform 1 0 2364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9220
timestamp 1680363874
transform 1 0 2404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9340
timestamp 1680363874
transform 1 0 2332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8375
timestamp 1680363874
transform 1 0 2284 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9341
timestamp 1680363874
transform 1 0 2356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9342
timestamp 1680363874
transform 1 0 2444 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8376
timestamp 1680363874
transform 1 0 2444 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8270
timestamp 1680363874
transform 1 0 2532 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9221
timestamp 1680363874
transform 1 0 2492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9222
timestamp 1680363874
transform 1 0 2548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9343
timestamp 1680363874
transform 1 0 2468 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8377
timestamp 1680363874
transform 1 0 2468 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8378
timestamp 1680363874
transform 1 0 2532 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8325
timestamp 1680363874
transform 1 0 2572 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9223
timestamp 1680363874
transform 1 0 2636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9344
timestamp 1680363874
transform 1 0 2588 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8347
timestamp 1680363874
transform 1 0 2612 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8379
timestamp 1680363874
transform 1 0 2588 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8380
timestamp 1680363874
transform 1 0 2676 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9224
timestamp 1680363874
transform 1 0 2700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9345
timestamp 1680363874
transform 1 0 2708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9225
timestamp 1680363874
transform 1 0 2740 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8348
timestamp 1680363874
transform 1 0 2740 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8271
timestamp 1680363874
transform 1 0 2764 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9154
timestamp 1680363874
transform 1 0 2764 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8326
timestamp 1680363874
transform 1 0 2764 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8272
timestamp 1680363874
transform 1 0 2796 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9155
timestamp 1680363874
transform 1 0 2796 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9226
timestamp 1680363874
transform 1 0 2780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9346
timestamp 1680363874
transform 1 0 2764 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9347
timestamp 1680363874
transform 1 0 2772 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8349
timestamp 1680363874
transform 1 0 2780 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8327
timestamp 1680363874
transform 1 0 2836 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9227
timestamp 1680363874
transform 1 0 2844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9348
timestamp 1680363874
transform 1 0 2828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9228
timestamp 1680363874
transform 1 0 2860 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8273
timestamp 1680363874
transform 1 0 2924 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8300
timestamp 1680363874
transform 1 0 2940 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8301
timestamp 1680363874
transform 1 0 2980 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9229
timestamp 1680363874
transform 1 0 2892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9230
timestamp 1680363874
transform 1 0 2908 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8328
timestamp 1680363874
transform 1 0 2916 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9231
timestamp 1680363874
transform 1 0 2924 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8329
timestamp 1680363874
transform 1 0 2932 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9232
timestamp 1680363874
transform 1 0 2940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9233
timestamp 1680363874
transform 1 0 2948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9234
timestamp 1680363874
transform 1 0 2980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9349
timestamp 1680363874
transform 1 0 2900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9350
timestamp 1680363874
transform 1 0 2916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9351
timestamp 1680363874
transform 1 0 2924 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8381
timestamp 1680363874
transform 1 0 2900 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9352
timestamp 1680363874
transform 1 0 3028 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8382
timestamp 1680363874
transform 1 0 2948 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8274
timestamp 1680363874
transform 1 0 3132 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8302
timestamp 1680363874
transform 1 0 3100 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8303
timestamp 1680363874
transform 1 0 3140 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8330
timestamp 1680363874
transform 1 0 3052 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9235
timestamp 1680363874
transform 1 0 3100 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8331
timestamp 1680363874
transform 1 0 3116 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9236
timestamp 1680363874
transform 1 0 3132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9237
timestamp 1680363874
transform 1 0 3140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9353
timestamp 1680363874
transform 1 0 3052 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8383
timestamp 1680363874
transform 1 0 3052 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8384
timestamp 1680363874
transform 1 0 3084 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8275
timestamp 1680363874
transform 1 0 3164 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9238
timestamp 1680363874
transform 1 0 3148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9239
timestamp 1680363874
transform 1 0 3156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9240
timestamp 1680363874
transform 1 0 3172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9241
timestamp 1680363874
transform 1 0 3188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9354
timestamp 1680363874
transform 1 0 3156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9355
timestamp 1680363874
transform 1 0 3164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9356
timestamp 1680363874
transform 1 0 3180 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8350
timestamp 1680363874
transform 1 0 3196 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9357
timestamp 1680363874
transform 1 0 3220 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8304
timestamp 1680363874
transform 1 0 3276 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9242
timestamp 1680363874
transform 1 0 3284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9358
timestamp 1680363874
transform 1 0 3268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9359
timestamp 1680363874
transform 1 0 3276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9360
timestamp 1680363874
transform 1 0 3292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9361
timestamp 1680363874
transform 1 0 3300 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8305
timestamp 1680363874
transform 1 0 3324 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9243
timestamp 1680363874
transform 1 0 3324 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8252
timestamp 1680363874
transform 1 0 3340 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9244
timestamp 1680363874
transform 1 0 3364 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8351
timestamp 1680363874
transform 1 0 3364 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8404
timestamp 1680363874
transform 1 0 3364 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8276
timestamp 1680363874
transform 1 0 3404 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8306
timestamp 1680363874
transform 1 0 3412 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9245
timestamp 1680363874
transform 1 0 3396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9246
timestamp 1680363874
transform 1 0 3412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9362
timestamp 1680363874
transform 1 0 3388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9363
timestamp 1680363874
transform 1 0 3404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9364
timestamp 1680363874
transform 1 0 3412 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8277
timestamp 1680363874
transform 1 0 3452 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8307
timestamp 1680363874
transform 1 0 3444 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8308
timestamp 1680363874
transform 1 0 3484 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9247
timestamp 1680363874
transform 1 0 3444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9248
timestamp 1680363874
transform 1 0 3452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9249
timestamp 1680363874
transform 1 0 3484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9365
timestamp 1680363874
transform 1 0 3532 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8278
timestamp 1680363874
transform 1 0 3580 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8279
timestamp 1680363874
transform 1 0 3596 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8309
timestamp 1680363874
transform 1 0 3572 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8310
timestamp 1680363874
transform 1 0 3612 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8332
timestamp 1680363874
transform 1 0 3564 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9250
timestamp 1680363874
transform 1 0 3572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9251
timestamp 1680363874
transform 1 0 3580 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8333
timestamp 1680363874
transform 1 0 3588 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9252
timestamp 1680363874
transform 1 0 3612 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8334
timestamp 1680363874
transform 1 0 3660 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9366
timestamp 1680363874
transform 1 0 3564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9253
timestamp 1680363874
transform 1 0 3684 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8335
timestamp 1680363874
transform 1 0 3716 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9254
timestamp 1680363874
transform 1 0 3724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9367
timestamp 1680363874
transform 1 0 3660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9368
timestamp 1680363874
transform 1 0 3676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9369
timestamp 1680363874
transform 1 0 3692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9370
timestamp 1680363874
transform 1 0 3708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8385
timestamp 1680363874
transform 1 0 3684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8352
timestamp 1680363874
transform 1 0 3724 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8336
timestamp 1680363874
transform 1 0 3740 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9255
timestamp 1680363874
transform 1 0 3788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9256
timestamp 1680363874
transform 1 0 3820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9371
timestamp 1680363874
transform 1 0 3740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8353
timestamp 1680363874
transform 1 0 3764 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8386
timestamp 1680363874
transform 1 0 3780 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8337
timestamp 1680363874
transform 1 0 3828 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8311
timestamp 1680363874
transform 1 0 3900 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8338
timestamp 1680363874
transform 1 0 3852 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8312
timestamp 1680363874
transform 1 0 3940 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9257
timestamp 1680363874
transform 1 0 3900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9258
timestamp 1680363874
transform 1 0 3932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9259
timestamp 1680363874
transform 1 0 3940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9372
timestamp 1680363874
transform 1 0 3852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9373
timestamp 1680363874
transform 1 0 3948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9374
timestamp 1680363874
transform 1 0 3972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9260
timestamp 1680363874
transform 1 0 3988 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9261
timestamp 1680363874
transform 1 0 4020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9262
timestamp 1680363874
transform 1 0 4036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9263
timestamp 1680363874
transform 1 0 4092 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8339
timestamp 1680363874
transform 1 0 4116 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9375
timestamp 1680363874
transform 1 0 4012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9376
timestamp 1680363874
transform 1 0 4028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9377
timestamp 1680363874
transform 1 0 4116 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8405
timestamp 1680363874
transform 1 0 4052 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9264
timestamp 1680363874
transform 1 0 4132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9378
timestamp 1680363874
transform 1 0 4188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9265
timestamp 1680363874
transform 1 0 4196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9379
timestamp 1680363874
transform 1 0 4196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9266
timestamp 1680363874
transform 1 0 4236 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8354
timestamp 1680363874
transform 1 0 4220 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9380
timestamp 1680363874
transform 1 0 4228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8406
timestamp 1680363874
transform 1 0 4236 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9267
timestamp 1680363874
transform 1 0 4252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9268
timestamp 1680363874
transform 1 0 4268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9269
timestamp 1680363874
transform 1 0 4292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9381
timestamp 1680363874
transform 1 0 4276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9382
timestamp 1680363874
transform 1 0 4284 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8355
timestamp 1680363874
transform 1 0 4292 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9383
timestamp 1680363874
transform 1 0 4300 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8387
timestamp 1680363874
transform 1 0 4276 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8388
timestamp 1680363874
transform 1 0 4300 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9270
timestamp 1680363874
transform 1 0 4316 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8356
timestamp 1680363874
transform 1 0 4316 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8389
timestamp 1680363874
transform 1 0 4316 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8407
timestamp 1680363874
transform 1 0 4308 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8390
timestamp 1680363874
transform 1 0 4356 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8280
timestamp 1680363874
transform 1 0 4404 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9271
timestamp 1680363874
transform 1 0 4396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9384
timestamp 1680363874
transform 1 0 4444 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8391
timestamp 1680363874
transform 1 0 4428 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9272
timestamp 1680363874
transform 1 0 4468 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8392
timestamp 1680363874
transform 1 0 4460 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9273
timestamp 1680363874
transform 1 0 4508 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8340
timestamp 1680363874
transform 1 0 4532 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8341
timestamp 1680363874
transform 1 0 4556 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9385
timestamp 1680363874
transform 1 0 4556 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8408
timestamp 1680363874
transform 1 0 4508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8281
timestamp 1680363874
transform 1 0 4572 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9274
timestamp 1680363874
transform 1 0 4572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9386
timestamp 1680363874
transform 1 0 4588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9275
timestamp 1680363874
transform 1 0 4620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9387
timestamp 1680363874
transform 1 0 4612 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8409
timestamp 1680363874
transform 1 0 4596 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9388
timestamp 1680363874
transform 1 0 4644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9276
timestamp 1680363874
transform 1 0 4668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9277
timestamp 1680363874
transform 1 0 4748 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9389
timestamp 1680363874
transform 1 0 4780 0 1 405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_86
timestamp 1680363874
transform 1 0 48 0 1 370
box -10 -3 10 3
use FILL  FILL_10216
timestamp 1680363874
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_10217
timestamp 1680363874
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_10218
timestamp 1680363874
transform 1 0 88 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_175
timestamp 1680363874
transform 1 0 96 0 1 370
box -8 -3 34 105
use FILL  FILL_10219
timestamp 1680363874
transform 1 0 128 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_63
timestamp 1680363874
transform 1 0 136 0 1 370
box -8 -3 32 105
use INVX2  INVX2_648
timestamp 1680363874
transform 1 0 160 0 1 370
box -9 -3 26 105
use FILL  FILL_10220
timestamp 1680363874
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_10223
timestamp 1680363874
transform 1 0 184 0 1 370
box -8 -3 16 105
use INVX2  INVX2_649
timestamp 1680363874
transform 1 0 192 0 1 370
box -9 -3 26 105
use FILL  FILL_10225
timestamp 1680363874
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_10229
timestamp 1680363874
transform 1 0 216 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_176
timestamp 1680363874
transform 1 0 224 0 1 370
box -8 -3 34 105
use NAND2X1  NAND2X1_64
timestamp 1680363874
transform -1 0 280 0 1 370
box -8 -3 32 105
use FILL  FILL_10231
timestamp 1680363874
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_10235
timestamp 1680363874
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_10237
timestamp 1680363874
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_10239
timestamp 1680363874
transform 1 0 304 0 1 370
box -8 -3 16 105
use FILL  FILL_10241
timestamp 1680363874
transform 1 0 312 0 1 370
box -8 -3 16 105
use FILL  FILL_10243
timestamp 1680363874
transform 1 0 320 0 1 370
box -8 -3 16 105
use FILL  FILL_10245
timestamp 1680363874
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_10247
timestamp 1680363874
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_10249
timestamp 1680363874
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_10250
timestamp 1680363874
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_10251
timestamp 1680363874
transform 1 0 360 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_373
timestamp 1680363874
transform 1 0 368 0 1 370
box -8 -3 46 105
use INVX2  INVX2_650
timestamp 1680363874
transform -1 0 424 0 1 370
box -9 -3 26 105
use FILL  FILL_10252
timestamp 1680363874
transform 1 0 424 0 1 370
box -8 -3 16 105
use FILL  FILL_10253
timestamp 1680363874
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_10254
timestamp 1680363874
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_10255
timestamp 1680363874
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_10256
timestamp 1680363874
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_10257
timestamp 1680363874
transform 1 0 464 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_566
timestamp 1680363874
transform -1 0 568 0 1 370
box -8 -3 104 105
use FILL  FILL_10258
timestamp 1680363874
transform 1 0 568 0 1 370
box -8 -3 16 105
use FILL  FILL_10259
timestamp 1680363874
transform 1 0 576 0 1 370
box -8 -3 16 105
use INVX2  INVX2_651
timestamp 1680363874
transform 1 0 584 0 1 370
box -9 -3 26 105
use FILL  FILL_10260
timestamp 1680363874
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_10261
timestamp 1680363874
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_10262
timestamp 1680363874
transform 1 0 616 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8410
timestamp 1680363874
transform 1 0 644 0 1 375
box -3 -3 3 3
use INVX2  INVX2_652
timestamp 1680363874
transform 1 0 624 0 1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_403
timestamp 1680363874
transform -1 0 680 0 1 370
box -8 -3 46 105
use FILL  FILL_10263
timestamp 1680363874
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_10271
timestamp 1680363874
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_10272
timestamp 1680363874
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_10273
timestamp 1680363874
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_10274
timestamp 1680363874
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_10275
timestamp 1680363874
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_10276
timestamp 1680363874
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_10278
timestamp 1680363874
transform 1 0 736 0 1 370
box -8 -3 16 105
use FILL  FILL_10280
timestamp 1680363874
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_10282
timestamp 1680363874
transform 1 0 752 0 1 370
box -8 -3 16 105
use FILL  FILL_10283
timestamp 1680363874
transform 1 0 760 0 1 370
box -8 -3 16 105
use INVX2  INVX2_654
timestamp 1680363874
transform 1 0 768 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_374
timestamp 1680363874
transform -1 0 824 0 1 370
box -8 -3 46 105
use FILL  FILL_10284
timestamp 1680363874
transform 1 0 824 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_75
timestamp 1680363874
transform 1 0 832 0 1 370
box -8 -3 40 105
use FILL  FILL_10290
timestamp 1680363874
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_10292
timestamp 1680363874
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_10294
timestamp 1680363874
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_10296
timestamp 1680363874
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_10298
timestamp 1680363874
transform 1 0 896 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8411
timestamp 1680363874
transform 1 0 940 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_407
timestamp 1680363874
transform 1 0 904 0 1 370
box -8 -3 46 105
use FILL  FILL_10300
timestamp 1680363874
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_10301
timestamp 1680363874
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_10302
timestamp 1680363874
transform 1 0 960 0 1 370
box -8 -3 16 105
use FILL  FILL_10303
timestamp 1680363874
transform 1 0 968 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_77
timestamp 1680363874
transform 1 0 976 0 1 370
box -8 -3 40 105
use OAI22X1  OAI22X1_408
timestamp 1680363874
transform 1 0 1008 0 1 370
box -8 -3 46 105
use FILL  FILL_10304
timestamp 1680363874
transform 1 0 1048 0 1 370
box -8 -3 16 105
use FILL  FILL_10305
timestamp 1680363874
transform 1 0 1056 0 1 370
box -8 -3 16 105
use FILL  FILL_10306
timestamp 1680363874
transform 1 0 1064 0 1 370
box -8 -3 16 105
use FILL  FILL_10307
timestamp 1680363874
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_10308
timestamp 1680363874
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_10309
timestamp 1680363874
transform 1 0 1088 0 1 370
box -8 -3 16 105
use INVX2  INVX2_655
timestamp 1680363874
transform 1 0 1096 0 1 370
box -9 -3 26 105
use FILL  FILL_10310
timestamp 1680363874
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_10311
timestamp 1680363874
transform 1 0 1120 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8412
timestamp 1680363874
transform 1 0 1140 0 1 375
box -3 -3 3 3
use FILL  FILL_10312
timestamp 1680363874
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_10313
timestamp 1680363874
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_10314
timestamp 1680363874
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_10315
timestamp 1680363874
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_10316
timestamp 1680363874
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_10317
timestamp 1680363874
transform 1 0 1168 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8413
timestamp 1680363874
transform 1 0 1196 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_376
timestamp 1680363874
transform 1 0 1176 0 1 370
box -8 -3 46 105
use FILL  FILL_10318
timestamp 1680363874
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_10326
timestamp 1680363874
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_10327
timestamp 1680363874
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_10328
timestamp 1680363874
transform 1 0 1240 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8414
timestamp 1680363874
transform 1 0 1292 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8415
timestamp 1680363874
transform 1 0 1340 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_570
timestamp 1680363874
transform 1 0 1248 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_8416
timestamp 1680363874
transform 1 0 1356 0 1 375
box -3 -3 3 3
use FILL  FILL_10329
timestamp 1680363874
transform 1 0 1344 0 1 370
box -8 -3 16 105
use FILL  FILL_10339
timestamp 1680363874
transform 1 0 1352 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_411
timestamp 1680363874
transform -1 0 1400 0 1 370
box -8 -3 46 105
use FILL  FILL_10340
timestamp 1680363874
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_10341
timestamp 1680363874
transform 1 0 1408 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8417
timestamp 1680363874
transform 1 0 1444 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_379
timestamp 1680363874
transform -1 0 1456 0 1 370
box -8 -3 46 105
use FILL  FILL_10342
timestamp 1680363874
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_10343
timestamp 1680363874
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_10344
timestamp 1680363874
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_10345
timestamp 1680363874
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_10346
timestamp 1680363874
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_10347
timestamp 1680363874
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_10348
timestamp 1680363874
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_10349
timestamp 1680363874
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_10350
timestamp 1680363874
transform 1 0 1520 0 1 370
box -8 -3 16 105
use INVX2  INVX2_661
timestamp 1680363874
transform 1 0 1528 0 1 370
box -9 -3 26 105
use FILL  FILL_10354
timestamp 1680363874
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_10355
timestamp 1680363874
transform 1 0 1552 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_380
timestamp 1680363874
transform 1 0 1560 0 1 370
box -8 -3 46 105
use FILL  FILL_10356
timestamp 1680363874
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_10357
timestamp 1680363874
transform 1 0 1608 0 1 370
box -8 -3 16 105
use FILL  FILL_10358
timestamp 1680363874
transform 1 0 1616 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_413
timestamp 1680363874
transform -1 0 1664 0 1 370
box -8 -3 46 105
use FILL  FILL_10359
timestamp 1680363874
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_10360
timestamp 1680363874
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_10361
timestamp 1680363874
transform 1 0 1680 0 1 370
box -8 -3 16 105
use FILL  FILL_10362
timestamp 1680363874
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_10363
timestamp 1680363874
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_10364
timestamp 1680363874
transform 1 0 1704 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_414
timestamp 1680363874
transform -1 0 1752 0 1 370
box -8 -3 46 105
use FILL  FILL_10365
timestamp 1680363874
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_10366
timestamp 1680363874
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_10367
timestamp 1680363874
transform 1 0 1768 0 1 370
box -8 -3 16 105
use FILL  FILL_10368
timestamp 1680363874
transform 1 0 1776 0 1 370
box -8 -3 16 105
use FILL  FILL_10369
timestamp 1680363874
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_10370
timestamp 1680363874
transform 1 0 1792 0 1 370
box -8 -3 16 105
use FILL  FILL_10374
timestamp 1680363874
transform 1 0 1800 0 1 370
box -8 -3 16 105
use FILL  FILL_10376
timestamp 1680363874
transform 1 0 1808 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_416
timestamp 1680363874
transform -1 0 1856 0 1 370
box -8 -3 46 105
use FILL  FILL_10378
timestamp 1680363874
transform 1 0 1856 0 1 370
box -8 -3 16 105
use FILL  FILL_10380
timestamp 1680363874
transform 1 0 1864 0 1 370
box -8 -3 16 105
use BUFX2  BUFX2_116
timestamp 1680363874
transform 1 0 1872 0 1 370
box -5 -3 28 105
use FILL  FILL_10382
timestamp 1680363874
transform 1 0 1896 0 1 370
box -8 -3 16 105
use FILL  FILL_10383
timestamp 1680363874
transform 1 0 1904 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_574
timestamp 1680363874
transform 1 0 1912 0 1 370
box -8 -3 104 105
use FILL  FILL_10384
timestamp 1680363874
transform 1 0 2008 0 1 370
box -8 -3 16 105
use FILL  FILL_10385
timestamp 1680363874
transform 1 0 2016 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_382
timestamp 1680363874
transform 1 0 2024 0 1 370
box -8 -3 46 105
use FILL  FILL_10393
timestamp 1680363874
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_10400
timestamp 1680363874
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_10402
timestamp 1680363874
transform 1 0 2080 0 1 370
box -8 -3 16 105
use INVX2  INVX2_664
timestamp 1680363874
transform -1 0 2104 0 1 370
box -9 -3 26 105
use FILL  FILL_10403
timestamp 1680363874
transform 1 0 2104 0 1 370
box -8 -3 16 105
use FILL  FILL_10408
timestamp 1680363874
transform 1 0 2112 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_419
timestamp 1680363874
transform 1 0 2120 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_8418
timestamp 1680363874
transform 1 0 2180 0 1 375
box -3 -3 3 3
use FILL  FILL_10410
timestamp 1680363874
transform 1 0 2160 0 1 370
box -8 -3 16 105
use FILL  FILL_10411
timestamp 1680363874
transform 1 0 2168 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8419
timestamp 1680363874
transform 1 0 2220 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_420
timestamp 1680363874
transform 1 0 2176 0 1 370
box -8 -3 46 105
use FILL  FILL_10417
timestamp 1680363874
transform 1 0 2216 0 1 370
box -8 -3 16 105
use FILL  FILL_10418
timestamp 1680363874
transform 1 0 2224 0 1 370
box -8 -3 16 105
use FILL  FILL_10419
timestamp 1680363874
transform 1 0 2232 0 1 370
box -8 -3 16 105
use FILL  FILL_10420
timestamp 1680363874
transform 1 0 2240 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_575
timestamp 1680363874
transform -1 0 2344 0 1 370
box -8 -3 104 105
use INVX2  INVX2_666
timestamp 1680363874
transform -1 0 2360 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_576
timestamp 1680363874
transform -1 0 2456 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_577
timestamp 1680363874
transform 1 0 2456 0 1 370
box -8 -3 104 105
use FILL  FILL_10421
timestamp 1680363874
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_10422
timestamp 1680363874
transform 1 0 2560 0 1 370
box -8 -3 16 105
use FILL  FILL_10423
timestamp 1680363874
transform 1 0 2568 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8420
timestamp 1680363874
transform 1 0 2644 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_578
timestamp 1680363874
transform 1 0 2576 0 1 370
box -8 -3 104 105
use FILL  FILL_10424
timestamp 1680363874
transform 1 0 2672 0 1 370
box -8 -3 16 105
use FILL  FILL_10425
timestamp 1680363874
transform 1 0 2680 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8421
timestamp 1680363874
transform 1 0 2700 0 1 375
box -3 -3 3 3
use INVX2  INVX2_667
timestamp 1680363874
transform 1 0 2688 0 1 370
box -9 -3 26 105
use FILL  FILL_10426
timestamp 1680363874
transform 1 0 2704 0 1 370
box -8 -3 16 105
use FILL  FILL_10427
timestamp 1680363874
transform 1 0 2712 0 1 370
box -8 -3 16 105
use FILL  FILL_10428
timestamp 1680363874
transform 1 0 2720 0 1 370
box -8 -3 16 105
use FILL  FILL_10440
timestamp 1680363874
transform 1 0 2728 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_177
timestamp 1680363874
transform 1 0 2736 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1680363874
transform 1 0 2768 0 1 370
box -8 -3 34 105
use FILL  FILL_10442
timestamp 1680363874
transform 1 0 2800 0 1 370
box -8 -3 16 105
use FILL  FILL_10443
timestamp 1680363874
transform 1 0 2808 0 1 370
box -8 -3 16 105
use FILL  FILL_10444
timestamp 1680363874
transform 1 0 2816 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_179
timestamp 1680363874
transform -1 0 2856 0 1 370
box -8 -3 34 105
use FILL  FILL_10445
timestamp 1680363874
transform 1 0 2856 0 1 370
box -8 -3 16 105
use FILL  FILL_10446
timestamp 1680363874
transform 1 0 2864 0 1 370
box -8 -3 16 105
use FILL  FILL_10447
timestamp 1680363874
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_10448
timestamp 1680363874
transform 1 0 2880 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_384
timestamp 1680363874
transform -1 0 2928 0 1 370
box -8 -3 46 105
use INVX2  INVX2_670
timestamp 1680363874
transform 1 0 2928 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_582
timestamp 1680363874
transform -1 0 3040 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_583
timestamp 1680363874
transform 1 0 3040 0 1 370
box -8 -3 104 105
use INVX2  INVX2_671
timestamp 1680363874
transform -1 0 3152 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_385
timestamp 1680363874
transform -1 0 3192 0 1 370
box -8 -3 46 105
use FILL  FILL_10449
timestamp 1680363874
transform 1 0 3192 0 1 370
box -8 -3 16 105
use FILL  FILL_10450
timestamp 1680363874
transform 1 0 3200 0 1 370
box -8 -3 16 105
use FILL  FILL_10451
timestamp 1680363874
transform 1 0 3208 0 1 370
box -8 -3 16 105
use FILL  FILL_10452
timestamp 1680363874
transform 1 0 3216 0 1 370
box -8 -3 16 105
use FILL  FILL_10453
timestamp 1680363874
transform 1 0 3224 0 1 370
box -8 -3 16 105
use FILL  FILL_10454
timestamp 1680363874
transform 1 0 3232 0 1 370
box -8 -3 16 105
use FILL  FILL_10473
timestamp 1680363874
transform 1 0 3240 0 1 370
box -8 -3 16 105
use FILL  FILL_10475
timestamp 1680363874
transform 1 0 3248 0 1 370
box -8 -3 16 105
use FILL  FILL_10477
timestamp 1680363874
transform 1 0 3256 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_389
timestamp 1680363874
transform 1 0 3264 0 1 370
box -8 -3 46 105
use FILL  FILL_10478
timestamp 1680363874
transform 1 0 3304 0 1 370
box -8 -3 16 105
use FILL  FILL_10479
timestamp 1680363874
transform 1 0 3312 0 1 370
box -8 -3 16 105
use FILL  FILL_10480
timestamp 1680363874
transform 1 0 3320 0 1 370
box -8 -3 16 105
use FILL  FILL_10481
timestamp 1680363874
transform 1 0 3328 0 1 370
box -8 -3 16 105
use FILL  FILL_10482
timestamp 1680363874
transform 1 0 3336 0 1 370
box -8 -3 16 105
use FILL  FILL_10483
timestamp 1680363874
transform 1 0 3344 0 1 370
box -8 -3 16 105
use FILL  FILL_10484
timestamp 1680363874
transform 1 0 3352 0 1 370
box -8 -3 16 105
use FILL  FILL_10485
timestamp 1680363874
transform 1 0 3360 0 1 370
box -8 -3 16 105
use FILL  FILL_10486
timestamp 1680363874
transform 1 0 3368 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_390
timestamp 1680363874
transform 1 0 3376 0 1 370
box -8 -3 46 105
use FILL  FILL_10488
timestamp 1680363874
transform 1 0 3416 0 1 370
box -8 -3 16 105
use INVX2  INVX2_674
timestamp 1680363874
transform 1 0 3424 0 1 370
box -9 -3 26 105
use FILL  FILL_10490
timestamp 1680363874
transform 1 0 3440 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_586
timestamp 1680363874
transform -1 0 3544 0 1 370
box -8 -3 104 105
use FILL  FILL_10491
timestamp 1680363874
transform 1 0 3544 0 1 370
box -8 -3 16 105
use FILL  FILL_10492
timestamp 1680363874
transform 1 0 3552 0 1 370
box -8 -3 16 105
use INVX2  INVX2_675
timestamp 1680363874
transform 1 0 3560 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_587
timestamp 1680363874
transform -1 0 3672 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_8422
timestamp 1680363874
transform 1 0 3716 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_424
timestamp 1680363874
transform -1 0 3712 0 1 370
box -8 -3 46 105
use FILL  FILL_10493
timestamp 1680363874
transform 1 0 3712 0 1 370
box -8 -3 16 105
use FILL  FILL_10502
timestamp 1680363874
transform 1 0 3720 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8423
timestamp 1680363874
transform 1 0 3748 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_589
timestamp 1680363874
transform 1 0 3728 0 1 370
box -8 -3 104 105
use FILL  FILL_10504
timestamp 1680363874
transform 1 0 3824 0 1 370
box -8 -3 16 105
use FILL  FILL_10505
timestamp 1680363874
transform 1 0 3832 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_590
timestamp 1680363874
transform 1 0 3840 0 1 370
box -8 -3 104 105
use FILL  FILL_10506
timestamp 1680363874
transform 1 0 3936 0 1 370
box -8 -3 16 105
use FILL  FILL_10507
timestamp 1680363874
transform 1 0 3944 0 1 370
box -8 -3 16 105
use INVX2  INVX2_677
timestamp 1680363874
transform 1 0 3952 0 1 370
box -9 -3 26 105
use FILL  FILL_10508
timestamp 1680363874
transform 1 0 3968 0 1 370
box -8 -3 16 105
use FILL  FILL_10509
timestamp 1680363874
transform 1 0 3976 0 1 370
box -8 -3 16 105
use FILL  FILL_10516
timestamp 1680363874
transform 1 0 3984 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_426
timestamp 1680363874
transform 1 0 3992 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_8424
timestamp 1680363874
transform 1 0 4108 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_591
timestamp 1680363874
transform -1 0 4128 0 1 370
box -8 -3 104 105
use FILL  FILL_10518
timestamp 1680363874
transform 1 0 4128 0 1 370
box -8 -3 16 105
use FILL  FILL_10519
timestamp 1680363874
transform 1 0 4136 0 1 370
box -8 -3 16 105
use FILL  FILL_10520
timestamp 1680363874
transform 1 0 4144 0 1 370
box -8 -3 16 105
use FILL  FILL_10521
timestamp 1680363874
transform 1 0 4152 0 1 370
box -8 -3 16 105
use FILL  FILL_10522
timestamp 1680363874
transform 1 0 4160 0 1 370
box -8 -3 16 105
use INVX2  INVX2_681
timestamp 1680363874
transform -1 0 4184 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_8425
timestamp 1680363874
transform 1 0 4196 0 1 375
box -3 -3 3 3
use FILL  FILL_10523
timestamp 1680363874
transform 1 0 4184 0 1 370
box -8 -3 16 105
use FILL  FILL_10524
timestamp 1680363874
transform 1 0 4192 0 1 370
box -8 -3 16 105
use FILL  FILL_10525
timestamp 1680363874
transform 1 0 4200 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_427
timestamp 1680363874
transform 1 0 4208 0 1 370
box -8 -3 46 105
use FILL  FILL_10526
timestamp 1680363874
transform 1 0 4248 0 1 370
box -8 -3 16 105
use FILL  FILL_10532
timestamp 1680363874
transform 1 0 4256 0 1 370
box -8 -3 16 105
use FILL  FILL_10533
timestamp 1680363874
transform 1 0 4264 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8426
timestamp 1680363874
transform 1 0 4284 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_400
timestamp 1680363874
transform 1 0 4272 0 1 370
box -8 -3 46 105
use FILL  FILL_10534
timestamp 1680363874
transform 1 0 4312 0 1 370
box -8 -3 16 105
use FILL  FILL_10535
timestamp 1680363874
transform 1 0 4320 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8427
timestamp 1680363874
transform 1 0 4340 0 1 375
box -3 -3 3 3
use FILL  FILL_10536
timestamp 1680363874
transform 1 0 4328 0 1 370
box -8 -3 16 105
use FILL  FILL_10537
timestamp 1680363874
transform 1 0 4336 0 1 370
box -8 -3 16 105
use FILL  FILL_10539
timestamp 1680363874
transform 1 0 4344 0 1 370
box -8 -3 16 105
use FILL  FILL_10541
timestamp 1680363874
transform 1 0 4352 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8428
timestamp 1680363874
transform 1 0 4436 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_593
timestamp 1680363874
transform -1 0 4456 0 1 370
box -8 -3 104 105
use FILL  FILL_10542
timestamp 1680363874
transform 1 0 4456 0 1 370
box -8 -3 16 105
use FILL  FILL_10543
timestamp 1680363874
transform 1 0 4464 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8429
timestamp 1680363874
transform 1 0 4532 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8430
timestamp 1680363874
transform 1 0 4572 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_594
timestamp 1680363874
transform -1 0 4568 0 1 370
box -8 -3 104 105
use FILL  FILL_10544
timestamp 1680363874
transform 1 0 4568 0 1 370
box -8 -3 16 105
use FILL  FILL_10556
timestamp 1680363874
transform 1 0 4576 0 1 370
box -8 -3 16 105
use FILL  FILL_10558
timestamp 1680363874
transform 1 0 4584 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_431
timestamp 1680363874
transform 1 0 4592 0 1 370
box -8 -3 46 105
use FILL  FILL_10560
timestamp 1680363874
transform 1 0 4632 0 1 370
box -8 -3 16 105
use FILL  FILL_10561
timestamp 1680363874
transform 1 0 4640 0 1 370
box -8 -3 16 105
use FILL  FILL_10564
timestamp 1680363874
transform 1 0 4648 0 1 370
box -8 -3 16 105
use FILL  FILL_10566
timestamp 1680363874
transform 1 0 4656 0 1 370
box -8 -3 16 105
use FILL  FILL_10568
timestamp 1680363874
transform 1 0 4664 0 1 370
box -8 -3 16 105
use FILL  FILL_10570
timestamp 1680363874
transform 1 0 4672 0 1 370
box -8 -3 16 105
use FILL  FILL_10572
timestamp 1680363874
transform 1 0 4680 0 1 370
box -8 -3 16 105
use FILL  FILL_10573
timestamp 1680363874
transform 1 0 4688 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_595
timestamp 1680363874
transform -1 0 4792 0 1 370
box -8 -3 104 105
use FILL  FILL_10574
timestamp 1680363874
transform 1 0 4792 0 1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_87
timestamp 1680363874
transform 1 0 4827 0 1 370
box -10 -3 10 3
use M3_M2  M3_M2_8501
timestamp 1680363874
transform 1 0 84 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8502
timestamp 1680363874
transform 1 0 140 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9393
timestamp 1680363874
transform 1 0 164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9521
timestamp 1680363874
transform 1 0 84 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9522
timestamp 1680363874
transform 1 0 132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8449
timestamp 1680363874
transform 1 0 260 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9394
timestamp 1680363874
transform 1 0 236 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9395
timestamp 1680363874
transform 1 0 252 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8531
timestamp 1680363874
transform 1 0 236 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9523
timestamp 1680363874
transform 1 0 244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9524
timestamp 1680363874
transform 1 0 260 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8532
timestamp 1680363874
transform 1 0 268 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9525
timestamp 1680363874
transform 1 0 276 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8450
timestamp 1680363874
transform 1 0 284 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8469
timestamp 1680363874
transform 1 0 324 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9396
timestamp 1680363874
transform 1 0 316 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8533
timestamp 1680363874
transform 1 0 308 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8431
timestamp 1680363874
transform 1 0 356 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8451
timestamp 1680363874
transform 1 0 372 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8470
timestamp 1680363874
transform 1 0 348 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9397
timestamp 1680363874
transform 1 0 348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9398
timestamp 1680363874
transform 1 0 364 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8534
timestamp 1680363874
transform 1 0 348 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9399
timestamp 1680363874
transform 1 0 388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9526
timestamp 1680363874
transform 1 0 372 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8535
timestamp 1680363874
transform 1 0 380 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9527
timestamp 1680363874
transform 1 0 388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9400
timestamp 1680363874
transform 1 0 404 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8452
timestamp 1680363874
transform 1 0 484 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9401
timestamp 1680363874
transform 1 0 436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9528
timestamp 1680363874
transform 1 0 484 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8503
timestamp 1680363874
transform 1 0 532 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9529
timestamp 1680363874
transform 1 0 532 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8471
timestamp 1680363874
transform 1 0 596 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9402
timestamp 1680363874
transform 1 0 548 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8504
timestamp 1680363874
transform 1 0 572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8505
timestamp 1680363874
transform 1 0 636 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8432
timestamp 1680363874
transform 1 0 652 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8453
timestamp 1680363874
transform 1 0 660 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9403
timestamp 1680363874
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9404
timestamp 1680363874
transform 1 0 660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9530
timestamp 1680363874
transform 1 0 596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9531
timestamp 1680363874
transform 1 0 628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9532
timestamp 1680363874
transform 1 0 652 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8536
timestamp 1680363874
transform 1 0 660 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9533
timestamp 1680363874
transform 1 0 668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9405
timestamp 1680363874
transform 1 0 684 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8472
timestamp 1680363874
transform 1 0 708 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9406
timestamp 1680363874
transform 1 0 708 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8506
timestamp 1680363874
transform 1 0 716 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9407
timestamp 1680363874
transform 1 0 724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9534
timestamp 1680363874
transform 1 0 700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9535
timestamp 1680363874
transform 1 0 716 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8507
timestamp 1680363874
transform 1 0 732 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9408
timestamp 1680363874
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9536
timestamp 1680363874
transform 1 0 732 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8607
timestamp 1680363874
transform 1 0 740 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9409
timestamp 1680363874
transform 1 0 780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9537
timestamp 1680363874
transform 1 0 772 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8537
timestamp 1680363874
transform 1 0 780 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9538
timestamp 1680363874
transform 1 0 788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8565
timestamp 1680363874
transform 1 0 788 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9670
timestamp 1680363874
transform 1 0 796 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8608
timestamp 1680363874
transform 1 0 796 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9539
timestamp 1680363874
transform 1 0 844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9674
timestamp 1680363874
transform 1 0 852 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_9410
timestamp 1680363874
transform 1 0 884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9671
timestamp 1680363874
transform 1 0 892 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8454
timestamp 1680363874
transform 1 0 916 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9390
timestamp 1680363874
transform 1 0 932 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9540
timestamp 1680363874
transform 1 0 940 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8566
timestamp 1680363874
transform 1 0 940 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8473
timestamp 1680363874
transform 1 0 988 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8508
timestamp 1680363874
transform 1 0 980 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9411
timestamp 1680363874
transform 1 0 988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9541
timestamp 1680363874
transform 1 0 964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9542
timestamp 1680363874
transform 1 0 980 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8433
timestamp 1680363874
transform 1 0 1020 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8434
timestamp 1680363874
transform 1 0 1044 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8474
timestamp 1680363874
transform 1 0 1036 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9412
timestamp 1680363874
transform 1 0 1004 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9413
timestamp 1680363874
transform 1 0 1092 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8509
timestamp 1680363874
transform 1 0 1108 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8455
timestamp 1680363874
transform 1 0 1172 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9414
timestamp 1680363874
transform 1 0 1116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9415
timestamp 1680363874
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9416
timestamp 1680363874
transform 1 0 1140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9417
timestamp 1680363874
transform 1 0 1164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9418
timestamp 1680363874
transform 1 0 1180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9543
timestamp 1680363874
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9544
timestamp 1680363874
transform 1 0 1084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9545
timestamp 1680363874
transform 1 0 1100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9546
timestamp 1680363874
transform 1 0 1108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9547
timestamp 1680363874
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9548
timestamp 1680363874
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9549
timestamp 1680363874
transform 1 0 1156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9550
timestamp 1680363874
transform 1 0 1172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8567
timestamp 1680363874
transform 1 0 1100 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8568
timestamp 1680363874
transform 1 0 1132 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8569
timestamp 1680363874
transform 1 0 1156 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8609
timestamp 1680363874
transform 1 0 1140 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8630
timestamp 1680363874
transform 1 0 1180 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9419
timestamp 1680363874
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8610
timestamp 1680363874
transform 1 0 1212 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9551
timestamp 1680363874
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9420
timestamp 1680363874
transform 1 0 1244 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8456
timestamp 1680363874
transform 1 0 1324 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9421
timestamp 1680363874
transform 1 0 1292 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8510
timestamp 1680363874
transform 1 0 1300 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9422
timestamp 1680363874
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9423
timestamp 1680363874
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9552
timestamp 1680363874
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9553
timestamp 1680363874
transform 1 0 1308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9554
timestamp 1680363874
transform 1 0 1324 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8475
timestamp 1680363874
transform 1 0 1348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8435
timestamp 1680363874
transform 1 0 1372 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8457
timestamp 1680363874
transform 1 0 1388 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8476
timestamp 1680363874
transform 1 0 1404 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9424
timestamp 1680363874
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9425
timestamp 1680363874
transform 1 0 1388 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8511
timestamp 1680363874
transform 1 0 1396 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9426
timestamp 1680363874
transform 1 0 1404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9555
timestamp 1680363874
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9556
timestamp 1680363874
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9557
timestamp 1680363874
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8611
timestamp 1680363874
transform 1 0 1380 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8436
timestamp 1680363874
transform 1 0 1420 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8437
timestamp 1680363874
transform 1 0 1436 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8458
timestamp 1680363874
transform 1 0 1484 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8477
timestamp 1680363874
transform 1 0 1516 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9427
timestamp 1680363874
transform 1 0 1420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9428
timestamp 1680363874
transform 1 0 1436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9558
timestamp 1680363874
transform 1 0 1484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9559
timestamp 1680363874
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8438
timestamp 1680363874
transform 1 0 1620 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8478
timestamp 1680363874
transform 1 0 1540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8479
timestamp 1680363874
transform 1 0 1588 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9429
timestamp 1680363874
transform 1 0 1540 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8512
timestamp 1680363874
transform 1 0 1564 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8538
timestamp 1680363874
transform 1 0 1540 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9560
timestamp 1680363874
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8539
timestamp 1680363874
transform 1 0 1612 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9430
timestamp 1680363874
transform 1 0 1628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9561
timestamp 1680363874
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8570
timestamp 1680363874
transform 1 0 1604 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8459
timestamp 1680363874
transform 1 0 1644 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8460
timestamp 1680363874
transform 1 0 1660 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8612
timestamp 1680363874
transform 1 0 1636 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8480
timestamp 1680363874
transform 1 0 1660 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8513
timestamp 1680363874
transform 1 0 1652 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9431
timestamp 1680363874
transform 1 0 1660 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8514
timestamp 1680363874
transform 1 0 1668 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8439
timestamp 1680363874
transform 1 0 1692 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9432
timestamp 1680363874
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9433
timestamp 1680363874
transform 1 0 1692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9562
timestamp 1680363874
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8540
timestamp 1680363874
transform 1 0 1660 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9563
timestamp 1680363874
transform 1 0 1668 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8571
timestamp 1680363874
transform 1 0 1652 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8613
timestamp 1680363874
transform 1 0 1668 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9564
timestamp 1680363874
transform 1 0 1732 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8481
timestamp 1680363874
transform 1 0 1796 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9434
timestamp 1680363874
transform 1 0 1796 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9565
timestamp 1680363874
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9435
timestamp 1680363874
transform 1 0 1836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9566
timestamp 1680363874
transform 1 0 1828 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9567
timestamp 1680363874
transform 1 0 1844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9568
timestamp 1680363874
transform 1 0 1852 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8572
timestamp 1680363874
transform 1 0 1828 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8573
timestamp 1680363874
transform 1 0 1852 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8614
timestamp 1680363874
transform 1 0 1844 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9436
timestamp 1680363874
transform 1 0 1876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9437
timestamp 1680363874
transform 1 0 1884 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8541
timestamp 1680363874
transform 1 0 1876 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9438
timestamp 1680363874
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9569
timestamp 1680363874
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9570
timestamp 1680363874
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8542
timestamp 1680363874
transform 1 0 1956 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9439
timestamp 1680363874
transform 1 0 1972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9571
timestamp 1680363874
transform 1 0 1964 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8482
timestamp 1680363874
transform 1 0 2012 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9440
timestamp 1680363874
transform 1 0 1996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9441
timestamp 1680363874
transform 1 0 2012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9572
timestamp 1680363874
transform 1 0 1980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9573
timestamp 1680363874
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8574
timestamp 1680363874
transform 1 0 1972 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8575
timestamp 1680363874
transform 1 0 2004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8615
timestamp 1680363874
transform 1 0 1980 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8576
timestamp 1680363874
transform 1 0 2036 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8515
timestamp 1680363874
transform 1 0 2108 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8516
timestamp 1680363874
transform 1 0 2140 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9442
timestamp 1680363874
transform 1 0 2156 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8440
timestamp 1680363874
transform 1 0 2172 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9443
timestamp 1680363874
transform 1 0 2172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9574
timestamp 1680363874
transform 1 0 2164 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8543
timestamp 1680363874
transform 1 0 2172 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9575
timestamp 1680363874
transform 1 0 2188 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8441
timestamp 1680363874
transform 1 0 2212 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8461
timestamp 1680363874
transform 1 0 2228 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9444
timestamp 1680363874
transform 1 0 2212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9445
timestamp 1680363874
transform 1 0 2228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9576
timestamp 1680363874
transform 1 0 2204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9577
timestamp 1680363874
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8544
timestamp 1680363874
transform 1 0 2228 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9578
timestamp 1680363874
transform 1 0 2236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9446
timestamp 1680363874
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8483
timestamp 1680363874
transform 1 0 2284 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8484
timestamp 1680363874
transform 1 0 2332 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9447
timestamp 1680363874
transform 1 0 2284 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8517
timestamp 1680363874
transform 1 0 2308 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9579
timestamp 1680363874
transform 1 0 2308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9580
timestamp 1680363874
transform 1 0 2364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9448
timestamp 1680363874
transform 1 0 2396 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8485
timestamp 1680363874
transform 1 0 2500 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8462
timestamp 1680363874
transform 1 0 2516 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9391
timestamp 1680363874
transform 1 0 2516 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9449
timestamp 1680363874
transform 1 0 2500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9450
timestamp 1680363874
transform 1 0 2508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9581
timestamp 1680363874
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9582
timestamp 1680363874
transform 1 0 2476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9583
timestamp 1680363874
transform 1 0 2484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9584
timestamp 1680363874
transform 1 0 2500 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8577
timestamp 1680363874
transform 1 0 2444 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8578
timestamp 1680363874
transform 1 0 2484 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8616
timestamp 1680363874
transform 1 0 2476 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9451
timestamp 1680363874
transform 1 0 2532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9452
timestamp 1680363874
transform 1 0 2620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9453
timestamp 1680363874
transform 1 0 2636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9585
timestamp 1680363874
transform 1 0 2580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9586
timestamp 1680363874
transform 1 0 2620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9587
timestamp 1680363874
transform 1 0 2628 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8579
timestamp 1680363874
transform 1 0 2580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8545
timestamp 1680363874
transform 1 0 2636 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9588
timestamp 1680363874
transform 1 0 2644 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8631
timestamp 1680363874
transform 1 0 2644 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8639
timestamp 1680363874
transform 1 0 2612 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8640
timestamp 1680363874
transform 1 0 2628 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9454
timestamp 1680363874
transform 1 0 2660 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8546
timestamp 1680363874
transform 1 0 2660 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8580
timestamp 1680363874
transform 1 0 2668 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9455
timestamp 1680363874
transform 1 0 2676 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8486
timestamp 1680363874
transform 1 0 2700 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9456
timestamp 1680363874
transform 1 0 2716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9457
timestamp 1680363874
transform 1 0 2724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9458
timestamp 1680363874
transform 1 0 2732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9589
timestamp 1680363874
transform 1 0 2684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9590
timestamp 1680363874
transform 1 0 2700 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8581
timestamp 1680363874
transform 1 0 2684 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8617
timestamp 1680363874
transform 1 0 2676 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8547
timestamp 1680363874
transform 1 0 2724 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8518
timestamp 1680363874
transform 1 0 2748 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9591
timestamp 1680363874
transform 1 0 2740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9672
timestamp 1680363874
transform 1 0 2748 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9673
timestamp 1680363874
transform 1 0 2780 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9459
timestamp 1680363874
transform 1 0 2804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9592
timestamp 1680363874
transform 1 0 2820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9593
timestamp 1680363874
transform 1 0 2828 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8582
timestamp 1680363874
transform 1 0 2828 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8442
timestamp 1680363874
transform 1 0 2900 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8487
timestamp 1680363874
transform 1 0 2868 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8488
timestamp 1680363874
transform 1 0 2916 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8489
timestamp 1680363874
transform 1 0 2996 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9460
timestamp 1680363874
transform 1 0 2868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9461
timestamp 1680363874
transform 1 0 2884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9462
timestamp 1680363874
transform 1 0 2892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9594
timestamp 1680363874
transform 1 0 2860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9595
timestamp 1680363874
transform 1 0 2876 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8548
timestamp 1680363874
transform 1 0 2884 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9463
timestamp 1680363874
transform 1 0 2996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9596
timestamp 1680363874
transform 1 0 2900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9597
timestamp 1680363874
transform 1 0 2908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9598
timestamp 1680363874
transform 1 0 2916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8549
timestamp 1680363874
transform 1 0 2932 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9599
timestamp 1680363874
transform 1 0 2948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9600
timestamp 1680363874
transform 1 0 3012 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8583
timestamp 1680363874
transform 1 0 2908 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8584
timestamp 1680363874
transform 1 0 2948 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8490
timestamp 1680363874
transform 1 0 3028 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9464
timestamp 1680363874
transform 1 0 3028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9392
timestamp 1680363874
transform 1 0 3076 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8519
timestamp 1680363874
transform 1 0 3076 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8463
timestamp 1680363874
transform 1 0 3100 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9465
timestamp 1680363874
transform 1 0 3084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9466
timestamp 1680363874
transform 1 0 3100 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8550
timestamp 1680363874
transform 1 0 3084 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9601
timestamp 1680363874
transform 1 0 3092 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9602
timestamp 1680363874
transform 1 0 3108 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8585
timestamp 1680363874
transform 1 0 3116 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8632
timestamp 1680363874
transform 1 0 3108 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8641
timestamp 1680363874
transform 1 0 3092 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9603
timestamp 1680363874
transform 1 0 3140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9604
timestamp 1680363874
transform 1 0 3148 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8618
timestamp 1680363874
transform 1 0 3148 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8443
timestamp 1680363874
transform 1 0 3188 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8491
timestamp 1680363874
transform 1 0 3188 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9467
timestamp 1680363874
transform 1 0 3180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9468
timestamp 1680363874
transform 1 0 3220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9469
timestamp 1680363874
transform 1 0 3228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9605
timestamp 1680363874
transform 1 0 3172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9606
timestamp 1680363874
transform 1 0 3188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9607
timestamp 1680363874
transform 1 0 3196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9608
timestamp 1680363874
transform 1 0 3212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9609
timestamp 1680363874
transform 1 0 3228 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8586
timestamp 1680363874
transform 1 0 3220 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8619
timestamp 1680363874
transform 1 0 3228 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8633
timestamp 1680363874
transform 1 0 3204 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8444
timestamp 1680363874
transform 1 0 3268 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9470
timestamp 1680363874
transform 1 0 3284 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8520
timestamp 1680363874
transform 1 0 3332 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8492
timestamp 1680363874
transform 1 0 3372 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9610
timestamp 1680363874
transform 1 0 3268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9611
timestamp 1680363874
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9612
timestamp 1680363874
transform 1 0 3364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9613
timestamp 1680363874
transform 1 0 3372 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8587
timestamp 1680363874
transform 1 0 3268 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8588
timestamp 1680363874
transform 1 0 3308 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8620
timestamp 1680363874
transform 1 0 3364 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8634
timestamp 1680363874
transform 1 0 3324 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8642
timestamp 1680363874
transform 1 0 3292 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8643
timestamp 1680363874
transform 1 0 3316 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8644
timestamp 1680363874
transform 1 0 3340 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9471
timestamp 1680363874
transform 1 0 3388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9472
timestamp 1680363874
transform 1 0 3404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9473
timestamp 1680363874
transform 1 0 3412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9614
timestamp 1680363874
transform 1 0 3396 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8551
timestamp 1680363874
transform 1 0 3404 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9615
timestamp 1680363874
transform 1 0 3420 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8521
timestamp 1680363874
transform 1 0 3460 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9474
timestamp 1680363874
transform 1 0 3548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9616
timestamp 1680363874
transform 1 0 3460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9617
timestamp 1680363874
transform 1 0 3468 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8552
timestamp 1680363874
transform 1 0 3476 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9618
timestamp 1680363874
transform 1 0 3500 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8589
timestamp 1680363874
transform 1 0 3460 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8590
timestamp 1680363874
transform 1 0 3500 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9475
timestamp 1680363874
transform 1 0 3564 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8522
timestamp 1680363874
transform 1 0 3580 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9619
timestamp 1680363874
transform 1 0 3572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9620
timestamp 1680363874
transform 1 0 3588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8591
timestamp 1680363874
transform 1 0 3572 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8464
timestamp 1680363874
transform 1 0 3676 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8465
timestamp 1680363874
transform 1 0 3708 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9476
timestamp 1680363874
transform 1 0 3636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9477
timestamp 1680363874
transform 1 0 3644 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8523
timestamp 1680363874
transform 1 0 3652 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9478
timestamp 1680363874
transform 1 0 3676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9479
timestamp 1680363874
transform 1 0 3684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9480
timestamp 1680363874
transform 1 0 3700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9481
timestamp 1680363874
transform 1 0 3708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9621
timestamp 1680363874
transform 1 0 3628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9622
timestamp 1680363874
transform 1 0 3636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9623
timestamp 1680363874
transform 1 0 3652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9624
timestamp 1680363874
transform 1 0 3668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9625
timestamp 1680363874
transform 1 0 3676 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9626
timestamp 1680363874
transform 1 0 3692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9627
timestamp 1680363874
transform 1 0 3708 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8621
timestamp 1680363874
transform 1 0 3620 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8592
timestamp 1680363874
transform 1 0 3668 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8645
timestamp 1680363874
transform 1 0 3636 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8622
timestamp 1680363874
transform 1 0 3676 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8635
timestamp 1680363874
transform 1 0 3700 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8646
timestamp 1680363874
transform 1 0 3708 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8553
timestamp 1680363874
transform 1 0 3724 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9628
timestamp 1680363874
transform 1 0 3732 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8493
timestamp 1680363874
transform 1 0 3796 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8494
timestamp 1680363874
transform 1 0 3828 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9482
timestamp 1680363874
transform 1 0 3756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9483
timestamp 1680363874
transform 1 0 3772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9484
timestamp 1680363874
transform 1 0 3796 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9485
timestamp 1680363874
transform 1 0 3804 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8554
timestamp 1680363874
transform 1 0 3756 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8524
timestamp 1680363874
transform 1 0 3812 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9486
timestamp 1680363874
transform 1 0 3820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9487
timestamp 1680363874
transform 1 0 3828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9629
timestamp 1680363874
transform 1 0 3764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9630
timestamp 1680363874
transform 1 0 3780 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9631
timestamp 1680363874
transform 1 0 3796 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8555
timestamp 1680363874
transform 1 0 3804 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9632
timestamp 1680363874
transform 1 0 3812 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8593
timestamp 1680363874
transform 1 0 3796 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8647
timestamp 1680363874
transform 1 0 3788 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8495
timestamp 1680363874
transform 1 0 3852 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8496
timestamp 1680363874
transform 1 0 3892 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9488
timestamp 1680363874
transform 1 0 3868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9489
timestamp 1680363874
transform 1 0 3876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9633
timestamp 1680363874
transform 1 0 3844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9634
timestamp 1680363874
transform 1 0 3860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8623
timestamp 1680363874
transform 1 0 3836 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9675
timestamp 1680363874
transform 1 0 3836 0 1 295
box -2 -2 2 2
use M3_M2  M3_M2_8648
timestamp 1680363874
transform 1 0 3836 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8556
timestamp 1680363874
transform 1 0 3868 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8525
timestamp 1680363874
transform 1 0 3892 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9490
timestamp 1680363874
transform 1 0 3900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9635
timestamp 1680363874
transform 1 0 3876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9636
timestamp 1680363874
transform 1 0 3884 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8636
timestamp 1680363874
transform 1 0 3868 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8649
timestamp 1680363874
transform 1 0 3852 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8650
timestamp 1680363874
transform 1 0 3876 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9637
timestamp 1680363874
transform 1 0 3900 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8594
timestamp 1680363874
transform 1 0 3900 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9491
timestamp 1680363874
transform 1 0 3924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9492
timestamp 1680363874
transform 1 0 3940 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8526
timestamp 1680363874
transform 1 0 3948 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9493
timestamp 1680363874
transform 1 0 3972 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8527
timestamp 1680363874
transform 1 0 3980 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9638
timestamp 1680363874
transform 1 0 3940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9639
timestamp 1680363874
transform 1 0 3956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9640
timestamp 1680363874
transform 1 0 3972 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8595
timestamp 1680363874
transform 1 0 3972 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9494
timestamp 1680363874
transform 1 0 3996 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8528
timestamp 1680363874
transform 1 0 4004 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9495
timestamp 1680363874
transform 1 0 4012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9496
timestamp 1680363874
transform 1 0 4020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9497
timestamp 1680363874
transform 1 0 4036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9641
timestamp 1680363874
transform 1 0 4004 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8557
timestamp 1680363874
transform 1 0 4020 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9642
timestamp 1680363874
transform 1 0 4028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9643
timestamp 1680363874
transform 1 0 4044 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8596
timestamp 1680363874
transform 1 0 3996 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8597
timestamp 1680363874
transform 1 0 4028 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9498
timestamp 1680363874
transform 1 0 4060 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8598
timestamp 1680363874
transform 1 0 4052 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8624
timestamp 1680363874
transform 1 0 4044 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8445
timestamp 1680363874
transform 1 0 4204 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9499
timestamp 1680363874
transform 1 0 4084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9500
timestamp 1680363874
transform 1 0 4172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9501
timestamp 1680363874
transform 1 0 4196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9644
timestamp 1680363874
transform 1 0 4132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9645
timestamp 1680363874
transform 1 0 4164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9646
timestamp 1680363874
transform 1 0 4172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9647
timestamp 1680363874
transform 1 0 4188 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8558
timestamp 1680363874
transform 1 0 4196 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9648
timestamp 1680363874
transform 1 0 4204 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8625
timestamp 1680363874
transform 1 0 4172 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9649
timestamp 1680363874
transform 1 0 4220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9650
timestamp 1680363874
transform 1 0 4236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8626
timestamp 1680363874
transform 1 0 4220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8497
timestamp 1680363874
transform 1 0 4284 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9502
timestamp 1680363874
transform 1 0 4260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9503
timestamp 1680363874
transform 1 0 4268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9504
timestamp 1680363874
transform 1 0 4284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9651
timestamp 1680363874
transform 1 0 4260 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8559
timestamp 1680363874
transform 1 0 4268 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9505
timestamp 1680363874
transform 1 0 4316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9506
timestamp 1680363874
transform 1 0 4332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9652
timestamp 1680363874
transform 1 0 4276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9653
timestamp 1680363874
transform 1 0 4292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9654
timestamp 1680363874
transform 1 0 4308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9655
timestamp 1680363874
transform 1 0 4324 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8599
timestamp 1680363874
transform 1 0 4260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8600
timestamp 1680363874
transform 1 0 4300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8627
timestamp 1680363874
transform 1 0 4292 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8529
timestamp 1680363874
transform 1 0 4364 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8498
timestamp 1680363874
transform 1 0 4420 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9507
timestamp 1680363874
transform 1 0 4412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9508
timestamp 1680363874
transform 1 0 4428 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8560
timestamp 1680363874
transform 1 0 4412 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8530
timestamp 1680363874
transform 1 0 4444 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9509
timestamp 1680363874
transform 1 0 4452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9656
timestamp 1680363874
transform 1 0 4420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9657
timestamp 1680363874
transform 1 0 4436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9658
timestamp 1680363874
transform 1 0 4444 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8601
timestamp 1680363874
transform 1 0 4404 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8602
timestamp 1680363874
transform 1 0 4436 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9659
timestamp 1680363874
transform 1 0 4468 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8628
timestamp 1680363874
transform 1 0 4468 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8446
timestamp 1680363874
transform 1 0 4492 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8447
timestamp 1680363874
transform 1 0 4516 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9510
timestamp 1680363874
transform 1 0 4484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9511
timestamp 1680363874
transform 1 0 4492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9512
timestamp 1680363874
transform 1 0 4508 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8561
timestamp 1680363874
transform 1 0 4492 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9513
timestamp 1680363874
transform 1 0 4524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9660
timestamp 1680363874
transform 1 0 4500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9661
timestamp 1680363874
transform 1 0 4516 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8448
timestamp 1680363874
transform 1 0 4548 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8466
timestamp 1680363874
transform 1 0 4540 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8467
timestamp 1680363874
transform 1 0 4556 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8499
timestamp 1680363874
transform 1 0 4556 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9514
timestamp 1680363874
transform 1 0 4548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9662
timestamp 1680363874
transform 1 0 4532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9663
timestamp 1680363874
transform 1 0 4556 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8603
timestamp 1680363874
transform 1 0 4540 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9515
timestamp 1680363874
transform 1 0 4572 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8562
timestamp 1680363874
transform 1 0 4572 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9664
timestamp 1680363874
transform 1 0 4580 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8604
timestamp 1680363874
transform 1 0 4580 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9516
timestamp 1680363874
transform 1 0 4596 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8468
timestamp 1680363874
transform 1 0 4620 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9517
timestamp 1680363874
transform 1 0 4612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9518
timestamp 1680363874
transform 1 0 4628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9519
timestamp 1680363874
transform 1 0 4636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9665
timestamp 1680363874
transform 1 0 4620 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8563
timestamp 1680363874
transform 1 0 4628 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9666
timestamp 1680363874
transform 1 0 4636 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8629
timestamp 1680363874
transform 1 0 4636 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8637
timestamp 1680363874
transform 1 0 4612 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8638
timestamp 1680363874
transform 1 0 4660 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8500
timestamp 1680363874
transform 1 0 4708 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9520
timestamp 1680363874
transform 1 0 4708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9667
timestamp 1680363874
transform 1 0 4692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9668
timestamp 1680363874
transform 1 0 4732 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8564
timestamp 1680363874
transform 1 0 4780 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9669
timestamp 1680363874
transform 1 0 4788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8605
timestamp 1680363874
transform 1 0 4692 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8606
timestamp 1680363874
transform 1 0 4732 0 1 315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_88
timestamp 1680363874
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_10221
timestamp 1680363874
transform 1 0 72 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_565
timestamp 1680363874
transform -1 0 176 0 -1 370
box -8 -3 104 105
use FILL  FILL_10222
timestamp 1680363874
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_10224
timestamp 1680363874
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10226
timestamp 1680363874
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_10227
timestamp 1680363874
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_10228
timestamp 1680363874
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_10230
timestamp 1680363874
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_10232
timestamp 1680363874
transform 1 0 224 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_402
timestamp 1680363874
transform 1 0 232 0 -1 370
box -8 -3 46 105
use FILL  FILL_10233
timestamp 1680363874
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_10234
timestamp 1680363874
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_10236
timestamp 1680363874
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_10238
timestamp 1680363874
transform 1 0 296 0 -1 370
box -8 -3 16 105
use FILL  FILL_10240
timestamp 1680363874
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_10242
timestamp 1680363874
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_10244
timestamp 1680363874
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_10246
timestamp 1680363874
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_10248
timestamp 1680363874
transform 1 0 336 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_404
timestamp 1680363874
transform 1 0 344 0 -1 370
box -8 -3 46 105
use FILL  FILL_10264
timestamp 1680363874
transform 1 0 384 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_653
timestamp 1680363874
transform -1 0 408 0 -1 370
box -9 -3 26 105
use FILL  FILL_10265
timestamp 1680363874
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_10266
timestamp 1680363874
transform 1 0 416 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_567
timestamp 1680363874
transform 1 0 424 0 -1 370
box -8 -3 104 105
use FILL  FILL_10267
timestamp 1680363874
transform 1 0 520 0 -1 370
box -8 -3 16 105
use FILL  FILL_10268
timestamp 1680363874
transform 1 0 528 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_568
timestamp 1680363874
transform 1 0 536 0 -1 370
box -8 -3 104 105
use FILL  FILL_10269
timestamp 1680363874
transform 1 0 632 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_405
timestamp 1680363874
transform -1 0 680 0 -1 370
box -8 -3 46 105
use FILL  FILL_10270
timestamp 1680363874
transform 1 0 680 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_406
timestamp 1680363874
transform 1 0 688 0 -1 370
box -8 -3 46 105
use FILL  FILL_10277
timestamp 1680363874
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_10279
timestamp 1680363874
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_10281
timestamp 1680363874
transform 1 0 744 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_375
timestamp 1680363874
transform 1 0 752 0 -1 370
box -8 -3 46 105
use FILL  FILL_10285
timestamp 1680363874
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_10286
timestamp 1680363874
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_10287
timestamp 1680363874
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_10288
timestamp 1680363874
transform 1 0 816 0 -1 370
box -8 -3 16 105
use FILL  FILL_10289
timestamp 1680363874
transform 1 0 824 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8651
timestamp 1680363874
transform 1 0 852 0 1 275
box -3 -3 3 3
use NAND3X1  NAND3X1_76
timestamp 1680363874
transform 1 0 832 0 -1 370
box -8 -3 40 105
use FILL  FILL_10291
timestamp 1680363874
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_10293
timestamp 1680363874
transform 1 0 872 0 -1 370
box -8 -3 16 105
use FILL  FILL_10295
timestamp 1680363874
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_10297
timestamp 1680363874
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_10299
timestamp 1680363874
transform 1 0 896 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_656
timestamp 1680363874
transform 1 0 904 0 -1 370
box -9 -3 26 105
use FILL  FILL_10319
timestamp 1680363874
transform 1 0 920 0 -1 370
box -8 -3 16 105
use FILL  FILL_10320
timestamp 1680363874
transform 1 0 928 0 -1 370
box -8 -3 16 105
use FILL  FILL_10321
timestamp 1680363874
transform 1 0 936 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_377
timestamp 1680363874
transform -1 0 984 0 -1 370
box -8 -3 46 105
use FILL  FILL_10322
timestamp 1680363874
transform 1 0 984 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_569
timestamp 1680363874
transform 1 0 992 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_657
timestamp 1680363874
transform 1 0 1088 0 -1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_378
timestamp 1680363874
transform 1 0 1104 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_409
timestamp 1680363874
transform -1 0 1184 0 -1 370
box -8 -3 46 105
use FILL  FILL_10323
timestamp 1680363874
transform 1 0 1184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10324
timestamp 1680363874
transform 1 0 1192 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_658
timestamp 1680363874
transform 1 0 1200 0 -1 370
box -9 -3 26 105
use FILL  FILL_10325
timestamp 1680363874
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_10330
timestamp 1680363874
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_659
timestamp 1680363874
transform -1 0 1248 0 -1 370
box -9 -3 26 105
use FILL  FILL_10331
timestamp 1680363874
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_10332
timestamp 1680363874
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_10333
timestamp 1680363874
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_10334
timestamp 1680363874
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_10335
timestamp 1680363874
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_10336
timestamp 1680363874
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_410
timestamp 1680363874
transform -1 0 1336 0 -1 370
box -8 -3 46 105
use FILL  FILL_10337
timestamp 1680363874
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_10338
timestamp 1680363874
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_10351
timestamp 1680363874
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_10352
timestamp 1680363874
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_412
timestamp 1680363874
transform 1 0 1368 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_660
timestamp 1680363874
transform -1 0 1424 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_571
timestamp 1680363874
transform 1 0 1424 0 -1 370
box -8 -3 104 105
use FILL  FILL_10353
timestamp 1680363874
transform 1 0 1520 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_572
timestamp 1680363874
transform 1 0 1528 0 -1 370
box -8 -3 104 105
use FILL  FILL_10371
timestamp 1680363874
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_10372
timestamp 1680363874
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_415
timestamp 1680363874
transform -1 0 1680 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_573
timestamp 1680363874
transform 1 0 1680 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_662
timestamp 1680363874
transform 1 0 1776 0 -1 370
box -9 -3 26 105
use FILL  FILL_10373
timestamp 1680363874
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_10375
timestamp 1680363874
transform 1 0 1800 0 -1 370
box -8 -3 16 105
use FILL  FILL_10377
timestamp 1680363874
transform 1 0 1808 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_417
timestamp 1680363874
transform -1 0 1856 0 -1 370
box -8 -3 46 105
use FILL  FILL_10379
timestamp 1680363874
transform 1 0 1856 0 -1 370
box -8 -3 16 105
use FILL  FILL_10381
timestamp 1680363874
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_10386
timestamp 1680363874
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_663
timestamp 1680363874
transform 1 0 1880 0 -1 370
box -9 -3 26 105
use FILL  FILL_10387
timestamp 1680363874
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_381
timestamp 1680363874
transform -1 0 1944 0 -1 370
box -8 -3 46 105
use FILL  FILL_10388
timestamp 1680363874
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_10389
timestamp 1680363874
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_10390
timestamp 1680363874
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_10391
timestamp 1680363874
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_418
timestamp 1680363874
transform 1 0 1976 0 -1 370
box -8 -3 46 105
use FILL  FILL_10392
timestamp 1680363874
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_10394
timestamp 1680363874
transform 1 0 2024 0 -1 370
box -8 -3 16 105
use FILL  FILL_10395
timestamp 1680363874
transform 1 0 2032 0 -1 370
box -8 -3 16 105
use FILL  FILL_10396
timestamp 1680363874
transform 1 0 2040 0 -1 370
box -8 -3 16 105
use FILL  FILL_10397
timestamp 1680363874
transform 1 0 2048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10398
timestamp 1680363874
transform 1 0 2056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10399
timestamp 1680363874
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_10401
timestamp 1680363874
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10404
timestamp 1680363874
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_10405
timestamp 1680363874
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use FILL  FILL_10406
timestamp 1680363874
transform 1 0 2096 0 -1 370
box -8 -3 16 105
use FILL  FILL_10407
timestamp 1680363874
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_10409
timestamp 1680363874
transform 1 0 2112 0 -1 370
box -8 -3 16 105
use FILL  FILL_10412
timestamp 1680363874
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use FILL  FILL_10413
timestamp 1680363874
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_10414
timestamp 1680363874
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_10415
timestamp 1680363874
transform 1 0 2144 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_665
timestamp 1680363874
transform 1 0 2152 0 -1 370
box -9 -3 26 105
use FILL  FILL_10416
timestamp 1680363874
transform 1 0 2168 0 -1 370
box -8 -3 16 105
use FILL  FILL_10429
timestamp 1680363874
transform 1 0 2176 0 -1 370
box -8 -3 16 105
use FILL  FILL_10430
timestamp 1680363874
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_421
timestamp 1680363874
transform -1 0 2232 0 -1 370
box -8 -3 46 105
use FILL  FILL_10431
timestamp 1680363874
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_668
timestamp 1680363874
transform -1 0 2256 0 -1 370
box -9 -3 26 105
use FILL  FILL_10432
timestamp 1680363874
transform 1 0 2256 0 -1 370
box -8 -3 16 105
use FILL  FILL_10433
timestamp 1680363874
transform 1 0 2264 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_579
timestamp 1680363874
transform 1 0 2272 0 -1 370
box -8 -3 104 105
use FILL  FILL_10434
timestamp 1680363874
transform 1 0 2368 0 -1 370
box -8 -3 16 105
use FILL  FILL_10435
timestamp 1680363874
transform 1 0 2376 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_580
timestamp 1680363874
transform 1 0 2384 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_8652
timestamp 1680363874
transform 1 0 2492 0 1 275
box -3 -3 3 3
use INVX2  INVX2_669
timestamp 1680363874
transform -1 0 2496 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_116
timestamp 1680363874
transform -1 0 2520 0 -1 370
box -8 -3 32 105
use M3_M2  M3_M2_8653
timestamp 1680363874
transform 1 0 2572 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_581
timestamp 1680363874
transform 1 0 2520 0 -1 370
box -8 -3 104 105
use OAI22X1  OAI22X1_422
timestamp 1680363874
transform 1 0 2616 0 -1 370
box -8 -3 46 105
use FILL  FILL_10436
timestamp 1680363874
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_10437
timestamp 1680363874
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_10438
timestamp 1680363874
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_383
timestamp 1680363874
transform -1 0 2720 0 -1 370
box -8 -3 46 105
use FILL  FILL_10439
timestamp 1680363874
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_10441
timestamp 1680363874
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_10455
timestamp 1680363874
transform 1 0 2736 0 -1 370
box -8 -3 16 105
use FILL  FILL_10456
timestamp 1680363874
transform 1 0 2744 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_180
timestamp 1680363874
transform 1 0 2752 0 -1 370
box -8 -3 34 105
use FILL  FILL_10457
timestamp 1680363874
transform 1 0 2784 0 -1 370
box -8 -3 16 105
use FILL  FILL_10458
timestamp 1680363874
transform 1 0 2792 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_181
timestamp 1680363874
transform -1 0 2832 0 -1 370
box -8 -3 34 105
use FILL  FILL_10459
timestamp 1680363874
transform 1 0 2832 0 -1 370
box -8 -3 16 105
use FILL  FILL_10460
timestamp 1680363874
transform 1 0 2840 0 -1 370
box -8 -3 16 105
use FILL  FILL_10461
timestamp 1680363874
transform 1 0 2848 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_386
timestamp 1680363874
transform -1 0 2896 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_672
timestamp 1680363874
transform 1 0 2896 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_584
timestamp 1680363874
transform -1 0 3008 0 -1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_117
timestamp 1680363874
transform -1 0 3032 0 -1 370
box -8 -3 32 105
use FILL  FILL_10462
timestamp 1680363874
transform 1 0 3032 0 -1 370
box -8 -3 16 105
use FILL  FILL_10463
timestamp 1680363874
transform 1 0 3040 0 -1 370
box -8 -3 16 105
use FILL  FILL_10464
timestamp 1680363874
transform 1 0 3048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10465
timestamp 1680363874
transform 1 0 3056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10466
timestamp 1680363874
transform 1 0 3064 0 -1 370
box -8 -3 16 105
use FILL  FILL_10467
timestamp 1680363874
transform 1 0 3072 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_423
timestamp 1680363874
transform 1 0 3080 0 -1 370
box -8 -3 46 105
use FILL  FILL_10468
timestamp 1680363874
transform 1 0 3120 0 -1 370
box -8 -3 16 105
use FILL  FILL_10469
timestamp 1680363874
transform 1 0 3128 0 -1 370
box -8 -3 16 105
use FILL  FILL_10470
timestamp 1680363874
transform 1 0 3136 0 -1 370
box -8 -3 16 105
use FILL  FILL_10471
timestamp 1680363874
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_387
timestamp 1680363874
transform -1 0 3192 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_388
timestamp 1680363874
transform 1 0 3192 0 -1 370
box -8 -3 46 105
use FILL  FILL_10472
timestamp 1680363874
transform 1 0 3232 0 -1 370
box -8 -3 16 105
use FILL  FILL_10474
timestamp 1680363874
transform 1 0 3240 0 -1 370
box -8 -3 16 105
use FILL  FILL_10476
timestamp 1680363874
transform 1 0 3248 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_673
timestamp 1680363874
transform 1 0 3256 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_585
timestamp 1680363874
transform 1 0 3272 0 -1 370
box -8 -3 104 105
use FILL  FILL_10487
timestamp 1680363874
transform 1 0 3368 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_391
timestamp 1680363874
transform 1 0 3376 0 -1 370
box -8 -3 46 105
use FILL  FILL_10489
timestamp 1680363874
transform 1 0 3416 0 -1 370
box -8 -3 16 105
use FILL  FILL_10494
timestamp 1680363874
transform 1 0 3424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10495
timestamp 1680363874
transform 1 0 3432 0 -1 370
box -8 -3 16 105
use FILL  FILL_10496
timestamp 1680363874
transform 1 0 3440 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_676
timestamp 1680363874
transform 1 0 3448 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_588
timestamp 1680363874
transform -1 0 3560 0 -1 370
box -8 -3 104 105
use FILL  FILL_10497
timestamp 1680363874
transform 1 0 3560 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_392
timestamp 1680363874
transform -1 0 3608 0 -1 370
box -8 -3 46 105
use FILL  FILL_10498
timestamp 1680363874
transform 1 0 3608 0 -1 370
box -8 -3 16 105
use FILL  FILL_10499
timestamp 1680363874
transform 1 0 3616 0 -1 370
box -8 -3 16 105
use FILL  FILL_10500
timestamp 1680363874
transform 1 0 3624 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_393
timestamp 1680363874
transform 1 0 3632 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_394
timestamp 1680363874
transform -1 0 3712 0 -1 370
box -8 -3 46 105
use FILL  FILL_10501
timestamp 1680363874
transform 1 0 3712 0 -1 370
box -8 -3 16 105
use FILL  FILL_10503
timestamp 1680363874
transform 1 0 3720 0 -1 370
box -8 -3 16 105
use FILL  FILL_10510
timestamp 1680363874
transform 1 0 3728 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_678
timestamp 1680363874
transform 1 0 3736 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_425
timestamp 1680363874
transform 1 0 3752 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_8654
timestamp 1680363874
transform 1 0 3836 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_395
timestamp 1680363874
transform -1 0 3832 0 -1 370
box -8 -3 46 105
use FILL  FILL_10511
timestamp 1680363874
transform 1 0 3832 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_396
timestamp 1680363874
transform -1 0 3880 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_679
timestamp 1680363874
transform 1 0 3880 0 -1 370
box -9 -3 26 105
use FILL  FILL_10512
timestamp 1680363874
transform 1 0 3896 0 -1 370
box -8 -3 16 105
use FILL  FILL_10513
timestamp 1680363874
transform 1 0 3904 0 -1 370
box -8 -3 16 105
use FILL  FILL_10514
timestamp 1680363874
transform 1 0 3912 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8655
timestamp 1680363874
transform 1 0 3932 0 1 275
box -3 -3 3 3
use INVX2  INVX2_680
timestamp 1680363874
transform 1 0 3920 0 -1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_397
timestamp 1680363874
transform 1 0 3936 0 -1 370
box -8 -3 46 105
use FILL  FILL_10515
timestamp 1680363874
transform 1 0 3976 0 -1 370
box -8 -3 16 105
use FILL  FILL_10517
timestamp 1680363874
transform 1 0 3984 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_682
timestamp 1680363874
transform 1 0 3992 0 -1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_398
timestamp 1680363874
transform 1 0 4008 0 -1 370
box -8 -3 46 105
use FILL  FILL_10527
timestamp 1680363874
transform 1 0 4048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10528
timestamp 1680363874
transform 1 0 4056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10529
timestamp 1680363874
transform 1 0 4064 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8656
timestamp 1680363874
transform 1 0 4092 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_592
timestamp 1680363874
transform 1 0 4072 0 -1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_399
timestamp 1680363874
transform -1 0 4208 0 -1 370
box -8 -3 46 105
use FILL  FILL_10530
timestamp 1680363874
transform 1 0 4208 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_683
timestamp 1680363874
transform 1 0 4216 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_684
timestamp 1680363874
transform -1 0 4248 0 -1 370
box -9 -3 26 105
use FILL  FILL_10531
timestamp 1680363874
transform 1 0 4248 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_401
timestamp 1680363874
transform 1 0 4256 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_428
timestamp 1680363874
transform -1 0 4336 0 -1 370
box -8 -3 46 105
use FILL  FILL_10538
timestamp 1680363874
transform 1 0 4336 0 -1 370
box -8 -3 16 105
use FILL  FILL_10540
timestamp 1680363874
transform 1 0 4344 0 -1 370
box -8 -3 16 105
use FILL  FILL_10545
timestamp 1680363874
transform 1 0 4352 0 -1 370
box -8 -3 16 105
use FILL  FILL_10546
timestamp 1680363874
transform 1 0 4360 0 -1 370
box -8 -3 16 105
use FILL  FILL_10547
timestamp 1680363874
transform 1 0 4368 0 -1 370
box -8 -3 16 105
use FILL  FILL_10548
timestamp 1680363874
transform 1 0 4376 0 -1 370
box -8 -3 16 105
use FILL  FILL_10549
timestamp 1680363874
transform 1 0 4384 0 -1 370
box -8 -3 16 105
use FILL  FILL_10550
timestamp 1680363874
transform 1 0 4392 0 -1 370
box -8 -3 16 105
use FILL  FILL_10551
timestamp 1680363874
transform 1 0 4400 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_429
timestamp 1680363874
transform -1 0 4448 0 -1 370
box -8 -3 46 105
use FILL  FILL_10552
timestamp 1680363874
transform 1 0 4448 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_685
timestamp 1680363874
transform -1 0 4472 0 -1 370
box -9 -3 26 105
use FILL  FILL_10553
timestamp 1680363874
transform 1 0 4472 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_402
timestamp 1680363874
transform -1 0 4520 0 -1 370
box -8 -3 46 105
use FILL  FILL_10554
timestamp 1680363874
transform 1 0 4520 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_430
timestamp 1680363874
transform 1 0 4528 0 -1 370
box -8 -3 46 105
use FILL  FILL_10555
timestamp 1680363874
transform 1 0 4568 0 -1 370
box -8 -3 16 105
use FILL  FILL_10557
timestamp 1680363874
transform 1 0 4576 0 -1 370
box -8 -3 16 105
use FILL  FILL_10559
timestamp 1680363874
transform 1 0 4584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10562
timestamp 1680363874
transform 1 0 4592 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_403
timestamp 1680363874
transform 1 0 4600 0 -1 370
box -8 -3 46 105
use FILL  FILL_10563
timestamp 1680363874
transform 1 0 4640 0 -1 370
box -8 -3 16 105
use FILL  FILL_10565
timestamp 1680363874
transform 1 0 4648 0 -1 370
box -8 -3 16 105
use FILL  FILL_10567
timestamp 1680363874
transform 1 0 4656 0 -1 370
box -8 -3 16 105
use FILL  FILL_10569
timestamp 1680363874
transform 1 0 4664 0 -1 370
box -8 -3 16 105
use FILL  FILL_10571
timestamp 1680363874
transform 1 0 4672 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_686
timestamp 1680363874
transform 1 0 4680 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_596
timestamp 1680363874
transform 1 0 4696 0 -1 370
box -8 -3 104 105
use FILL  FILL_10575
timestamp 1680363874
transform 1 0 4792 0 -1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_89
timestamp 1680363874
transform 1 0 4851 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_8713
timestamp 1680363874
transform 1 0 220 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8714
timestamp 1680363874
transform 1 0 252 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8732
timestamp 1680363874
transform 1 0 172 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9681
timestamp 1680363874
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9820
timestamp 1680363874
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9682
timestamp 1680363874
transform 1 0 268 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8733
timestamp 1680363874
transform 1 0 324 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9683
timestamp 1680363874
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9684
timestamp 1680363874
transform 1 0 404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9821
timestamp 1680363874
transform 1 0 324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8779
timestamp 1680363874
transform 1 0 324 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9822
timestamp 1680363874
transform 1 0 412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8780
timestamp 1680363874
transform 1 0 412 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8685
timestamp 1680363874
transform 1 0 476 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9685
timestamp 1680363874
transform 1 0 476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9686
timestamp 1680363874
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9823
timestamp 1680363874
transform 1 0 492 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8781
timestamp 1680363874
transform 1 0 540 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8715
timestamp 1680363874
transform 1 0 596 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9687
timestamp 1680363874
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9824
timestamp 1680363874
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9688
timestamp 1680363874
transform 1 0 636 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8686
timestamp 1680363874
transform 1 0 652 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8716
timestamp 1680363874
transform 1 0 652 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9689
timestamp 1680363874
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9690
timestamp 1680363874
transform 1 0 668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9825
timestamp 1680363874
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9826
timestamp 1680363874
transform 1 0 660 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8820
timestamp 1680363874
transform 1 0 636 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8782
timestamp 1680363874
transform 1 0 660 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8821
timestamp 1680363874
transform 1 0 660 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8671
timestamp 1680363874
transform 1 0 684 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9827
timestamp 1680363874
transform 1 0 692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9828
timestamp 1680363874
transform 1 0 708 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8783
timestamp 1680363874
transform 1 0 700 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8687
timestamp 1680363874
transform 1 0 724 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8717
timestamp 1680363874
transform 1 0 748 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9691
timestamp 1680363874
transform 1 0 724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9692
timestamp 1680363874
transform 1 0 740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9829
timestamp 1680363874
transform 1 0 732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9830
timestamp 1680363874
transform 1 0 748 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8784
timestamp 1680363874
transform 1 0 748 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8688
timestamp 1680363874
transform 1 0 820 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9693
timestamp 1680363874
transform 1 0 788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9694
timestamp 1680363874
transform 1 0 804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9695
timestamp 1680363874
transform 1 0 820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9831
timestamp 1680363874
transform 1 0 788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9832
timestamp 1680363874
transform 1 0 812 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8822
timestamp 1680363874
transform 1 0 788 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8718
timestamp 1680363874
transform 1 0 836 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9833
timestamp 1680363874
transform 1 0 836 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8657
timestamp 1680363874
transform 1 0 972 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9696
timestamp 1680363874
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9697
timestamp 1680363874
transform 1 0 924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9834
timestamp 1680363874
transform 1 0 964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9835
timestamp 1680363874
transform 1 0 996 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8689
timestamp 1680363874
transform 1 0 1044 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9698
timestamp 1680363874
transform 1 0 1020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9699
timestamp 1680363874
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9836
timestamp 1680363874
transform 1 0 1028 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8785
timestamp 1680363874
transform 1 0 1020 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8786
timestamp 1680363874
transform 1 0 1044 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8734
timestamp 1680363874
transform 1 0 1060 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9837
timestamp 1680363874
transform 1 0 1060 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9700
timestamp 1680363874
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9701
timestamp 1680363874
transform 1 0 1156 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8735
timestamp 1680363874
transform 1 0 1180 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9838
timestamp 1680363874
transform 1 0 1180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8787
timestamp 1680363874
transform 1 0 1116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8788
timestamp 1680363874
transform 1 0 1180 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8823
timestamp 1680363874
transform 1 0 1204 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8690
timestamp 1680363874
transform 1 0 1228 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8736
timestamp 1680363874
transform 1 0 1236 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9702
timestamp 1680363874
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9703
timestamp 1680363874
transform 1 0 1308 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8737
timestamp 1680363874
transform 1 0 1332 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8691
timestamp 1680363874
transform 1 0 1372 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9704
timestamp 1680363874
transform 1 0 1356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9705
timestamp 1680363874
transform 1 0 1372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9839
timestamp 1680363874
transform 1 0 1332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9840
timestamp 1680363874
transform 1 0 1348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9841
timestamp 1680363874
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8789
timestamp 1680363874
transform 1 0 1260 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8790
timestamp 1680363874
transform 1 0 1332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8763
timestamp 1680363874
transform 1 0 1372 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8692
timestamp 1680363874
transform 1 0 1388 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9842
timestamp 1680363874
transform 1 0 1380 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8824
timestamp 1680363874
transform 1 0 1348 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8693
timestamp 1680363874
transform 1 0 1452 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9706
timestamp 1680363874
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9707
timestamp 1680363874
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9843
timestamp 1680363874
transform 1 0 1500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8791
timestamp 1680363874
transform 1 0 1516 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9844
timestamp 1680363874
transform 1 0 1524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8825
timestamp 1680363874
transform 1 0 1524 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9708
timestamp 1680363874
transform 1 0 1540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9709
timestamp 1680363874
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9845
timestamp 1680363874
transform 1 0 1548 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8764
timestamp 1680363874
transform 1 0 1556 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8792
timestamp 1680363874
transform 1 0 1556 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8826
timestamp 1680363874
transform 1 0 1572 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9846
timestamp 1680363874
transform 1 0 1588 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8827
timestamp 1680363874
transform 1 0 1588 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9710
timestamp 1680363874
transform 1 0 1604 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8738
timestamp 1680363874
transform 1 0 1612 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8694
timestamp 1680363874
transform 1 0 1628 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8739
timestamp 1680363874
transform 1 0 1636 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9711
timestamp 1680363874
transform 1 0 1644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9712
timestamp 1680363874
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8740
timestamp 1680363874
transform 1 0 1660 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9713
timestamp 1680363874
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8741
timestamp 1680363874
transform 1 0 1676 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9714
timestamp 1680363874
transform 1 0 1684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9847
timestamp 1680363874
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9848
timestamp 1680363874
transform 1 0 1628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9849
timestamp 1680363874
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8765
timestamp 1680363874
transform 1 0 1652 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9850
timestamp 1680363874
transform 1 0 1660 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8828
timestamp 1680363874
transform 1 0 1644 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8695
timestamp 1680363874
transform 1 0 1692 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9851
timestamp 1680363874
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8793
timestamp 1680363874
transform 1 0 1684 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8829
timestamp 1680363874
transform 1 0 1692 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8742
timestamp 1680363874
transform 1 0 1740 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8662
timestamp 1680363874
transform 1 0 1780 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9715
timestamp 1680363874
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9716
timestamp 1680363874
transform 1 0 1780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9852
timestamp 1680363874
transform 1 0 1740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9853
timestamp 1680363874
transform 1 0 1756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9854
timestamp 1680363874
transform 1 0 1772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9855
timestamp 1680363874
transform 1 0 1780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8830
timestamp 1680363874
transform 1 0 1772 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8663
timestamp 1680363874
transform 1 0 1812 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9717
timestamp 1680363874
transform 1 0 1836 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9718
timestamp 1680363874
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9856
timestamp 1680363874
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9857
timestamp 1680363874
transform 1 0 1892 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8794
timestamp 1680363874
transform 1 0 1804 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8831
timestamp 1680363874
transform 1 0 1788 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8832
timestamp 1680363874
transform 1 0 1868 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8795
timestamp 1680363874
transform 1 0 1900 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9719
timestamp 1680363874
transform 1 0 1916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9858
timestamp 1680363874
transform 1 0 1916 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8833
timestamp 1680363874
transform 1 0 1916 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9720
timestamp 1680363874
transform 1 0 1932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9721
timestamp 1680363874
transform 1 0 1948 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8696
timestamp 1680363874
transform 1 0 2116 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9722
timestamp 1680363874
transform 1 0 1996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9723
timestamp 1680363874
transform 1 0 2052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9724
timestamp 1680363874
transform 1 0 2116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9725
timestamp 1680363874
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9726
timestamp 1680363874
transform 1 0 2164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9727
timestamp 1680363874
transform 1 0 2180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9728
timestamp 1680363874
transform 1 0 2196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9859
timestamp 1680363874
transform 1 0 1940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9860
timestamp 1680363874
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9861
timestamp 1680363874
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8796
timestamp 1680363874
transform 1 0 1972 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9862
timestamp 1680363874
transform 1 0 2068 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8766
timestamp 1680363874
transform 1 0 2148 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9863
timestamp 1680363874
transform 1 0 2156 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8767
timestamp 1680363874
transform 1 0 2164 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9864
timestamp 1680363874
transform 1 0 2172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9865
timestamp 1680363874
transform 1 0 2188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9866
timestamp 1680363874
transform 1 0 2196 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8834
timestamp 1680363874
transform 1 0 2188 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8697
timestamp 1680363874
transform 1 0 2212 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9729
timestamp 1680363874
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9730
timestamp 1680363874
transform 1 0 2220 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8768
timestamp 1680363874
transform 1 0 2212 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8797
timestamp 1680363874
transform 1 0 2212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8743
timestamp 1680363874
transform 1 0 2236 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9731
timestamp 1680363874
transform 1 0 2260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9732
timestamp 1680363874
transform 1 0 2276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9867
timestamp 1680363874
transform 1 0 2228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9868
timestamp 1680363874
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9869
timestamp 1680363874
transform 1 0 2252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9870
timestamp 1680363874
transform 1 0 2268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9871
timestamp 1680363874
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8835
timestamp 1680363874
transform 1 0 2228 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8798
timestamp 1680363874
transform 1 0 2276 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8836
timestamp 1680363874
transform 1 0 2268 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9733
timestamp 1680363874
transform 1 0 2356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9872
timestamp 1680363874
transform 1 0 2308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8799
timestamp 1680363874
transform 1 0 2356 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9734
timestamp 1680363874
transform 1 0 2420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9735
timestamp 1680363874
transform 1 0 2436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9736
timestamp 1680363874
transform 1 0 2452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9873
timestamp 1680363874
transform 1 0 2428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9874
timestamp 1680363874
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8769
timestamp 1680363874
transform 1 0 2452 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8800
timestamp 1680363874
transform 1 0 2444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8837
timestamp 1680363874
transform 1 0 2428 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8838
timestamp 1680363874
transform 1 0 2460 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9875
timestamp 1680363874
transform 1 0 2476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9876
timestamp 1680363874
transform 1 0 2484 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8664
timestamp 1680363874
transform 1 0 2500 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9737
timestamp 1680363874
transform 1 0 2500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9877
timestamp 1680363874
transform 1 0 2516 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8698
timestamp 1680363874
transform 1 0 2540 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9676
timestamp 1680363874
transform 1 0 2540 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9738
timestamp 1680363874
transform 1 0 2556 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8672
timestamp 1680363874
transform 1 0 2572 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9878
timestamp 1680363874
transform 1 0 2564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9879
timestamp 1680363874
transform 1 0 2572 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8673
timestamp 1680363874
transform 1 0 2596 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9739
timestamp 1680363874
transform 1 0 2596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9740
timestamp 1680363874
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8744
timestamp 1680363874
transform 1 0 2620 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9741
timestamp 1680363874
transform 1 0 2628 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8770
timestamp 1680363874
transform 1 0 2612 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9880
timestamp 1680363874
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9881
timestamp 1680363874
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9882
timestamp 1680363874
transform 1 0 2644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8801
timestamp 1680363874
transform 1 0 2628 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8839
timestamp 1680363874
transform 1 0 2636 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9742
timestamp 1680363874
transform 1 0 2660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9743
timestamp 1680363874
transform 1 0 2676 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8771
timestamp 1680363874
transform 1 0 2660 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9744
timestamp 1680363874
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9883
timestamp 1680363874
transform 1 0 2668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9884
timestamp 1680363874
transform 1 0 2684 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8840
timestamp 1680363874
transform 1 0 2684 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8745
timestamp 1680363874
transform 1 0 2700 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9885
timestamp 1680363874
transform 1 0 2700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9886
timestamp 1680363874
transform 1 0 2724 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8802
timestamp 1680363874
transform 1 0 2724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8674
timestamp 1680363874
transform 1 0 2740 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8658
timestamp 1680363874
transform 1 0 2804 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8675
timestamp 1680363874
transform 1 0 2764 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8676
timestamp 1680363874
transform 1 0 2780 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8677
timestamp 1680363874
transform 1 0 2796 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8699
timestamp 1680363874
transform 1 0 2764 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8700
timestamp 1680363874
transform 1 0 2780 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8719
timestamp 1680363874
transform 1 0 2756 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9677
timestamp 1680363874
transform 1 0 2764 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9745
timestamp 1680363874
transform 1 0 2732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9746
timestamp 1680363874
transform 1 0 2740 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8746
timestamp 1680363874
transform 1 0 2764 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8701
timestamp 1680363874
transform 1 0 2804 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9678
timestamp 1680363874
transform 1 0 2796 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9747
timestamp 1680363874
transform 1 0 2772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9887
timestamp 1680363874
transform 1 0 2764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9888
timestamp 1680363874
transform 1 0 2772 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8803
timestamp 1680363874
transform 1 0 2756 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9748
timestamp 1680363874
transform 1 0 2812 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8665
timestamp 1680363874
transform 1 0 2852 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9679
timestamp 1680363874
transform 1 0 2836 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8720
timestamp 1680363874
transform 1 0 2860 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8747
timestamp 1680363874
transform 1 0 2836 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9749
timestamp 1680363874
transform 1 0 2852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9750
timestamp 1680363874
transform 1 0 2860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9751
timestamp 1680363874
transform 1 0 2884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9889
timestamp 1680363874
transform 1 0 2804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9890
timestamp 1680363874
transform 1 0 2812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9891
timestamp 1680363874
transform 1 0 2828 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8804
timestamp 1680363874
transform 1 0 2812 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9949
timestamp 1680363874
transform 1 0 2828 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_8841
timestamp 1680363874
transform 1 0 2828 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8748
timestamp 1680363874
transform 1 0 2892 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8721
timestamp 1680363874
transform 1 0 2908 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9752
timestamp 1680363874
transform 1 0 2900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9753
timestamp 1680363874
transform 1 0 2908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9892
timestamp 1680363874
transform 1 0 2860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9893
timestamp 1680363874
transform 1 0 2892 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8772
timestamp 1680363874
transform 1 0 2900 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8666
timestamp 1680363874
transform 1 0 2972 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8678
timestamp 1680363874
transform 1 0 2964 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9754
timestamp 1680363874
transform 1 0 2948 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8749
timestamp 1680363874
transform 1 0 2956 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9755
timestamp 1680363874
transform 1 0 2964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9756
timestamp 1680363874
transform 1 0 2972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9894
timestamp 1680363874
transform 1 0 2940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9895
timestamp 1680363874
transform 1 0 2956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9896
timestamp 1680363874
transform 1 0 2964 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8805
timestamp 1680363874
transform 1 0 2940 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8806
timestamp 1680363874
transform 1 0 2964 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8702
timestamp 1680363874
transform 1 0 3004 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9680
timestamp 1680363874
transform 1 0 3004 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9897
timestamp 1680363874
transform 1 0 3012 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8722
timestamp 1680363874
transform 1 0 3108 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8723
timestamp 1680363874
transform 1 0 3148 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9757
timestamp 1680363874
transform 1 0 3108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9758
timestamp 1680363874
transform 1 0 3140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9759
timestamp 1680363874
transform 1 0 3148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9760
timestamp 1680363874
transform 1 0 3156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9898
timestamp 1680363874
transform 1 0 3060 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8807
timestamp 1680363874
transform 1 0 3076 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8773
timestamp 1680363874
transform 1 0 3156 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8703
timestamp 1680363874
transform 1 0 3188 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8679
timestamp 1680363874
transform 1 0 3260 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9761
timestamp 1680363874
transform 1 0 3188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9762
timestamp 1680363874
transform 1 0 3204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9763
timestamp 1680363874
transform 1 0 3228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9899
timestamp 1680363874
transform 1 0 3172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9900
timestamp 1680363874
transform 1 0 3180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8750
timestamp 1680363874
transform 1 0 3236 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9764
timestamp 1680363874
transform 1 0 3244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9765
timestamp 1680363874
transform 1 0 3260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9766
timestamp 1680363874
transform 1 0 3276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9767
timestamp 1680363874
transform 1 0 3292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9901
timestamp 1680363874
transform 1 0 3196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9902
timestamp 1680363874
transform 1 0 3220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9903
timestamp 1680363874
transform 1 0 3236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9904
timestamp 1680363874
transform 1 0 3252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9905
timestamp 1680363874
transform 1 0 3260 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8808
timestamp 1680363874
transform 1 0 3196 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8809
timestamp 1680363874
transform 1 0 3252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8774
timestamp 1680363874
transform 1 0 3276 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9906
timestamp 1680363874
transform 1 0 3284 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8751
timestamp 1680363874
transform 1 0 3316 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8667
timestamp 1680363874
transform 1 0 3348 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9768
timestamp 1680363874
transform 1 0 3324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9769
timestamp 1680363874
transform 1 0 3340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9907
timestamp 1680363874
transform 1 0 3308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9908
timestamp 1680363874
transform 1 0 3316 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8810
timestamp 1680363874
transform 1 0 3308 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8842
timestamp 1680363874
transform 1 0 3284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8775
timestamp 1680363874
transform 1 0 3324 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8724
timestamp 1680363874
transform 1 0 3364 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8704
timestamp 1680363874
transform 1 0 3396 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9770
timestamp 1680363874
transform 1 0 3364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9771
timestamp 1680363874
transform 1 0 3380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9909
timestamp 1680363874
transform 1 0 3332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9910
timestamp 1680363874
transform 1 0 3348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9911
timestamp 1680363874
transform 1 0 3356 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8811
timestamp 1680363874
transform 1 0 3356 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8843
timestamp 1680363874
transform 1 0 3348 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8752
timestamp 1680363874
transform 1 0 3388 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9772
timestamp 1680363874
transform 1 0 3396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9912
timestamp 1680363874
transform 1 0 3372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9913
timestamp 1680363874
transform 1 0 3388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9914
timestamp 1680363874
transform 1 0 3396 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8776
timestamp 1680363874
transform 1 0 3404 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8725
timestamp 1680363874
transform 1 0 3420 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8680
timestamp 1680363874
transform 1 0 3452 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8726
timestamp 1680363874
transform 1 0 3452 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9773
timestamp 1680363874
transform 1 0 3412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9774
timestamp 1680363874
transform 1 0 3420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9775
timestamp 1680363874
transform 1 0 3436 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8753
timestamp 1680363874
transform 1 0 3444 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9776
timestamp 1680363874
transform 1 0 3452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9915
timestamp 1680363874
transform 1 0 3420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9916
timestamp 1680363874
transform 1 0 3444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9917
timestamp 1680363874
transform 1 0 3452 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8844
timestamp 1680363874
transform 1 0 3420 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8845
timestamp 1680363874
transform 1 0 3476 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8681
timestamp 1680363874
transform 1 0 3500 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8682
timestamp 1680363874
transform 1 0 3564 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8705
timestamp 1680363874
transform 1 0 3556 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8706
timestamp 1680363874
transform 1 0 3596 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9777
timestamp 1680363874
transform 1 0 3492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9778
timestamp 1680363874
transform 1 0 3500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9779
timestamp 1680363874
transform 1 0 3556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9780
timestamp 1680363874
transform 1 0 3596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9918
timestamp 1680363874
transform 1 0 3580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9919
timestamp 1680363874
transform 1 0 3596 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8812
timestamp 1680363874
transform 1 0 3580 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8813
timestamp 1680363874
transform 1 0 3620 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9781
timestamp 1680363874
transform 1 0 3644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9920
timestamp 1680363874
transform 1 0 3636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9782
timestamp 1680363874
transform 1 0 3676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9783
timestamp 1680363874
transform 1 0 3732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9921
timestamp 1680363874
transform 1 0 3756 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8814
timestamp 1680363874
transform 1 0 3756 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8754
timestamp 1680363874
transform 1 0 3788 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9922
timestamp 1680363874
transform 1 0 3788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9784
timestamp 1680363874
transform 1 0 3804 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8755
timestamp 1680363874
transform 1 0 3812 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9785
timestamp 1680363874
transform 1 0 3828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9786
timestamp 1680363874
transform 1 0 3884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9923
timestamp 1680363874
transform 1 0 3908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9787
timestamp 1680363874
transform 1 0 3932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9924
timestamp 1680363874
transform 1 0 3956 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8659
timestamp 1680363874
transform 1 0 3972 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8668
timestamp 1680363874
transform 1 0 4084 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8660
timestamp 1680363874
transform 1 0 4116 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9788
timestamp 1680363874
transform 1 0 4004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9789
timestamp 1680363874
transform 1 0 4060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9790
timestamp 1680363874
transform 1 0 4068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9791
timestamp 1680363874
transform 1 0 4084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9925
timestamp 1680363874
transform 1 0 3980 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8815
timestamp 1680363874
transform 1 0 3980 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8756
timestamp 1680363874
transform 1 0 4092 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9792
timestamp 1680363874
transform 1 0 4100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9793
timestamp 1680363874
transform 1 0 4116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9926
timestamp 1680363874
transform 1 0 4084 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9927
timestamp 1680363874
transform 1 0 4092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9928
timestamp 1680363874
transform 1 0 4108 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8816
timestamp 1680363874
transform 1 0 4076 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9929
timestamp 1680363874
transform 1 0 4132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9794
timestamp 1680363874
transform 1 0 4156 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8757
timestamp 1680363874
transform 1 0 4164 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8669
timestamp 1680363874
transform 1 0 4252 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9795
timestamp 1680363874
transform 1 0 4180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9796
timestamp 1680363874
transform 1 0 4188 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8758
timestamp 1680363874
transform 1 0 4204 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8727
timestamp 1680363874
transform 1 0 4292 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9797
timestamp 1680363874
transform 1 0 4236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9798
timestamp 1680363874
transform 1 0 4284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9930
timestamp 1680363874
transform 1 0 4148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9931
timestamp 1680363874
transform 1 0 4164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9932
timestamp 1680363874
transform 1 0 4172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9933
timestamp 1680363874
transform 1 0 4204 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8817
timestamp 1680363874
transform 1 0 4204 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9799
timestamp 1680363874
transform 1 0 4300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9934
timestamp 1680363874
transform 1 0 4292 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8661
timestamp 1680363874
transform 1 0 4340 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8707
timestamp 1680363874
transform 1 0 4340 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9800
timestamp 1680363874
transform 1 0 4324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9801
timestamp 1680363874
transform 1 0 4340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9935
timestamp 1680363874
transform 1 0 4332 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8818
timestamp 1680363874
transform 1 0 4316 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8819
timestamp 1680363874
transform 1 0 4332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8670
timestamp 1680363874
transform 1 0 4372 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8708
timestamp 1680363874
transform 1 0 4452 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8728
timestamp 1680363874
transform 1 0 4412 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8729
timestamp 1680363874
transform 1 0 4444 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8759
timestamp 1680363874
transform 1 0 4364 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8683
timestamp 1680363874
transform 1 0 4484 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9802
timestamp 1680363874
transform 1 0 4412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9803
timestamp 1680363874
transform 1 0 4444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9804
timestamp 1680363874
transform 1 0 4452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9805
timestamp 1680363874
transform 1 0 4468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9936
timestamp 1680363874
transform 1 0 4364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8760
timestamp 1680363874
transform 1 0 4476 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9806
timestamp 1680363874
transform 1 0 4484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9937
timestamp 1680363874
transform 1 0 4460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9938
timestamp 1680363874
transform 1 0 4476 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8709
timestamp 1680363874
transform 1 0 4500 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9807
timestamp 1680363874
transform 1 0 4500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9939
timestamp 1680363874
transform 1 0 4500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8684
timestamp 1680363874
transform 1 0 4516 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9808
timestamp 1680363874
transform 1 0 4524 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8761
timestamp 1680363874
transform 1 0 4532 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9809
timestamp 1680363874
transform 1 0 4540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9810
timestamp 1680363874
transform 1 0 4556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9940
timestamp 1680363874
transform 1 0 4516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9941
timestamp 1680363874
transform 1 0 4532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9942
timestamp 1680363874
transform 1 0 4540 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8710
timestamp 1680363874
transform 1 0 4580 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9811
timestamp 1680363874
transform 1 0 4580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9943
timestamp 1680363874
transform 1 0 4588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9812
timestamp 1680363874
transform 1 0 4612 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8762
timestamp 1680363874
transform 1 0 4620 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8711
timestamp 1680363874
transform 1 0 4644 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9813
timestamp 1680363874
transform 1 0 4628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9814
timestamp 1680363874
transform 1 0 4636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9815
timestamp 1680363874
transform 1 0 4652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9944
timestamp 1680363874
transform 1 0 4620 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8777
timestamp 1680363874
transform 1 0 4628 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9816
timestamp 1680363874
transform 1 0 4676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9945
timestamp 1680363874
transform 1 0 4644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9946
timestamp 1680363874
transform 1 0 4660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9947
timestamp 1680363874
transform 1 0 4668 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8778
timestamp 1680363874
transform 1 0 4676 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8712
timestamp 1680363874
transform 1 0 4796 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8730
timestamp 1680363874
transform 1 0 4700 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8731
timestamp 1680363874
transform 1 0 4740 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9817
timestamp 1680363874
transform 1 0 4700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9818
timestamp 1680363874
transform 1 0 4740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9819
timestamp 1680363874
transform 1 0 4796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9948
timestamp 1680363874
transform 1 0 4716 0 1 205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_90
timestamp 1680363874
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_10576
timestamp 1680363874
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_10578
timestamp 1680363874
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_10580
timestamp 1680363874
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_10582
timestamp 1680363874
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_10584
timestamp 1680363874
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_10586
timestamp 1680363874
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_10588
timestamp 1680363874
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_10590
timestamp 1680363874
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_10592
timestamp 1680363874
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_10594
timestamp 1680363874
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_10596
timestamp 1680363874
transform 1 0 152 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_597
timestamp 1680363874
transform 1 0 160 0 1 170
box -8 -3 104 105
use INVX2  INVX2_687
timestamp 1680363874
transform 1 0 256 0 1 170
box -9 -3 26 105
use FILL  FILL_10598
timestamp 1680363874
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_10614
timestamp 1680363874
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_10616
timestamp 1680363874
transform 1 0 288 0 1 170
box -8 -3 16 105
use FILL  FILL_10618
timestamp 1680363874
transform 1 0 296 0 1 170
box -8 -3 16 105
use FILL  FILL_10620
timestamp 1680363874
transform 1 0 304 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_598
timestamp 1680363874
transform 1 0 312 0 1 170
box -8 -3 104 105
use FILL  FILL_10622
timestamp 1680363874
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_10623
timestamp 1680363874
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_10626
timestamp 1680363874
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_10627
timestamp 1680363874
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_10628
timestamp 1680363874
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_10629
timestamp 1680363874
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_10630
timestamp 1680363874
transform 1 0 456 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8846
timestamp 1680363874
transform 1 0 492 0 1 175
box -3 -3 3 3
use INVX2  INVX2_688
timestamp 1680363874
transform 1 0 464 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_600
timestamp 1680363874
transform 1 0 480 0 1 170
box -8 -3 104 105
use INVX2  INVX2_689
timestamp 1680363874
transform 1 0 576 0 1 170
box -9 -3 26 105
use INVX2  INVX2_690
timestamp 1680363874
transform 1 0 592 0 1 170
box -9 -3 26 105
use FILL  FILL_10631
timestamp 1680363874
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_10632
timestamp 1680363874
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_10633
timestamp 1680363874
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_10634
timestamp 1680363874
transform 1 0 632 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_432
timestamp 1680363874
transform -1 0 680 0 1 170
box -8 -3 46 105
use FILL  FILL_10635
timestamp 1680363874
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_10636
timestamp 1680363874
transform 1 0 688 0 1 170
box -8 -3 16 105
use FILL  FILL_10642
timestamp 1680363874
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_10644
timestamp 1680363874
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_10645
timestamp 1680363874
transform 1 0 712 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_404
timestamp 1680363874
transform 1 0 720 0 1 170
box -8 -3 46 105
use FILL  FILL_10646
timestamp 1680363874
transform 1 0 760 0 1 170
box -8 -3 16 105
use FILL  FILL_10648
timestamp 1680363874
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_10650
timestamp 1680363874
transform 1 0 776 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_405
timestamp 1680363874
transform -1 0 824 0 1 170
box -8 -3 46 105
use FILL  FILL_10651
timestamp 1680363874
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_10652
timestamp 1680363874
transform 1 0 832 0 1 170
box -8 -3 16 105
use INVX2  INVX2_692
timestamp 1680363874
transform 1 0 840 0 1 170
box -9 -3 26 105
use FILL  FILL_10653
timestamp 1680363874
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_10654
timestamp 1680363874
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_10655
timestamp 1680363874
transform 1 0 872 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8847
timestamp 1680363874
transform 1 0 964 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_603
timestamp 1680363874
transform -1 0 976 0 1 170
box -8 -3 104 105
use FILL  FILL_10656
timestamp 1680363874
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_10657
timestamp 1680363874
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_10658
timestamp 1680363874
transform 1 0 992 0 1 170
box -8 -3 16 105
use FILL  FILL_10659
timestamp 1680363874
transform 1 0 1000 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_435
timestamp 1680363874
transform -1 0 1048 0 1 170
box -8 -3 46 105
use FILL  FILL_10660
timestamp 1680363874
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_10665
timestamp 1680363874
transform 1 0 1056 0 1 170
box -8 -3 16 105
use FILL  FILL_10667
timestamp 1680363874
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_10669
timestamp 1680363874
transform 1 0 1072 0 1 170
box -8 -3 16 105
use FILL  FILL_10670
timestamp 1680363874
transform 1 0 1080 0 1 170
box -8 -3 16 105
use FILL  FILL_10671
timestamp 1680363874
transform 1 0 1088 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_606
timestamp 1680363874
transform -1 0 1192 0 1 170
box -8 -3 104 105
use FILL  FILL_10672
timestamp 1680363874
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_10673
timestamp 1680363874
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_10674
timestamp 1680363874
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_10675
timestamp 1680363874
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_10676
timestamp 1680363874
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_10677
timestamp 1680363874
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_10678
timestamp 1680363874
transform 1 0 1240 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_607
timestamp 1680363874
transform -1 0 1344 0 1 170
box -8 -3 104 105
use OAI22X1  OAI22X1_437
timestamp 1680363874
transform -1 0 1384 0 1 170
box -8 -3 46 105
use FILL  FILL_10679
timestamp 1680363874
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_10687
timestamp 1680363874
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_10689
timestamp 1680363874
transform 1 0 1400 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8848
timestamp 1680363874
transform 1 0 1500 0 1 175
box -3 -3 3 3
use FILL  FILL_10691
timestamp 1680363874
transform 1 0 1408 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_610
timestamp 1680363874
transform -1 0 1512 0 1 170
box -8 -3 104 105
use FILL  FILL_10692
timestamp 1680363874
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_10693
timestamp 1680363874
transform 1 0 1520 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_439
timestamp 1680363874
transform -1 0 1568 0 1 170
box -8 -3 46 105
use FILL  FILL_10694
timestamp 1680363874
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_10695
timestamp 1680363874
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_10696
timestamp 1680363874
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_10697
timestamp 1680363874
transform 1 0 1592 0 1 170
box -8 -3 16 105
use INVX2  INVX2_696
timestamp 1680363874
transform -1 0 1616 0 1 170
box -9 -3 26 105
use FILL  FILL_10698
timestamp 1680363874
transform 1 0 1616 0 1 170
box -8 -3 16 105
use INVX2  INVX2_697
timestamp 1680363874
transform 1 0 1624 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_440
timestamp 1680363874
transform 1 0 1640 0 1 170
box -8 -3 46 105
use FILL  FILL_10699
timestamp 1680363874
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_10700
timestamp 1680363874
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_10701
timestamp 1680363874
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_10702
timestamp 1680363874
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_10703
timestamp 1680363874
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_10704
timestamp 1680363874
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_10705
timestamp 1680363874
transform 1 0 1728 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_441
timestamp 1680363874
transform 1 0 1736 0 1 170
box -8 -3 46 105
use INVX2  INVX2_698
timestamp 1680363874
transform 1 0 1776 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_611
timestamp 1680363874
transform 1 0 1792 0 1 170
box -8 -3 104 105
use INVX2  INVX2_699
timestamp 1680363874
transform 1 0 1888 0 1 170
box -9 -3 26 105
use FILL  FILL_10706
timestamp 1680363874
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_10707
timestamp 1680363874
transform 1 0 1912 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8849
timestamp 1680363874
transform 1 0 1948 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_442
timestamp 1680363874
transform -1 0 1960 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_8850
timestamp 1680363874
transform 1 0 2004 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_612
timestamp 1680363874
transform 1 0 1960 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_613
timestamp 1680363874
transform 1 0 2056 0 1 170
box -8 -3 104 105
use OAI22X1  OAI22X1_443
timestamp 1680363874
transform 1 0 2152 0 1 170
box -8 -3 46 105
use INVX2  INVX2_700
timestamp 1680363874
transform 1 0 2192 0 1 170
box -9 -3 26 105
use FILL  FILL_10708
timestamp 1680363874
transform 1 0 2208 0 1 170
box -8 -3 16 105
use INVX2  INVX2_701
timestamp 1680363874
transform -1 0 2232 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_444
timestamp 1680363874
transform 1 0 2232 0 1 170
box -8 -3 46 105
use FILL  FILL_10709
timestamp 1680363874
transform 1 0 2272 0 1 170
box -8 -3 16 105
use INVX2  INVX2_702
timestamp 1680363874
transform 1 0 2280 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_614
timestamp 1680363874
transform 1 0 2296 0 1 170
box -8 -3 104 105
use INVX2  INVX2_703
timestamp 1680363874
transform 1 0 2392 0 1 170
box -9 -3 26 105
use FILL  FILL_10710
timestamp 1680363874
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_10711
timestamp 1680363874
transform 1 0 2416 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_445
timestamp 1680363874
transform -1 0 2464 0 1 170
box -8 -3 46 105
use FILL  FILL_10712
timestamp 1680363874
transform 1 0 2464 0 1 170
box -8 -3 16 105
use FILL  FILL_10736
timestamp 1680363874
transform 1 0 2472 0 1 170
box -8 -3 16 105
use FILL  FILL_10737
timestamp 1680363874
transform 1 0 2480 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8851
timestamp 1680363874
transform 1 0 2516 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_182
timestamp 1680363874
transform 1 0 2488 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_8852
timestamp 1680363874
transform 1 0 2532 0 1 175
box -3 -3 3 3
use FILL  FILL_10738
timestamp 1680363874
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_10739
timestamp 1680363874
transform 1 0 2528 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_183
timestamp 1680363874
transform -1 0 2568 0 1 170
box -8 -3 34 105
use FILL  FILL_10740
timestamp 1680363874
transform 1 0 2568 0 1 170
box -8 -3 16 105
use FILL  FILL_10741
timestamp 1680363874
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_10742
timestamp 1680363874
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_10743
timestamp 1680363874
transform 1 0 2592 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_448
timestamp 1680363874
transform 1 0 2600 0 1 170
box -8 -3 46 105
use FILL  FILL_10744
timestamp 1680363874
transform 1 0 2640 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_449
timestamp 1680363874
transform 1 0 2648 0 1 170
box -8 -3 46 105
use FILL  FILL_10751
timestamp 1680363874
transform 1 0 2688 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8853
timestamp 1680363874
transform 1 0 2708 0 1 175
box -3 -3 3 3
use FILL  FILL_10752
timestamp 1680363874
transform 1 0 2696 0 1 170
box -8 -3 16 105
use INVX2  INVX2_708
timestamp 1680363874
transform 1 0 2704 0 1 170
box -9 -3 26 105
use FILL  FILL_10753
timestamp 1680363874
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_10754
timestamp 1680363874
transform 1 0 2728 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_184
timestamp 1680363874
transform 1 0 2736 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1680363874
transform 1 0 2768 0 1 170
box -8 -3 34 105
use FILL  FILL_10755
timestamp 1680363874
transform 1 0 2800 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_118
timestamp 1680363874
transform -1 0 2832 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_186
timestamp 1680363874
transform -1 0 2864 0 1 170
box -8 -3 34 105
use AOI22X1  AOI22X1_406
timestamp 1680363874
transform -1 0 2904 0 1 170
box -8 -3 46 105
use FILL  FILL_10756
timestamp 1680363874
transform 1 0 2904 0 1 170
box -8 -3 16 105
use FILL  FILL_10757
timestamp 1680363874
transform 1 0 2912 0 1 170
box -8 -3 16 105
use FILL  FILL_10758
timestamp 1680363874
transform 1 0 2920 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_407
timestamp 1680363874
transform -1 0 2968 0 1 170
box -8 -3 46 105
use FILL  FILL_10759
timestamp 1680363874
transform 1 0 2968 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_187
timestamp 1680363874
transform 1 0 2976 0 1 170
box -8 -3 34 105
use FILL  FILL_10760
timestamp 1680363874
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_10761
timestamp 1680363874
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_10762
timestamp 1680363874
transform 1 0 3024 0 1 170
box -8 -3 16 105
use FILL  FILL_10763
timestamp 1680363874
transform 1 0 3032 0 1 170
box -8 -3 16 105
use FILL  FILL_10764
timestamp 1680363874
transform 1 0 3040 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8854
timestamp 1680363874
transform 1 0 3060 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_8855
timestamp 1680363874
transform 1 0 3124 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_624
timestamp 1680363874
transform 1 0 3048 0 1 170
box -8 -3 104 105
use INVX2  INVX2_709
timestamp 1680363874
transform -1 0 3160 0 1 170
box -9 -3 26 105
use FILL  FILL_10765
timestamp 1680363874
transform 1 0 3160 0 1 170
box -8 -3 16 105
use FILL  FILL_10766
timestamp 1680363874
transform 1 0 3168 0 1 170
box -8 -3 16 105
use FILL  FILL_10767
timestamp 1680363874
transform 1 0 3176 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8856
timestamp 1680363874
transform 1 0 3204 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_8857
timestamp 1680363874
transform 1 0 3220 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_408
timestamp 1680363874
transform 1 0 3184 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_8858
timestamp 1680363874
transform 1 0 3260 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_409
timestamp 1680363874
transform -1 0 3264 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_450
timestamp 1680363874
transform -1 0 3304 0 1 170
box -8 -3 46 105
use FILL  FILL_10768
timestamp 1680363874
transform 1 0 3304 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_451
timestamp 1680363874
transform -1 0 3352 0 1 170
box -8 -3 46 105
use FILL  FILL_10769
timestamp 1680363874
transform 1 0 3352 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_410
timestamp 1680363874
transform -1 0 3400 0 1 170
box -8 -3 46 105
use INVX2  INVX2_710
timestamp 1680363874
transform 1 0 3400 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_411
timestamp 1680363874
transform -1 0 3456 0 1 170
box -8 -3 46 105
use FILL  FILL_10770
timestamp 1680363874
transform 1 0 3456 0 1 170
box -8 -3 16 105
use FILL  FILL_10771
timestamp 1680363874
transform 1 0 3464 0 1 170
box -8 -3 16 105
use FILL  FILL_10772
timestamp 1680363874
transform 1 0 3472 0 1 170
box -8 -3 16 105
use INVX2  INVX2_716
timestamp 1680363874
transform 1 0 3480 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_631
timestamp 1680363874
transform -1 0 3592 0 1 170
box -8 -3 104 105
use INVX2  INVX2_717
timestamp 1680363874
transform 1 0 3592 0 1 170
box -9 -3 26 105
use FILL  FILL_10790
timestamp 1680363874
transform 1 0 3608 0 1 170
box -8 -3 16 105
use FILL  FILL_10791
timestamp 1680363874
transform 1 0 3616 0 1 170
box -8 -3 16 105
use FILL  FILL_10792
timestamp 1680363874
transform 1 0 3624 0 1 170
box -8 -3 16 105
use INVX2  INVX2_718
timestamp 1680363874
transform 1 0 3632 0 1 170
box -9 -3 26 105
use FILL  FILL_10793
timestamp 1680363874
transform 1 0 3648 0 1 170
box -8 -3 16 105
use FILL  FILL_10794
timestamp 1680363874
transform 1 0 3656 0 1 170
box -8 -3 16 105
use FILL  FILL_10795
timestamp 1680363874
transform 1 0 3664 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_632
timestamp 1680363874
transform -1 0 3768 0 1 170
box -8 -3 104 105
use FILL  FILL_10796
timestamp 1680363874
transform 1 0 3768 0 1 170
box -8 -3 16 105
use FILL  FILL_10797
timestamp 1680363874
transform 1 0 3776 0 1 170
box -8 -3 16 105
use INVX2  INVX2_719
timestamp 1680363874
transform 1 0 3784 0 1 170
box -9 -3 26 105
use FILL  FILL_10798
timestamp 1680363874
transform 1 0 3800 0 1 170
box -8 -3 16 105
use FILL  FILL_10799
timestamp 1680363874
transform 1 0 3808 0 1 170
box -8 -3 16 105
use FILL  FILL_10800
timestamp 1680363874
transform 1 0 3816 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_633
timestamp 1680363874
transform -1 0 3920 0 1 170
box -8 -3 104 105
use FILL  FILL_10801
timestamp 1680363874
transform 1 0 3920 0 1 170
box -8 -3 16 105
use FILL  FILL_10802
timestamp 1680363874
transform 1 0 3928 0 1 170
box -8 -3 16 105
use FILL  FILL_10803
timestamp 1680363874
transform 1 0 3936 0 1 170
box -8 -3 16 105
use INVX2  INVX2_720
timestamp 1680363874
transform -1 0 3960 0 1 170
box -9 -3 26 105
use FILL  FILL_10804
timestamp 1680363874
transform 1 0 3960 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_634
timestamp 1680363874
transform 1 0 3968 0 1 170
box -8 -3 104 105
use INVX2  INVX2_721
timestamp 1680363874
transform -1 0 4080 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_412
timestamp 1680363874
transform 1 0 4080 0 1 170
box -8 -3 46 105
use FILL  FILL_10805
timestamp 1680363874
transform 1 0 4120 0 1 170
box -8 -3 16 105
use FILL  FILL_10806
timestamp 1680363874
transform 1 0 4128 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_413
timestamp 1680363874
transform -1 0 4176 0 1 170
box -8 -3 46 105
use INVX2  INVX2_722
timestamp 1680363874
transform 1 0 4176 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_635
timestamp 1680363874
transform 1 0 4192 0 1 170
box -8 -3 104 105
use FILL  FILL_10807
timestamp 1680363874
transform 1 0 4288 0 1 170
box -8 -3 16 105
use FILL  FILL_10808
timestamp 1680363874
transform 1 0 4296 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_414
timestamp 1680363874
transform 1 0 4304 0 1 170
box -8 -3 46 105
use FILL  FILL_10809
timestamp 1680363874
transform 1 0 4344 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_643
timestamp 1680363874
transform 1 0 4352 0 1 170
box -8 -3 104 105
use AOI22X1  AOI22X1_415
timestamp 1680363874
transform -1 0 4488 0 1 170
box -8 -3 46 105
use FILL  FILL_10833
timestamp 1680363874
transform 1 0 4488 0 1 170
box -8 -3 16 105
use FILL  FILL_10834
timestamp 1680363874
transform 1 0 4496 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_416
timestamp 1680363874
transform -1 0 4544 0 1 170
box -8 -3 46 105
use INVX2  INVX2_724
timestamp 1680363874
transform 1 0 4544 0 1 170
box -9 -3 26 105
use FILL  FILL_10835
timestamp 1680363874
transform 1 0 4560 0 1 170
box -8 -3 16 105
use FILL  FILL_10836
timestamp 1680363874
transform 1 0 4568 0 1 170
box -8 -3 16 105
use FILL  FILL_10837
timestamp 1680363874
transform 1 0 4576 0 1 170
box -8 -3 16 105
use FILL  FILL_10838
timestamp 1680363874
transform 1 0 4584 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_417
timestamp 1680363874
transform -1 0 4632 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_418
timestamp 1680363874
transform -1 0 4672 0 1 170
box -8 -3 46 105
use FILL  FILL_10839
timestamp 1680363874
transform 1 0 4672 0 1 170
box -8 -3 16 105
use FILL  FILL_10840
timestamp 1680363874
transform 1 0 4680 0 1 170
box -8 -3 16 105
use INVX2  INVX2_725
timestamp 1680363874
transform 1 0 4688 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_644
timestamp 1680363874
transform 1 0 4704 0 1 170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_91
timestamp 1680363874
transform 1 0 4827 0 1 170
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_92
timestamp 1680363874
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_10577
timestamp 1680363874
transform 1 0 72 0 -1 170
box -8 -3 16 105
use FILL  FILL_10579
timestamp 1680363874
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_10581
timestamp 1680363874
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_10583
timestamp 1680363874
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_10585
timestamp 1680363874
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_10587
timestamp 1680363874
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_10589
timestamp 1680363874
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_10591
timestamp 1680363874
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_10593
timestamp 1680363874
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_10595
timestamp 1680363874
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_10597
timestamp 1680363874
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_10599
timestamp 1680363874
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_10600
timestamp 1680363874
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_10601
timestamp 1680363874
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_10602
timestamp 1680363874
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_10603
timestamp 1680363874
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_10604
timestamp 1680363874
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_10605
timestamp 1680363874
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_10606
timestamp 1680363874
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_10607
timestamp 1680363874
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_10608
timestamp 1680363874
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_10609
timestamp 1680363874
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_10610
timestamp 1680363874
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_10611
timestamp 1680363874
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_10612
timestamp 1680363874
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_10613
timestamp 1680363874
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_10615
timestamp 1680363874
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_10617
timestamp 1680363874
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_10619
timestamp 1680363874
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_10621
timestamp 1680363874
transform 1 0 304 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8898
timestamp 1680363874
transform 1 0 404 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9950
timestamp 1680363874
transform 1 0 404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10014
timestamp 1680363874
transform 1 0 324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10015
timestamp 1680363874
transform 1 0 356 0 1 125
box -2 -2 2 2
use FILL  FILL_10624
timestamp 1680363874
transform 1 0 312 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_599
timestamp 1680363874
transform -1 0 416 0 -1 170
box -8 -3 104 105
use FILL  FILL_10625
timestamp 1680363874
transform 1 0 416 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8859
timestamp 1680363874
transform 1 0 436 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8860
timestamp 1680363874
transform 1 0 492 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8879
timestamp 1680363874
transform 1 0 484 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8899
timestamp 1680363874
transform 1 0 436 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9951
timestamp 1680363874
transform 1 0 436 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10016
timestamp 1680363874
transform 1 0 484 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_601
timestamp 1680363874
transform 1 0 424 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8931
timestamp 1680363874
transform 1 0 532 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10017
timestamp 1680363874
transform 1 0 532 0 1 125
box -2 -2 2 2
use FILL  FILL_10637
timestamp 1680363874
transform 1 0 520 0 -1 170
box -8 -3 16 105
use FILL  FILL_10638
timestamp 1680363874
transform 1 0 528 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8861
timestamp 1680363874
transform 1 0 556 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9952
timestamp 1680363874
transform 1 0 548 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8932
timestamp 1680363874
transform 1 0 596 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10018
timestamp 1680363874
transform 1 0 596 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8949
timestamp 1680363874
transform 1 0 596 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_602
timestamp 1680363874
transform 1 0 536 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8900
timestamp 1680363874
transform 1 0 644 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8880
timestamp 1680363874
transform 1 0 668 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8901
timestamp 1680363874
transform 1 0 692 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9953
timestamp 1680363874
transform 1 0 652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9954
timestamp 1680363874
transform 1 0 668 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9955
timestamp 1680363874
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9956
timestamp 1680363874
transform 1 0 692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10019
timestamp 1680363874
transform 1 0 644 0 1 125
box -2 -2 2 2
use FILL  FILL_10639
timestamp 1680363874
transform 1 0 632 0 -1 170
box -8 -3 16 105
use FILL  FILL_10640
timestamp 1680363874
transform 1 0 640 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10020
timestamp 1680363874
transform 1 0 660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10021
timestamp 1680363874
transform 1 0 676 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8945
timestamp 1680363874
transform 1 0 684 0 1 125
box -3 -3 3 3
use OAI22X1  OAI22X1_433
timestamp 1680363874
transform -1 0 688 0 -1 170
box -8 -3 46 105
use FILL  FILL_10641
timestamp 1680363874
transform 1 0 688 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8902
timestamp 1680363874
transform 1 0 708 0 1 145
box -3 -3 3 3
use FILL  FILL_10643
timestamp 1680363874
transform 1 0 696 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8881
timestamp 1680363874
transform 1 0 724 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8903
timestamp 1680363874
transform 1 0 756 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9957
timestamp 1680363874
transform 1 0 724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9958
timestamp 1680363874
transform 1 0 740 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9959
timestamp 1680363874
transform 1 0 756 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9960
timestamp 1680363874
transform 1 0 764 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10022
timestamp 1680363874
transform 1 0 716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10023
timestamp 1680363874
transform 1 0 732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10024
timestamp 1680363874
transform 1 0 748 0 1 125
box -2 -2 2 2
use INVX2  INVX2_691
timestamp 1680363874
transform 1 0 704 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_8950
timestamp 1680363874
transform 1 0 740 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8946
timestamp 1680363874
transform 1 0 764 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8972
timestamp 1680363874
transform 1 0 764 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_8976
timestamp 1680363874
transform 1 0 756 0 1 75
box -3 -3 3 3
use OAI22X1  OAI22X1_434
timestamp 1680363874
transform -1 0 760 0 -1 170
box -8 -3 46 105
use FILL  FILL_10647
timestamp 1680363874
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_10649
timestamp 1680363874
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10661
timestamp 1680363874
transform 1 0 776 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8882
timestamp 1680363874
transform 1 0 820 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8904
timestamp 1680363874
transform 1 0 804 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9961
timestamp 1680363874
transform 1 0 804 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9962
timestamp 1680363874
transform 1 0 820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10025
timestamp 1680363874
transform 1 0 812 0 1 125
box -2 -2 2 2
use OAI22X1  OAI22X1_436
timestamp 1680363874
transform 1 0 784 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_8862
timestamp 1680363874
transform 1 0 916 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8905
timestamp 1680363874
transform 1 0 868 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9963
timestamp 1680363874
transform 1 0 916 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10026
timestamp 1680363874
transform 1 0 836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10027
timestamp 1680363874
transform 1 0 868 0 1 125
box -2 -2 2 2
use FILL  FILL_10662
timestamp 1680363874
transform 1 0 824 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_604
timestamp 1680363874
transform -1 0 928 0 -1 170
box -8 -3 104 105
use FILL  FILL_10663
timestamp 1680363874
transform 1 0 928 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8863
timestamp 1680363874
transform 1 0 948 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8864
timestamp 1680363874
transform 1 0 1004 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8883
timestamp 1680363874
transform 1 0 996 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9964
timestamp 1680363874
transform 1 0 948 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8933
timestamp 1680363874
transform 1 0 996 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8934
timestamp 1680363874
transform 1 0 1028 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10028
timestamp 1680363874
transform 1 0 996 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_605
timestamp 1680363874
transform 1 0 936 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10029
timestamp 1680363874
transform 1 0 1044 0 1 125
box -2 -2 2 2
use INVX2  INVX2_693
timestamp 1680363874
transform 1 0 1032 0 -1 170
box -9 -3 26 105
use FILL  FILL_10664
timestamp 1680363874
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_10666
timestamp 1680363874
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8865
timestamp 1680363874
transform 1 0 1084 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8884
timestamp 1680363874
transform 1 0 1076 0 1 155
box -3 -3 3 3
use FILL  FILL_10668
timestamp 1680363874
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8906
timestamp 1680363874
transform 1 0 1132 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9965
timestamp 1680363874
transform 1 0 1084 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10030
timestamp 1680363874
transform 1 0 1132 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_608
timestamp 1680363874
transform 1 0 1072 0 -1 170
box -8 -3 104 105
use FILL  FILL_10680
timestamp 1680363874
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use FILL  FILL_10681
timestamp 1680363874
transform 1 0 1176 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8885
timestamp 1680363874
transform 1 0 1204 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8907
timestamp 1680363874
transform 1 0 1220 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9966
timestamp 1680363874
transform 1 0 1204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9967
timestamp 1680363874
transform 1 0 1220 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9968
timestamp 1680363874
transform 1 0 1236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10031
timestamp 1680363874
transform 1 0 1196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10032
timestamp 1680363874
transform 1 0 1212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10033
timestamp 1680363874
transform 1 0 1228 0 1 125
box -2 -2 2 2
use INVX2  INVX2_694
timestamp 1680363874
transform 1 0 1184 0 -1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_438
timestamp 1680363874
transform -1 0 1240 0 -1 170
box -8 -3 46 105
use FILL  FILL_10682
timestamp 1680363874
transform 1 0 1240 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8866
timestamp 1680363874
transform 1 0 1260 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9969
timestamp 1680363874
transform 1 0 1260 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8935
timestamp 1680363874
transform 1 0 1308 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10034
timestamp 1680363874
transform 1 0 1308 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_609
timestamp 1680363874
transform 1 0 1248 0 -1 170
box -8 -3 104 105
use FILL  FILL_10683
timestamp 1680363874
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8936
timestamp 1680363874
transform 1 0 1364 0 1 135
box -3 -3 3 3
use FILL  FILL_10684
timestamp 1680363874
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10035
timestamp 1680363874
transform 1 0 1372 0 1 125
box -2 -2 2 2
use INVX2  INVX2_695
timestamp 1680363874
transform 1 0 1360 0 -1 170
box -9 -3 26 105
use FILL  FILL_10685
timestamp 1680363874
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_10686
timestamp 1680363874
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use FILL  FILL_10688
timestamp 1680363874
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_10690
timestamp 1680363874
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8867
timestamp 1680363874
transform 1 0 1420 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8868
timestamp 1680363874
transform 1 0 1468 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8908
timestamp 1680363874
transform 1 0 1420 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9970
timestamp 1680363874
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10036
timestamp 1680363874
transform 1 0 1468 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_615
timestamp 1680363874
transform 1 0 1408 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_704
timestamp 1680363874
transform 1 0 1504 0 -1 170
box -9 -3 26 105
use FILL  FILL_10713
timestamp 1680363874
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8869
timestamp 1680363874
transform 1 0 1548 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_10037
timestamp 1680363874
transform 1 0 1540 0 1 125
box -2 -2 2 2
use FILL  FILL_10714
timestamp 1680363874
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use FILL  FILL_10715
timestamp 1680363874
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8886
timestamp 1680363874
transform 1 0 1620 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9971
timestamp 1680363874
transform 1 0 1556 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8937
timestamp 1680363874
transform 1 0 1604 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10038
timestamp 1680363874
transform 1 0 1604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10039
timestamp 1680363874
transform 1 0 1636 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_616
timestamp 1680363874
transform 1 0 1544 0 -1 170
box -8 -3 104 105
use FILL  FILL_10716
timestamp 1680363874
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8938
timestamp 1680363874
transform 1 0 1660 0 1 135
box -3 -3 3 3
use FILL  FILL_10717
timestamp 1680363874
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_10718
timestamp 1680363874
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_10719
timestamp 1680363874
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9972
timestamp 1680363874
transform 1 0 1684 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8939
timestamp 1680363874
transform 1 0 1732 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8940
timestamp 1680363874
transform 1 0 1756 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10040
timestamp 1680363874
transform 1 0 1732 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_617
timestamp 1680363874
transform 1 0 1672 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10041
timestamp 1680363874
transform 1 0 1780 0 1 125
box -2 -2 2 2
use FILL  FILL_10720
timestamp 1680363874
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10721
timestamp 1680363874
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8909
timestamp 1680363874
transform 1 0 1796 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9973
timestamp 1680363874
transform 1 0 1796 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8941
timestamp 1680363874
transform 1 0 1844 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10042
timestamp 1680363874
transform 1 0 1844 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_618
timestamp 1680363874
transform 1 0 1784 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10043
timestamp 1680363874
transform 1 0 1892 0 1 125
box -2 -2 2 2
use FILL  FILL_10722
timestamp 1680363874
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_10723
timestamp 1680363874
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8870
timestamp 1680363874
transform 1 0 1916 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8910
timestamp 1680363874
transform 1 0 1908 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8911
timestamp 1680363874
transform 1 0 1988 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9974
timestamp 1680363874
transform 1 0 1908 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8942
timestamp 1680363874
transform 1 0 1940 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8871
timestamp 1680363874
transform 1 0 2028 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8912
timestamp 1680363874
transform 1 0 2036 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9975
timestamp 1680363874
transform 1 0 1996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9976
timestamp 1680363874
transform 1 0 2012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9977
timestamp 1680363874
transform 1 0 2028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9978
timestamp 1680363874
transform 1 0 2036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10044
timestamp 1680363874
transform 1 0 1948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10045
timestamp 1680363874
transform 1 0 1988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10046
timestamp 1680363874
transform 1 0 2004 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10047
timestamp 1680363874
transform 1 0 2020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10048
timestamp 1680363874
transform 1 0 2036 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8951
timestamp 1680363874
transform 1 0 1948 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8952
timestamp 1680363874
transform 1 0 2012 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8974
timestamp 1680363874
transform 1 0 1996 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_619
timestamp 1680363874
transform 1 0 1896 0 -1 170
box -8 -3 104 105
use OAI22X1  OAI22X1_446
timestamp 1680363874
transform 1 0 1992 0 -1 170
box -8 -3 46 105
use INVX2  INVX2_705
timestamp 1680363874
transform 1 0 2032 0 -1 170
box -9 -3 26 105
use FILL  FILL_10724
timestamp 1680363874
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8872
timestamp 1680363874
transform 1 0 2068 0 1 165
box -3 -3 3 3
use FILL  FILL_10725
timestamp 1680363874
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_10726
timestamp 1680363874
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_10727
timestamp 1680363874
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8873
timestamp 1680363874
transform 1 0 2092 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9979
timestamp 1680363874
transform 1 0 2092 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8943
timestamp 1680363874
transform 1 0 2140 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8944
timestamp 1680363874
transform 1 0 2172 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10049
timestamp 1680363874
transform 1 0 2140 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_620
timestamp 1680363874
transform 1 0 2080 0 -1 170
box -8 -3 104 105
use FILL  FILL_10728
timestamp 1680363874
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9980
timestamp 1680363874
transform 1 0 2196 0 1 135
box -2 -2 2 2
use FILL  FILL_10729
timestamp 1680363874
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_10730
timestamp 1680363874
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9981
timestamp 1680363874
transform 1 0 2292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10050
timestamp 1680363874
transform 1 0 2212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10051
timestamp 1680363874
transform 1 0 2252 0 1 125
box -2 -2 2 2
use FILL  FILL_10731
timestamp 1680363874
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_621
timestamp 1680363874
transform -1 0 2304 0 -1 170
box -8 -3 104 105
use FILL  FILL_10732
timestamp 1680363874
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_10733
timestamp 1680363874
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8874
timestamp 1680363874
transform 1 0 2332 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9982
timestamp 1680363874
transform 1 0 2332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10052
timestamp 1680363874
transform 1 0 2380 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8953
timestamp 1680363874
transform 1 0 2380 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8913
timestamp 1680363874
transform 1 0 2420 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8914
timestamp 1680363874
transform 1 0 2468 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9983
timestamp 1680363874
transform 1 0 2428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9984
timestamp 1680363874
transform 1 0 2444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9985
timestamp 1680363874
transform 1 0 2460 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9986
timestamp 1680363874
transform 1 0 2468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10053
timestamp 1680363874
transform 1 0 2420 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_622
timestamp 1680363874
transform 1 0 2320 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10054
timestamp 1680363874
transform 1 0 2436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10055
timestamp 1680363874
transform 1 0 2452 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8954
timestamp 1680363874
transform 1 0 2444 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8977
timestamp 1680363874
transform 1 0 2428 0 1 75
box -3 -3 3 3
use FILL  FILL_10734
timestamp 1680363874
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10056
timestamp 1680363874
transform 1 0 2468 0 1 125
box -2 -2 2 2
use OAI22X1  OAI22X1_447
timestamp 1680363874
transform 1 0 2424 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_8975
timestamp 1680363874
transform 1 0 2476 0 1 85
box -3 -3 3 3
use FILL  FILL_10735
timestamp 1680363874
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8875
timestamp 1680363874
transform 1 0 2500 0 1 165
box -3 -3 3 3
use INVX2  INVX2_706
timestamp 1680363874
transform 1 0 2472 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_10057
timestamp 1680363874
transform 1 0 2500 0 1 125
box -2 -2 2 2
use FILL  FILL_10745
timestamp 1680363874
transform 1 0 2488 0 -1 170
box -8 -3 16 105
use FILL  FILL_10746
timestamp 1680363874
transform 1 0 2496 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8876
timestamp 1680363874
transform 1 0 2564 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8915
timestamp 1680363874
transform 1 0 2564 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9987
timestamp 1680363874
transform 1 0 2516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10058
timestamp 1680363874
transform 1 0 2564 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8887
timestamp 1680363874
transform 1 0 2604 0 1 155
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_623
timestamp 1680363874
transform 1 0 2504 0 -1 170
box -8 -3 104 105
use FILL  FILL_10747
timestamp 1680363874
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8916
timestamp 1680363874
transform 1 0 2620 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8947
timestamp 1680363874
transform 1 0 2620 0 1 125
box -3 -3 3 3
use FILL  FILL_10748
timestamp 1680363874
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_10749
timestamp 1680363874
transform 1 0 2616 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9988
timestamp 1680363874
transform 1 0 2644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10059
timestamp 1680363874
transform 1 0 2636 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8948
timestamp 1680363874
transform 1 0 2652 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8917
timestamp 1680363874
transform 1 0 2676 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8918
timestamp 1680363874
transform 1 0 2732 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9989
timestamp 1680363874
transform 1 0 2676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9990
timestamp 1680363874
transform 1 0 2692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9991
timestamp 1680363874
transform 1 0 2708 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10060
timestamp 1680363874
transform 1 0 2660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10061
timestamp 1680363874
transform 1 0 2684 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8973
timestamp 1680363874
transform 1 0 2644 0 1 105
box -3 -3 3 3
use INVX2  INVX2_707
timestamp 1680363874
transform 1 0 2624 0 -1 170
box -9 -3 26 105
use FILL  FILL_10750
timestamp 1680363874
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_10773
timestamp 1680363874
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8955
timestamp 1680363874
transform 1 0 2684 0 1 115
box -3 -3 3 3
use OAI22X1  OAI22X1_452
timestamp 1680363874
transform 1 0 2656 0 -1 170
box -8 -3 46 105
use M2_M1  M2_M1_10062
timestamp 1680363874
transform 1 0 2732 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8956
timestamp 1680363874
transform 1 0 2772 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_625
timestamp 1680363874
transform 1 0 2696 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10063
timestamp 1680363874
transform 1 0 2804 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8957
timestamp 1680363874
transform 1 0 2804 0 1 115
box -3 -3 3 3
use INVX2  INVX2_711
timestamp 1680363874
transform 1 0 2792 0 -1 170
box -9 -3 26 105
use FILL  FILL_10774
timestamp 1680363874
transform 1 0 2808 0 -1 170
box -8 -3 16 105
use FILL  FILL_10775
timestamp 1680363874
transform 1 0 2816 0 -1 170
box -8 -3 16 105
use FILL  FILL_10776
timestamp 1680363874
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8877
timestamp 1680363874
transform 1 0 2844 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9992
timestamp 1680363874
transform 1 0 2844 0 1 135
box -2 -2 2 2
use FILL  FILL_10777
timestamp 1680363874
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8878
timestamp 1680363874
transform 1 0 2884 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8919
timestamp 1680363874
transform 1 0 2940 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9993
timestamp 1680363874
transform 1 0 2940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10064
timestamp 1680363874
transform 1 0 2852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10065
timestamp 1680363874
transform 1 0 2860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10066
timestamp 1680363874
transform 1 0 2892 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8958
timestamp 1680363874
transform 1 0 2852 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8959
timestamp 1680363874
transform 1 0 2892 0 1 115
box -3 -3 3 3
use INVX2  INVX2_712
timestamp 1680363874
transform 1 0 2840 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_9994
timestamp 1680363874
transform 1 0 2956 0 1 135
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_626
timestamp 1680363874
transform -1 0 2952 0 -1 170
box -8 -3 104 105
use FILL  FILL_10778
timestamp 1680363874
transform 1 0 2952 0 -1 170
box -8 -3 16 105
use FILL  FILL_10779
timestamp 1680363874
transform 1 0 2960 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8920
timestamp 1680363874
transform 1 0 2996 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9995
timestamp 1680363874
transform 1 0 2996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10067
timestamp 1680363874
transform 1 0 2980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10068
timestamp 1680363874
transform 1 0 3020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10069
timestamp 1680363874
transform 1 0 3076 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8960
timestamp 1680363874
transform 1 0 2980 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8961
timestamp 1680363874
transform 1 0 3020 0 1 115
box -3 -3 3 3
use INVX2  INVX2_713
timestamp 1680363874
transform 1 0 2968 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_627
timestamp 1680363874
transform 1 0 2984 0 -1 170
box -8 -3 104 105
use FILL  FILL_10780
timestamp 1680363874
transform 1 0 3080 0 -1 170
box -8 -3 16 105
use FILL  FILL_10781
timestamp 1680363874
transform 1 0 3088 0 -1 170
box -8 -3 16 105
use FILL  FILL_10782
timestamp 1680363874
transform 1 0 3096 0 -1 170
box -8 -3 16 105
use FILL  FILL_10783
timestamp 1680363874
transform 1 0 3104 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8921
timestamp 1680363874
transform 1 0 3124 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9996
timestamp 1680363874
transform 1 0 3124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9997
timestamp 1680363874
transform 1 0 3212 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10070
timestamp 1680363874
transform 1 0 3172 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10071
timestamp 1680363874
transform 1 0 3204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10072
timestamp 1680363874
transform 1 0 3212 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8962
timestamp 1680363874
transform 1 0 3172 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8963
timestamp 1680363874
transform 1 0 3212 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_628
timestamp 1680363874
transform 1 0 3112 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_714
timestamp 1680363874
transform 1 0 3208 0 -1 170
box -9 -3 26 105
use FILL  FILL_10784
timestamp 1680363874
transform 1 0 3224 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8922
timestamp 1680363874
transform 1 0 3268 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8923
timestamp 1680363874
transform 1 0 3316 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8924
timestamp 1680363874
transform 1 0 3348 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9998
timestamp 1680363874
transform 1 0 3244 0 1 135
box -2 -2 2 2
use FILL  FILL_10785
timestamp 1680363874
transform 1 0 3232 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9999
timestamp 1680363874
transform 1 0 3268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10073
timestamp 1680363874
transform 1 0 3252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10074
timestamp 1680363874
transform 1 0 3292 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10075
timestamp 1680363874
transform 1 0 3348 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8964
timestamp 1680363874
transform 1 0 3252 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8965
timestamp 1680363874
transform 1 0 3292 0 1 115
box -3 -3 3 3
use INVX2  INVX2_715
timestamp 1680363874
transform 1 0 3240 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_629
timestamp 1680363874
transform 1 0 3256 0 -1 170
box -8 -3 104 105
use FILL  FILL_10786
timestamp 1680363874
transform 1 0 3352 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10076
timestamp 1680363874
transform 1 0 3372 0 1 125
box -2 -2 2 2
use FILL  FILL_10787
timestamp 1680363874
transform 1 0 3360 0 -1 170
box -8 -3 16 105
use FILL  FILL_10788
timestamp 1680363874
transform 1 0 3368 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8888
timestamp 1680363874
transform 1 0 3460 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10000
timestamp 1680363874
transform 1 0 3460 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10077
timestamp 1680363874
transform 1 0 3412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10078
timestamp 1680363874
transform 1 0 3476 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_630
timestamp 1680363874
transform -1 0 3472 0 -1 170
box -8 -3 104 105
use FILL  FILL_10789
timestamp 1680363874
transform 1 0 3472 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8889
timestamp 1680363874
transform 1 0 3548 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8890
timestamp 1680363874
transform 1 0 3572 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8925
timestamp 1680363874
transform 1 0 3492 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8926
timestamp 1680363874
transform 1 0 3524 0 1 145
box -3 -3 3 3
use FILL  FILL_10810
timestamp 1680363874
transform 1 0 3480 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10001
timestamp 1680363874
transform 1 0 3572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10079
timestamp 1680363874
transform 1 0 3524 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_636
timestamp 1680363874
transform -1 0 3584 0 -1 170
box -8 -3 104 105
use FILL  FILL_10811
timestamp 1680363874
transform 1 0 3584 0 -1 170
box -8 -3 16 105
use FILL  FILL_10812
timestamp 1680363874
transform 1 0 3592 0 -1 170
box -8 -3 16 105
use FILL  FILL_10813
timestamp 1680363874
transform 1 0 3600 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8927
timestamp 1680363874
transform 1 0 3620 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_10002
timestamp 1680363874
transform 1 0 3620 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10080
timestamp 1680363874
transform 1 0 3644 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_637
timestamp 1680363874
transform 1 0 3608 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10081
timestamp 1680363874
transform 1 0 3716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10082
timestamp 1680363874
transform 1 0 3724 0 1 125
box -2 -2 2 2
use FILL  FILL_10814
timestamp 1680363874
transform 1 0 3704 0 -1 170
box -8 -3 16 105
use FILL  FILL_10815
timestamp 1680363874
transform 1 0 3712 0 -1 170
box -8 -3 16 105
use FILL  FILL_10816
timestamp 1680363874
transform 1 0 3720 0 -1 170
box -8 -3 16 105
use FILL  FILL_10817
timestamp 1680363874
transform 1 0 3728 0 -1 170
box -8 -3 16 105
use FILL  FILL_10818
timestamp 1680363874
transform 1 0 3736 0 -1 170
box -8 -3 16 105
use FILL  FILL_10819
timestamp 1680363874
transform 1 0 3744 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8891
timestamp 1680363874
transform 1 0 3836 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10003
timestamp 1680363874
transform 1 0 3836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10083
timestamp 1680363874
transform 1 0 3804 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_638
timestamp 1680363874
transform -1 0 3848 0 -1 170
box -8 -3 104 105
use FILL  FILL_10820
timestamp 1680363874
transform 1 0 3848 0 -1 170
box -8 -3 16 105
use FILL  FILL_10821
timestamp 1680363874
transform 1 0 3856 0 -1 170
box -8 -3 16 105
use FILL  FILL_10822
timestamp 1680363874
transform 1 0 3864 0 -1 170
box -8 -3 16 105
use FILL  FILL_10823
timestamp 1680363874
transform 1 0 3872 0 -1 170
box -8 -3 16 105
use FILL  FILL_10824
timestamp 1680363874
transform 1 0 3880 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8928
timestamp 1680363874
transform 1 0 3900 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_10004
timestamp 1680363874
transform 1 0 3900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10084
timestamp 1680363874
transform 1 0 3932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10085
timestamp 1680363874
transform 1 0 3980 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_639
timestamp 1680363874
transform 1 0 3888 0 -1 170
box -8 -3 104 105
use FILL  FILL_10825
timestamp 1680363874
transform 1 0 3984 0 -1 170
box -8 -3 16 105
use FILL  FILL_10826
timestamp 1680363874
transform 1 0 3992 0 -1 170
box -8 -3 16 105
use FILL  FILL_10827
timestamp 1680363874
transform 1 0 4000 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8892
timestamp 1680363874
transform 1 0 4020 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10005
timestamp 1680363874
transform 1 0 4020 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10086
timestamp 1680363874
transform 1 0 4068 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10087
timestamp 1680363874
transform 1 0 4108 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_640
timestamp 1680363874
transform 1 0 4008 0 -1 170
box -8 -3 104 105
use FILL  FILL_10828
timestamp 1680363874
transform 1 0 4104 0 -1 170
box -8 -3 16 105
use FILL  FILL_10829
timestamp 1680363874
transform 1 0 4112 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8893
timestamp 1680363874
transform 1 0 4212 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10006
timestamp 1680363874
transform 1 0 4212 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10088
timestamp 1680363874
transform 1 0 4132 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10089
timestamp 1680363874
transform 1 0 4188 0 1 125
box -2 -2 2 2
use FILL  FILL_10830
timestamp 1680363874
transform 1 0 4120 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_641
timestamp 1680363874
transform -1 0 4224 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8894
timestamp 1680363874
transform 1 0 4236 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10007
timestamp 1680363874
transform 1 0 4236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10008
timestamp 1680363874
transform 1 0 4324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10090
timestamp 1680363874
transform 1 0 4284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10091
timestamp 1680363874
transform 1 0 4316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10092
timestamp 1680363874
transform 1 0 4324 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8966
timestamp 1680363874
transform 1 0 4284 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8967
timestamp 1680363874
transform 1 0 4324 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_642
timestamp 1680363874
transform 1 0 4224 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_723
timestamp 1680363874
transform 1 0 4320 0 -1 170
box -9 -3 26 105
use FILL  FILL_10831
timestamp 1680363874
transform 1 0 4336 0 -1 170
box -8 -3 16 105
use FILL  FILL_10832
timestamp 1680363874
transform 1 0 4344 0 -1 170
box -8 -3 16 105
use FILL  FILL_10841
timestamp 1680363874
transform 1 0 4352 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8895
timestamp 1680363874
transform 1 0 4372 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10009
timestamp 1680363874
transform 1 0 4372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10010
timestamp 1680363874
transform 1 0 4468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10093
timestamp 1680363874
transform 1 0 4420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10094
timestamp 1680363874
transform 1 0 4452 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10095
timestamp 1680363874
transform 1 0 4460 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8968
timestamp 1680363874
transform 1 0 4420 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8969
timestamp 1680363874
transform 1 0 4460 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_645
timestamp 1680363874
transform 1 0 4360 0 -1 170
box -8 -3 104 105
use FILL  FILL_10842
timestamp 1680363874
transform 1 0 4456 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_726
timestamp 1680363874
transform 1 0 4464 0 -1 170
box -9 -3 26 105
use FILL  FILL_10843
timestamp 1680363874
transform 1 0 4480 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8896
timestamp 1680363874
transform 1 0 4588 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8929
timestamp 1680363874
transform 1 0 4580 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8897
timestamp 1680363874
transform 1 0 4700 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8930
timestamp 1680363874
transform 1 0 4620 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_10011
timestamp 1680363874
transform 1 0 4580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10012
timestamp 1680363874
transform 1 0 4596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10096
timestamp 1680363874
transform 1 0 4500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10097
timestamp 1680363874
transform 1 0 4556 0 1 125
box -2 -2 2 2
use FILL  FILL_10844
timestamp 1680363874
transform 1 0 4488 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_646
timestamp 1680363874
transform -1 0 4592 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10013
timestamp 1680363874
transform 1 0 4620 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10098
timestamp 1680363874
transform 1 0 4604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10099
timestamp 1680363874
transform 1 0 4644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10100
timestamp 1680363874
transform 1 0 4700 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8970
timestamp 1680363874
transform 1 0 4604 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8971
timestamp 1680363874
transform 1 0 4644 0 1 115
box -3 -3 3 3
use INVX2  INVX2_727
timestamp 1680363874
transform 1 0 4592 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_647
timestamp 1680363874
transform 1 0 4608 0 -1 170
box -8 -3 104 105
use FILL  FILL_10845
timestamp 1680363874
transform 1 0 4704 0 -1 170
box -8 -3 16 105
use FILL  FILL_10846
timestamp 1680363874
transform 1 0 4712 0 -1 170
box -8 -3 16 105
use FILL  FILL_10847
timestamp 1680363874
transform 1 0 4720 0 -1 170
box -8 -3 16 105
use FILL  FILL_10848
timestamp 1680363874
transform 1 0 4728 0 -1 170
box -8 -3 16 105
use FILL  FILL_10849
timestamp 1680363874
transform 1 0 4736 0 -1 170
box -8 -3 16 105
use FILL  FILL_10850
timestamp 1680363874
transform 1 0 4744 0 -1 170
box -8 -3 16 105
use FILL  FILL_10851
timestamp 1680363874
transform 1 0 4752 0 -1 170
box -8 -3 16 105
use FILL  FILL_10852
timestamp 1680363874
transform 1 0 4760 0 -1 170
box -8 -3 16 105
use FILL  FILL_10853
timestamp 1680363874
transform 1 0 4768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10854
timestamp 1680363874
transform 1 0 4776 0 -1 170
box -8 -3 16 105
use FILL  FILL_10855
timestamp 1680363874
transform 1 0 4784 0 -1 170
box -8 -3 16 105
use FILL  FILL_10856
timestamp 1680363874
transform 1 0 4792 0 -1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_93
timestamp 1680363874
transform 1 0 4851 0 1 70
box -10 -3 10 3
use top_level_VIA1  top_level_VIA1_4
timestamp 1680363874
transform 1 0 48 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_8978
timestamp 1680363874
transform 1 0 1284 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_8979
timestamp 1680363874
transform 1 0 2788 0 1 55
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_6
timestamp 1680363874
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_8980
timestamp 1680363874
transform 1 0 1068 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_8981
timestamp 1680363874
transform 1 0 3028 0 1 35
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_5
timestamp 1680363874
transform 1 0 4827 0 1 47
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_7
timestamp 1680363874
transform 1 0 4851 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal3 2 2525 2 2525 4 clka
rlabel metal2 2228 4738 2228 4738 4 clkb
rlabel metal3 2 1155 2 1155 4 reset
rlabel metal2 2620 1 2620 1 4 we_ins
rlabel metal2 4052 4738 4052 4738 4 load[15]
rlabel metal2 3932 4738 3932 4738 4 load[14]
rlabel metal2 3820 4738 3820 4738 4 load[13]
rlabel metal2 3700 4738 3700 4738 4 load[12]
rlabel metal2 3684 4738 3684 4738 4 load[11]
rlabel metal2 3788 4738 3788 4738 4 load[10]
rlabel metal3 4875 3725 4875 3725 4 load[9]
rlabel metal2 4196 4738 4196 4738 4 load[8]
rlabel metal3 4875 4525 4875 4525 4 load[7]
rlabel metal3 4875 4615 4875 4615 4 load[6]
rlabel metal3 4875 3925 4875 3925 4 load[5]
rlabel metal3 4875 4125 4875 4125 4 load[4]
rlabel metal3 4875 4215 4875 4215 4 load[3]
rlabel metal3 4875 4415 4875 4415 4 load[2]
rlabel metal2 4644 4738 4644 4738 4 load[1]
rlabel metal2 3884 4738 3884 4738 4 load[0]
rlabel metal3 2 4375 2 4375 4 reg_0_out[7]
rlabel metal3 2 4135 2 4135 4 reg_0_out[6]
rlabel metal3 2 4215 2 4215 4 reg_0_out[5]
rlabel metal3 2 4575 2 4575 4 reg_0_out[4]
rlabel metal2 732 4738 732 4738 4 reg_0_out[3]
rlabel metal2 276 4738 276 4738 4 reg_0_out[2]
rlabel metal2 548 4738 548 4738 4 reg_0_out[1]
rlabel metal3 2 3965 2 3965 4 reg_0_out[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>

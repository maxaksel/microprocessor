magic
tech scmos
timestamp 1680464795
<< m2contact >>
rect -2 -2 2 2
<< end >>

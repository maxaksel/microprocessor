magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -7 48 39 105
<< ntransistor >>
rect 10 6 12 26
rect 15 6 17 26
rect 23 6 25 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 5 6 10 26
rect 12 6 15 26
rect 17 16 22 26
rect 17 6 23 16
rect 25 6 30 16
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 15 94
rect 17 54 23 94
rect 25 54 30 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 49 9 54
rect 6 47 10 49
rect 4 45 10 47
rect 4 29 6 45
rect 15 41 17 54
rect 10 37 17 41
rect 4 27 12 29
rect 10 26 12 27
rect 15 26 17 37
rect 23 23 25 54
rect 23 19 29 23
rect 23 16 25 19
rect 10 4 12 6
rect 15 4 17 6
rect 23 4 25 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 11 91 13 93
rect 3 89 5 91
rect 19 90 21 92
rect 27 90 29 92
rect 11 86 13 88
rect 3 84 5 86
rect 19 85 21 87
rect 27 85 29 87
rect 11 81 13 83
rect 3 79 5 81
rect 19 80 21 82
rect 27 80 29 82
rect 11 76 13 78
rect 3 74 5 76
rect 19 75 21 77
rect 27 75 29 77
rect 11 71 13 73
rect 3 69 5 71
rect 19 70 21 72
rect 27 70 29 72
rect 11 66 13 68
rect 3 64 5 66
rect 19 65 21 67
rect 27 65 29 67
rect 11 61 13 63
rect 3 59 5 61
rect 19 60 21 62
rect 27 60 29 62
rect 19 55 21 57
rect 27 55 29 57
rect 7 46 9 48
rect 11 38 13 40
rect 6 22 8 24
rect 19 22 21 24
rect 26 20 28 22
rect 6 17 8 19
rect 19 17 21 19
rect 6 12 8 14
rect 19 12 21 14
rect 27 12 29 14
rect 6 7 8 9
rect 19 7 21 9
rect 27 7 29 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 34 103
rect 2 57 6 94
rect 10 60 14 97
rect 18 57 22 94
rect 2 54 22 57
rect 26 54 30 94
rect 6 47 10 49
rect 26 47 29 54
rect 2 44 10 47
rect 18 44 30 47
rect 2 43 6 44
rect 10 33 14 41
rect 18 26 21 44
rect 26 43 30 44
rect 5 3 9 26
rect 18 6 22 26
rect 26 23 30 27
rect 25 19 29 23
rect 26 3 30 16
rect -2 -3 34 3
<< m1p >>
rect 2 43 6 47
rect 26 43 30 47
rect 10 33 14 37
rect 26 23 30 27
<< labels >>
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 45 4 45 6 A
rlabel metal1 12 35 12 35 6 B
rlabel metal1 28 45 28 45 6 Y
rlabel metal1 28 25 28 25 6 C
<< end >>

magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 16 105
<< psubstratepdiff >>
rect -2 -2 2 2
rect 6 -2 10 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 6 98 10 102
<< genericcontact >>
rect -1 99 1 101
rect 7 99 9 101
rect -1 -1 1 1
rect 7 -1 9 1
<< metal1 >>
rect -2 97 10 103
rect -2 -3 10 3
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
<< end >>

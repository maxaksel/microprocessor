magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 36
rect 12 6 14 36
rect 17 6 19 36
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
<< ndiffusion >>
rect 2 6 7 36
rect 9 6 12 36
rect 14 6 17 36
rect 19 6 24 36
<< pdiffusion >>
rect 2 74 7 94
rect 9 74 15 94
rect 17 74 23 94
rect 25 74 30 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 53 9 74
rect 15 73 17 74
rect 2 49 9 53
rect 7 36 9 49
rect 12 71 17 73
rect 12 47 14 71
rect 23 63 25 74
rect 18 59 25 63
rect 12 43 18 47
rect 12 36 14 43
rect 23 39 25 59
rect 17 37 25 39
rect 17 36 19 37
rect 7 4 9 6
rect 12 4 14 6
rect 17 4 19 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 11 90 13 92
rect 19 89 21 91
rect 27 90 29 92
rect 3 85 5 87
rect 11 85 13 87
rect 19 84 21 86
rect 27 85 29 87
rect 3 80 5 82
rect 11 80 13 82
rect 19 79 21 81
rect 27 80 29 82
rect 3 75 5 77
rect 11 75 13 77
rect 27 75 29 77
rect 19 60 21 62
rect 3 50 5 52
rect 15 44 17 46
rect 3 32 5 34
rect 21 32 23 34
rect 3 27 5 29
rect 21 27 23 29
rect 3 22 5 24
rect 21 22 23 24
rect 3 17 5 19
rect 21 17 23 19
rect 3 12 5 14
rect 21 12 23 14
rect 3 7 5 9
rect 21 7 23 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 34 103
rect 2 74 6 97
rect 10 74 14 94
rect 18 76 22 97
rect 11 73 14 74
rect 26 74 30 94
rect 26 73 29 74
rect 11 70 29 73
rect 18 59 22 67
rect 26 57 29 70
rect 2 49 6 57
rect 26 53 30 57
rect 10 43 18 47
rect 26 37 29 53
rect 21 36 29 37
rect 2 3 6 36
rect 20 34 29 36
rect 20 6 24 34
rect -2 -3 34 3
<< m1p >>
rect 18 63 22 67
rect 2 53 6 57
rect 26 53 30 57
rect 10 43 14 47
<< labels >>
rlabel metal1 12 45 12 45 6 B
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 55 4 55 6 A
rlabel metal1 20 65 20 65 6 C
rlabel metal1 28 55 28 55 6 Y
<< end >>

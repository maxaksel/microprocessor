magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
<< ndiffusion >>
rect 2 6 7 16
rect 9 6 15 16
rect 17 6 22 16
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 12 94
rect 14 54 19 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 7 23 9 54
rect 12 53 14 54
rect 12 51 17 53
rect 2 19 9 23
rect 7 16 9 19
rect 15 47 22 51
rect 15 16 17 47
rect 7 4 9 6
rect 15 4 17 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 16 90 18 92
rect 3 85 5 87
rect 16 85 18 87
rect 3 80 5 82
rect 16 80 18 82
rect 3 75 5 77
rect 16 75 18 77
rect 3 70 5 72
rect 16 70 18 72
rect 3 65 5 67
rect 16 65 18 67
rect 3 60 5 62
rect 16 60 18 62
rect 3 55 5 57
rect 16 55 18 57
rect 19 48 21 50
rect 3 20 5 22
rect 3 12 5 14
rect 11 12 13 14
rect 19 12 21 14
rect 3 7 5 9
rect 11 7 13 9
rect 19 7 21 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 26 103
rect 2 54 6 97
rect 15 58 19 94
rect 10 54 19 58
rect 11 37 14 54
rect 18 43 22 51
rect 10 33 14 37
rect 2 19 6 27
rect 11 16 14 33
rect 2 3 6 16
rect 10 6 14 16
rect 18 3 22 16
rect -2 -3 26 3
<< m1p >>
rect 18 43 22 47
rect 10 33 14 37
rect 2 23 6 27
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 20 45 20 45 6 B
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 12 35 12 35 6 Y
rlabel metal1 4 25 4 25 6 A
<< end >>

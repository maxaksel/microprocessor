magic
tech scmos
timestamp 1677622389
<< metal1 >>
rect 14 4707 4853 4727
rect 38 4683 4829 4703
rect 14 4667 4853 4673
rect 964 4623 981 4626
rect 2852 4623 2861 4626
rect 2892 4623 2901 4626
rect 2922 4623 2932 4626
rect 636 4613 661 4616
rect 698 4613 708 4616
rect 788 4613 813 4616
rect 850 4613 860 4616
rect 938 4613 948 4616
rect 1020 4613 1045 4616
rect 1090 4613 1100 4616
rect 1164 4613 1181 4616
rect 1218 4613 1244 4616
rect 1332 4613 1357 4616
rect 1444 4613 1469 4616
rect 1500 4613 1517 4616
rect 1604 4613 1613 4616
rect 1666 4613 1797 4616
rect 1836 4613 1861 4616
rect 1898 4613 1916 4616
rect 1980 4613 2005 4616
rect 2042 4613 2060 4616
rect 2164 4613 2189 4616
rect 2226 4613 2260 4616
rect 2322 4613 2348 4616
rect 2378 4613 2404 4616
rect 2540 4613 2565 4616
rect 2692 4613 2709 4616
rect 2850 4613 2876 4616
rect 866 4603 940 4606
rect 1092 4603 1101 4606
rect 1130 4603 1156 4606
rect 1514 4605 1517 4613
rect 2898 4606 2901 4623
rect 2948 4613 2957 4616
rect 3284 4613 3309 4616
rect 3442 4613 3452 4616
rect 3498 4613 3508 4616
rect 3660 4613 3669 4616
rect 3748 4613 3773 4616
rect 3804 4613 3813 4616
rect 3940 4613 3957 4616
rect 3996 4613 4021 4616
rect 4052 4613 4061 4616
rect 4100 4613 4125 4616
rect 4156 4613 4165 4616
rect 4244 4613 4261 4616
rect 4364 4613 4389 4616
rect 4420 4613 4437 4616
rect 4596 4613 4605 4616
rect 1898 4603 1908 4606
rect 2234 4603 2252 4606
rect 2298 4603 2308 4606
rect 2810 4603 2828 4606
rect 2898 4603 2932 4606
rect 2956 4603 3045 4606
rect 3306 4605 3309 4613
rect 3666 4605 3669 4613
rect 3810 4605 3813 4613
rect 4162 4605 4165 4613
rect 4434 4605 4437 4613
rect 4450 4603 4476 4606
rect 4508 4603 4525 4606
rect 38 4567 4829 4573
rect 866 4543 932 4546
rect 2714 4543 2788 4546
rect 2802 4543 2836 4546
rect 156 4533 197 4536
rect 234 4533 260 4536
rect 276 4533 309 4536
rect 324 4533 349 4536
rect 372 4533 396 4536
rect 412 4533 485 4536
rect 548 4533 565 4536
rect 818 4533 836 4536
rect 852 4533 861 4536
rect 898 4533 940 4536
rect 980 4533 989 4536
rect 1106 4533 1116 4536
rect 1132 4533 1165 4536
rect 1170 4533 1180 4536
rect 1210 4533 1236 4536
rect 1260 4533 1269 4536
rect 1300 4533 1309 4536
rect 1340 4533 1357 4536
rect 1372 4533 1381 4536
rect 1420 4533 1429 4536
rect 1434 4533 1492 4536
rect 1524 4533 1589 4536
rect 1628 4533 1653 4536
rect 1658 4533 1668 4536
rect 1690 4533 1724 4536
rect 1850 4533 1884 4536
rect 1900 4533 1909 4536
rect 1924 4533 1973 4536
rect 2034 4533 2060 4536
rect 2122 4533 2132 4536
rect 2164 4533 2220 4536
rect 2236 4533 2292 4536
rect 2308 4533 2325 4536
rect 2330 4533 2356 4536
rect 2394 4533 2444 4536
rect 2522 4533 2532 4536
rect 2548 4533 2661 4536
rect 2700 4533 2781 4536
rect 2796 4533 2829 4536
rect 2858 4533 2900 4536
rect 2930 4533 2940 4536
rect 2970 4533 2980 4536
rect 3004 4533 3021 4536
rect 3076 4533 3093 4536
rect 3108 4533 3141 4536
rect 3146 4533 3188 4536
rect 3220 4533 3268 4536
rect 3300 4533 3309 4536
rect 3458 4533 3484 4536
rect 3516 4533 3541 4536
rect 3546 4533 3556 4536
rect 3618 4533 3636 4536
rect 3658 4533 3708 4536
rect 3724 4533 3773 4536
rect 3812 4533 3852 4536
rect 3916 4533 3949 4536
rect 4108 4533 4141 4536
rect 4180 4533 4197 4536
rect 4202 4533 4244 4536
rect 4292 4533 4301 4536
rect 4306 4533 4340 4536
rect 4356 4533 4381 4536
rect 4394 4533 4404 4536
rect 4306 4526 4309 4533
rect 4570 4526 4573 4535
rect 164 4523 204 4526
rect 236 4523 245 4526
rect 306 4523 316 4526
rect 322 4523 348 4526
rect 500 4523 517 4526
rect 556 4523 565 4526
rect 618 4523 684 4526
rect 1044 4523 1053 4526
rect 1146 4523 1188 4526
rect 1346 4523 1364 4526
rect 1412 4523 1461 4526
rect 1626 4523 1676 4526
rect 1682 4523 1732 4526
rect 1788 4523 1813 4526
rect 1844 4523 1869 4526
rect 1930 4523 1972 4526
rect 2004 4523 2052 4526
rect 2178 4523 2212 4526
rect 2274 4523 2284 4526
rect 2322 4523 2364 4526
rect 2394 4523 2452 4526
rect 2482 4523 2524 4526
rect 2570 4523 2676 4526
rect 2708 4523 2741 4526
rect 2804 4523 2837 4526
rect 2874 4523 2908 4526
rect 2956 4523 2981 4526
rect 3042 4523 3052 4526
rect 3082 4523 3100 4526
rect 3146 4523 3196 4526
rect 3314 4523 3324 4526
rect 3452 4523 3485 4526
rect 3522 4523 3564 4526
rect 3660 4523 3693 4526
rect 3732 4523 3757 4526
rect 3930 4523 3964 4526
rect 4042 4523 4068 4526
rect 4082 4523 4100 4526
rect 4284 4523 4309 4526
rect 4364 4523 4397 4526
rect 4564 4523 4573 4526
rect 4626 4523 4660 4526
rect 980 4513 1005 4516
rect 1204 4513 1229 4516
rect 1266 4513 1276 4516
rect 1306 4513 1316 4516
rect 2924 4513 2933 4516
rect 2970 4513 2973 4523
rect 3364 4513 3373 4516
rect 3404 4513 3437 4516
rect 3388 4503 3397 4506
rect 14 4467 4853 4473
rect 1196 4423 1205 4426
rect 2908 4423 2917 4426
rect 2946 4423 2956 4426
rect 3402 4423 3412 4426
rect 3436 4423 3445 4426
rect 172 4413 197 4416
rect 300 4413 309 4416
rect 498 4413 508 4416
rect 538 4413 548 4416
rect 578 4406 581 4414
rect 586 4413 628 4416
rect 658 4413 692 4416
rect 748 4413 757 4416
rect 860 4413 869 4416
rect 916 4413 933 4416
rect 972 4413 989 4416
rect 1020 4413 1045 4416
rect 1058 4413 1084 4416
rect 1116 4413 1133 4416
rect 1202 4406 1205 4423
rect 1324 4413 1333 4416
rect 1458 4413 1508 4416
rect 1514 4413 1524 4416
rect 1724 4413 1749 4416
rect 1786 4413 1796 4416
rect 1802 4413 1844 4416
rect 1876 4413 1885 4416
rect 1954 4413 1972 4416
rect 2010 4413 2028 4416
rect 2066 4413 2100 4416
rect 2132 4413 2141 4416
rect 2172 4413 2181 4416
rect 2218 4413 2244 4416
rect 2356 4413 2381 4416
rect 2500 4413 2509 4416
rect 2564 4413 2581 4416
rect 2690 4413 2700 4416
rect 2732 4413 2741 4416
rect 2874 4413 2885 4416
rect 2978 4413 2989 4416
rect 3106 4413 3132 4416
rect 3308 4413 3333 4416
rect 3748 4413 3773 4416
rect 3804 4413 3829 4416
rect 3938 4413 3988 4416
rect 4196 4413 4213 4416
rect 4324 4413 4341 4416
rect 4380 4413 4389 4416
rect 4458 4413 4492 4416
rect 4620 4413 4629 4416
rect 4642 4413 4652 4416
rect 178 4403 204 4406
rect 516 4403 549 4406
rect 578 4403 605 4406
rect 610 4403 620 4406
rect 674 4403 684 4406
rect 754 4403 772 4406
rect 788 4403 813 4406
rect 964 4403 973 4406
rect 986 4403 1012 4406
rect 1060 4403 1085 4406
rect 1202 4403 1236 4406
rect 1260 4403 1301 4406
rect 1332 4403 1357 4406
rect 1474 4403 1500 4406
rect 1804 4403 1845 4406
rect 1868 4403 1908 4406
rect 1940 4403 1965 4406
rect 2090 4403 2108 4406
rect 2130 4403 2164 4406
rect 2282 4403 2292 4406
rect 2314 4403 2348 4406
rect 2508 4403 2524 4406
rect 2546 4403 2556 4406
rect 2682 4403 2708 4406
rect 2730 4403 2740 4406
rect 2874 4405 2877 4413
rect 2908 4403 2917 4406
rect 2932 4403 2941 4406
rect 2946 4403 2956 4406
rect 2986 4405 2989 4413
rect 3012 4403 3021 4406
rect 3826 4405 3829 4413
rect 3916 4403 3933 4406
rect 3946 4403 3980 4406
rect 4386 4405 4389 4413
rect 4436 4403 4477 4406
rect 4626 4405 4629 4413
rect 922 4393 956 4396
rect 978 4393 1004 4396
rect 1122 4393 1148 4396
rect 38 4367 4829 4373
rect 1018 4343 1060 4346
rect 2810 4343 2828 4346
rect 2898 4343 2908 4346
rect 2930 4343 2956 4346
rect 2970 4343 2997 4346
rect 2970 4336 2973 4343
rect 162 4333 204 4336
rect 236 4333 245 4336
rect 258 4333 268 4336
rect 324 4333 349 4336
rect 516 4333 549 4336
rect 610 4333 628 4336
rect 650 4333 660 4336
rect 810 4333 820 4336
rect 884 4333 909 4336
rect 932 4333 988 4336
rect 1068 4333 1085 4336
rect 1106 4333 1132 4336
rect 1162 4333 1204 4336
rect 1228 4333 1261 4336
rect 1362 4333 1396 4336
rect 1458 4333 1476 4336
rect 1508 4333 1541 4336
rect 1812 4333 1845 4336
rect 1868 4333 1916 4336
rect 1948 4333 1957 4336
rect 1988 4333 1997 4336
rect 2028 4333 2077 4336
rect 2098 4333 2108 4336
rect 2300 4333 2317 4336
rect 2378 4333 2388 4336
rect 2554 4333 2580 4336
rect 162 4323 165 4333
rect 250 4323 276 4326
rect 306 4323 316 4326
rect 322 4323 348 4326
rect 436 4323 461 4326
rect 498 4323 508 4326
rect 514 4323 548 4326
rect 580 4323 620 4326
rect 668 4323 701 4326
rect 802 4323 828 4326
rect 866 4323 876 4326
rect 882 4323 908 4326
rect 1076 4323 1125 4326
rect 1130 4323 1140 4326
rect 1162 4316 1165 4333
rect 1220 4323 1253 4326
rect 1300 4323 1325 4326
rect 1356 4323 1365 4326
rect 1370 4323 1469 4326
rect 1500 4323 1509 4326
rect 1578 4323 1604 4326
rect 1642 4323 1668 4326
rect 1674 4323 1692 4326
rect 1740 4323 1765 4326
rect 1810 4323 1844 4326
rect 1876 4323 1885 4326
rect 1914 4323 1924 4326
rect 1980 4323 1989 4326
rect 1994 4323 2004 4326
rect 2050 4323 2084 4326
rect 2116 4323 2149 4326
rect 2196 4323 2221 4326
rect 2258 4323 2292 4326
rect 2306 4323 2316 4326
rect 2348 4323 2389 4326
rect 2434 4323 2460 4326
rect 2546 4323 2572 4326
rect 2602 4325 2605 4336
rect 2626 4333 2644 4336
rect 2666 4333 2684 4336
rect 2850 4333 2868 4336
rect 2892 4333 2909 4336
rect 2916 4333 2957 4336
rect 2964 4333 2973 4336
rect 2978 4333 3004 4336
rect 3028 4333 3069 4336
rect 3114 4333 3172 4336
rect 3220 4333 3261 4336
rect 3458 4333 3492 4336
rect 3564 4333 3604 4336
rect 3676 4333 3685 4336
rect 3698 4333 3724 4336
rect 3746 4333 3788 4336
rect 3820 4333 3861 4336
rect 4026 4333 4052 4336
rect 4178 4333 4196 4336
rect 4266 4333 4276 4336
rect 4314 4333 4324 4336
rect 4356 4333 4365 4336
rect 4396 4333 4421 4336
rect 3698 4326 3701 4333
rect 4442 4326 4445 4336
rect 4468 4333 4509 4336
rect 4770 4333 4780 4336
rect 2610 4323 2636 4326
rect 2668 4323 2677 4326
rect 2692 4323 2709 4326
rect 2866 4323 2876 4326
rect 3234 4323 3268 4326
rect 3364 4323 3413 4326
rect 3444 4323 3493 4326
rect 3500 4323 3525 4326
rect 3556 4323 3565 4326
rect 3570 4323 3612 4326
rect 3642 4323 3701 4326
rect 3706 4323 3716 4326
rect 3748 4323 3789 4326
rect 3946 4323 3972 4326
rect 4026 4323 4060 4326
rect 4164 4323 4173 4326
rect 4178 4323 4204 4326
rect 4234 4323 4244 4326
rect 4250 4323 4284 4326
rect 4322 4323 4332 4326
rect 4362 4323 4372 4326
rect 4404 4325 4445 4326
rect 4404 4323 4444 4325
rect 4778 4323 4788 4326
rect 1012 4313 1053 4316
rect 1156 4313 1165 4316
rect 1194 4313 1204 4316
rect 1994 4313 1997 4323
rect 2892 4313 2901 4316
rect 2986 4313 3004 4316
rect 14 4267 4853 4273
rect 3404 4233 3413 4236
rect 4300 4233 4309 4236
rect 1194 4223 1260 4226
rect 1290 4223 1332 4226
rect 2852 4223 2869 4226
rect 2970 4223 2980 4226
rect 3386 4223 3396 4226
rect 3420 4223 3461 4226
rect 4282 4223 4292 4226
rect 4306 4223 4316 4226
rect 108 4213 117 4216
rect 242 4213 252 4216
rect 388 4213 397 4216
rect 444 4213 501 4216
rect 506 4213 532 4216
rect 564 4213 573 4216
rect 596 4213 613 4216
rect 732 4213 749 4216
rect 860 4213 869 4216
rect 916 4213 949 4216
rect 964 4213 1005 4216
rect 506 4206 509 4213
rect 1034 4206 1037 4214
rect 1106 4213 1116 4216
rect 1188 4213 1253 4216
rect 1276 4213 1333 4216
rect 1354 4213 1372 4216
rect 1420 4213 1429 4216
rect 1514 4213 1548 4216
rect 1562 4213 1588 4216
rect 1642 4213 1668 4216
rect 1764 4213 1789 4216
rect 1866 4213 1892 4216
rect 1906 4213 1932 4216
rect 1938 4213 1972 4216
rect 2002 4213 2028 4216
rect 2082 4213 2100 4216
rect 2146 4213 2156 4216
rect 2220 4213 2245 4216
rect 2602 4213 2620 4216
rect 2652 4213 2677 4216
rect 2692 4213 2709 4216
rect 2804 4213 2813 4216
rect 2818 4213 2836 4216
rect 2946 4213 2981 4216
rect 3082 4213 3092 4216
rect 3098 4213 3108 4216
rect 3146 4213 3164 4216
rect 3202 4213 3212 4216
rect 3252 4213 3261 4216
rect 3274 4213 3284 4216
rect 3314 4213 3340 4216
rect 3500 4213 3540 4216
rect 3578 4213 3612 4216
rect 3642 4213 3676 4216
rect 3682 4213 3692 4216
rect 3722 4213 3748 4216
rect 3786 4213 3804 4216
rect 3890 4213 3916 4216
rect 3930 4213 3972 4216
rect 4028 4213 4053 4216
rect 4090 4213 4100 4216
rect 4130 4213 4205 4216
rect 4210 4213 4228 4216
rect 4436 4213 4445 4216
rect 4468 4213 4492 4216
rect 2082 4206 2085 4213
rect 2810 4206 2813 4213
rect 458 4203 509 4206
rect 522 4203 540 4206
rect 562 4203 588 4206
rect 746 4203 764 4206
rect 956 4203 1005 4206
rect 1034 4203 1060 4206
rect 1084 4203 1093 4206
rect 1114 4203 1124 4206
rect 1146 4203 1180 4206
rect 1194 4203 1260 4206
rect 1284 4203 1325 4206
rect 1444 4203 1453 4206
rect 1458 4203 1484 4206
rect 1516 4203 1541 4206
rect 1570 4203 1580 4206
rect 1826 4203 1836 4206
rect 1954 4203 1964 4206
rect 1996 4203 2029 4206
rect 2052 4203 2085 4206
rect 2202 4203 2212 4206
rect 2410 4203 2444 4206
rect 2650 4203 2684 4206
rect 2810 4203 2828 4206
rect 2852 4203 2869 4206
rect 2898 4203 2924 4206
rect 2946 4205 2949 4213
rect 2954 4203 2980 4206
rect 3004 4203 3029 4206
rect 3068 4203 3085 4206
rect 3098 4205 3101 4213
rect 3218 4203 3228 4206
rect 3260 4203 3277 4206
rect 3434 4203 3476 4206
rect 3492 4203 3501 4206
rect 3522 4203 3548 4206
rect 3564 4203 3597 4206
rect 3636 4203 3653 4206
rect 3682 4205 3685 4213
rect 4202 4206 4205 4213
rect 3828 4203 3853 4206
rect 3980 4203 3989 4206
rect 4202 4203 4236 4206
rect 4252 4203 4277 4206
rect 4442 4205 4445 4213
rect 4562 4206 4565 4214
rect 4602 4213 4676 4216
rect 4706 4213 4740 4216
rect 4522 4203 4540 4206
rect 4562 4203 4573 4206
rect 4588 4203 4653 4206
rect 4658 4203 4668 4206
rect 4700 4203 4732 4206
rect 922 4193 948 4196
rect 962 4193 1020 4196
rect 2858 4193 2876 4196
rect 38 4167 4829 4173
rect 1122 4143 1156 4146
rect 132 4133 157 4136
rect 162 4133 172 4136
rect 188 4133 197 4136
rect 340 4133 349 4136
rect 436 4133 469 4136
rect 492 4133 501 4136
rect 506 4133 540 4136
rect 562 4133 588 4136
rect 892 4133 941 4136
rect 978 4133 1012 4136
rect 1036 4133 1045 4136
rect 1050 4133 1092 4136
rect 1116 4133 1157 4136
rect 1298 4133 1340 4136
rect 1364 4133 1389 4136
rect 1428 4133 1437 4136
rect 1562 4133 1604 4136
rect 1700 4133 1709 4136
rect 1810 4133 1868 4136
rect 1882 4133 1924 4136
rect 1956 4133 1997 4136
rect 2138 4133 2172 4136
rect 2202 4133 2244 4136
rect 2362 4133 2396 4136
rect 2556 4133 2597 4136
rect 2626 4133 2668 4136
rect 2690 4133 2708 4136
rect 2842 4133 2868 4136
rect 2898 4133 2948 4136
rect 2972 4133 3021 4136
rect 3036 4133 3101 4136
rect 3114 4133 3140 4136
rect 3172 4133 3205 4136
rect 1994 4126 1997 4133
rect 114 4123 124 4126
rect 202 4123 220 4126
rect 268 4123 293 4126
rect 394 4123 428 4126
rect 458 4123 468 4126
rect 596 4123 637 4126
rect 674 4123 700 4126
rect 770 4123 796 4126
rect 866 4123 884 4126
rect 890 4123 940 4126
rect 972 4123 1013 4126
rect 1186 4123 1204 4126
rect 1250 4123 1260 4126
rect 1420 4123 1445 4126
rect 1450 4123 1460 4126
rect 1498 4123 1516 4126
rect 1666 4123 1757 4126
rect 1796 4123 1861 4126
rect 1866 4123 1876 4126
rect 1914 4123 1932 4126
rect 1994 4123 2028 4126
rect 2122 4123 2164 4126
rect 2196 4123 2213 4126
rect 2290 4123 2316 4126
rect 2420 4123 2445 4126
rect 2554 4123 2596 4126
rect 2628 4123 2653 4126
rect 2692 4123 2701 4126
rect 2844 4123 2861 4126
rect 2866 4123 2876 4126
rect 2898 4116 2901 4133
rect 3338 4126 3341 4135
rect 3354 4133 3364 4136
rect 3530 4133 3556 4136
rect 3730 4126 3733 4135
rect 3850 4133 3876 4136
rect 3908 4133 3933 4136
rect 4130 4133 4164 4136
rect 4458 4126 4461 4135
rect 4554 4133 4564 4136
rect 4580 4133 4605 4136
rect 4602 4126 4605 4133
rect 2978 4123 3028 4126
rect 3042 4123 3148 4126
rect 3300 4123 3341 4126
rect 3380 4123 3397 4126
rect 3700 4123 3733 4126
rect 3746 4123 3756 4126
rect 3802 4123 3828 4126
rect 3874 4123 3884 4126
rect 4130 4123 4205 4126
rect 4436 4123 4461 4126
rect 4530 4123 4556 4126
rect 4602 4123 4637 4126
rect 4644 4123 4653 4126
rect 1036 4113 1077 4116
rect 1116 4113 1149 4116
rect 1314 4113 1340 4116
rect 2892 4113 2901 4116
rect 2922 4113 2948 4116
rect 3436 4113 3445 4116
rect 4482 4113 4492 4116
rect 14 4067 4853 4073
rect 2852 4023 2885 4026
rect 2916 4023 2925 4026
rect 108 4013 133 4016
rect 194 4013 204 4016
rect 242 4013 276 4016
rect 306 4013 332 4016
rect 412 4013 437 4016
rect 498 4013 516 4016
rect 562 4013 596 4016
rect 642 4013 660 4016
rect 706 4013 716 4016
rect 908 4013 933 4016
rect 964 4013 981 4016
rect 1020 4013 1045 4016
rect 1050 4013 1060 4016
rect 1098 4013 1132 4016
rect 1258 4013 1284 4016
rect 1396 4013 1421 4016
rect 1610 4013 1628 4016
rect 1716 4013 1741 4016
rect 1778 4013 1796 4016
rect 1802 4013 1812 4016
rect 1826 4013 1884 4016
rect 1954 4013 2004 4016
rect 2042 4013 2068 4016
rect 2106 4013 2132 4016
rect 2146 4013 2172 4016
rect 2204 4013 2213 4016
rect 2218 4013 2284 4016
rect 2330 4013 2348 4016
rect 2394 4013 2412 4016
rect 2506 4013 2532 4016
rect 2588 4013 2605 4016
rect 2642 4013 2668 4016
rect 2818 4013 2836 4016
rect 2850 4013 2900 4016
rect 642 4006 645 4013
rect 2922 4006 2925 4023
rect 2956 4013 2965 4016
rect 3044 4013 3053 4016
rect 3292 4013 3325 4016
rect 3458 4013 3500 4016
rect 3602 4013 3644 4016
rect 3682 4013 3700 4016
rect 3738 4013 3772 4016
rect 3916 4013 3941 4016
rect 3972 4013 3981 4016
rect 3988 4013 4029 4016
rect 4068 4013 4093 4016
rect 4124 4013 4173 4016
rect 4258 4013 4292 4016
rect 4436 4013 4461 4016
rect 4474 4013 4500 4016
rect 4620 4013 4669 4016
rect 4676 4013 4685 4016
rect 180 4003 205 4006
rect 300 4003 340 4006
rect 484 4003 517 4006
rect 540 4003 557 4006
rect 594 4003 604 4006
rect 620 4003 645 4006
rect 1012 4003 1021 4006
rect 1026 4003 1068 4006
rect 1084 4003 1140 4006
rect 1162 4003 1212 4006
rect 1458 4003 1484 4006
rect 1522 4003 1564 4006
rect 1636 4003 1645 4006
rect 1834 4003 1876 4006
rect 1956 4003 1997 4006
rect 2026 4003 2076 4006
rect 2098 4003 2124 4006
rect 2138 4003 2180 4006
rect 2196 4003 2261 4006
rect 2300 4003 2317 4006
rect 2346 4003 2356 4006
rect 2372 4003 2405 4006
rect 2434 4003 2460 4006
rect 2852 4003 2861 4006
rect 2922 4003 2940 4006
rect 2964 4003 3005 4006
rect 3322 4005 3325 4013
rect 3394 4003 3412 4006
rect 3516 4003 3549 4006
rect 3826 4003 3861 4006
rect 3978 4005 3981 4013
rect 4202 4003 4220 4006
rect 4236 4003 4253 4006
rect 4266 4003 4284 4006
rect 4316 4003 4325 4006
rect 4458 4005 4461 4013
rect 4666 4005 4669 4013
rect 978 3993 1004 3996
rect 38 3967 4829 3973
rect 1114 3953 1173 3956
rect 946 3943 972 3946
rect 2818 3943 2852 3946
rect 2866 3943 2892 3946
rect 180 3933 205 3936
rect 258 3926 261 3936
rect 290 3933 324 3936
rect 484 3933 533 3936
rect 586 3933 612 3936
rect 666 3933 684 3936
rect 748 3933 773 3936
rect 796 3933 845 3936
rect 1020 3933 1029 3936
rect 1250 3933 1292 3936
rect 1316 3933 1349 3936
rect 1450 3933 1460 3936
rect 108 3923 133 3926
rect 194 3923 204 3926
rect 236 3925 261 3926
rect 236 3923 260 3925
rect 292 3923 309 3926
rect 332 3923 365 3926
rect 402 3923 428 3926
rect 466 3923 476 3926
rect 498 3923 532 3926
rect 636 3923 645 3926
rect 692 3923 701 3926
rect 740 3923 765 3926
rect 804 3923 821 3926
rect 884 3923 893 3926
rect 940 3923 957 3926
rect 988 3923 997 3926
rect 1034 3923 1068 3926
rect 1218 3923 1228 3926
rect 1250 3916 1253 3933
rect 1490 3926 1493 3936
rect 1522 3926 1525 3935
rect 1722 3933 1748 3936
rect 1780 3933 1829 3936
rect 2026 3933 2052 3936
rect 2068 3933 2077 3936
rect 2106 3933 2132 3936
rect 2186 3933 2228 3936
rect 2290 3933 2348 3936
rect 2364 3933 2381 3936
rect 2394 3933 2428 3936
rect 2596 3933 2613 3936
rect 2626 3933 2652 3936
rect 2674 3933 2692 3936
rect 2812 3933 2821 3936
rect 2860 3933 2893 3936
rect 2906 3933 2940 3936
rect 2964 3933 3005 3936
rect 2026 3926 2029 3933
rect 2186 3926 2189 3933
rect 3106 3926 3109 3935
rect 3130 3933 3140 3936
rect 3178 3933 3220 3936
rect 3252 3933 3261 3936
rect 3362 3926 3365 3935
rect 3474 3933 3492 3936
rect 3508 3933 3549 3936
rect 4034 3933 4044 3936
rect 4148 3933 4165 3936
rect 4194 3933 4228 3936
rect 4244 3933 4285 3936
rect 4530 3933 4556 3936
rect 4588 3933 4613 3936
rect 4626 3933 4636 3936
rect 3546 3926 3549 3933
rect 4194 3926 4197 3933
rect 1308 3923 1317 3926
rect 1388 3923 1413 3926
rect 1458 3923 1493 3926
rect 1498 3923 1516 3926
rect 1522 3923 1572 3926
rect 1610 3923 1628 3926
rect 1698 3923 1756 3926
rect 1762 3923 1772 3926
rect 1802 3923 1828 3926
rect 1940 3923 1949 3926
rect 1996 3923 2029 3926
rect 2076 3923 2085 3926
rect 2148 3923 2189 3926
rect 2322 3923 2340 3926
rect 2436 3923 2445 3926
rect 2498 3923 2508 3926
rect 2554 3923 2572 3926
rect 2604 3923 2613 3926
rect 2618 3923 2644 3926
rect 2700 3923 2757 3926
rect 2770 3923 2796 3926
rect 2868 3923 2885 3926
rect 2908 3923 2917 3926
rect 3044 3923 3069 3926
rect 3100 3923 3109 3926
rect 3116 3923 3125 3926
rect 3300 3923 3325 3926
rect 3356 3923 3365 3926
rect 3372 3923 3397 3926
rect 3546 3923 3564 3926
rect 3852 3923 3885 3926
rect 4026 3923 4052 3926
rect 4090 3923 4124 3926
rect 4154 3923 4197 3926
rect 4210 3923 4220 3926
rect 4258 3923 4300 3926
rect 4372 3923 4397 3926
rect 4428 3923 4453 3926
rect 4602 3923 4628 3926
rect 4658 3925 4661 3936
rect 4668 3923 4677 3926
rect 1020 3913 1061 3916
rect 1244 3913 1253 3916
rect 1282 3913 1292 3916
rect 2812 3913 2829 3916
rect 2922 3913 2940 3916
rect 3428 3913 3477 3916
rect 4524 3913 4533 3916
rect 14 3867 4853 3873
rect 3642 3843 3661 3846
rect 996 3823 1029 3826
rect 1322 3823 1340 3826
rect 2884 3823 2893 3826
rect 2922 3823 2932 3826
rect 4010 3823 4028 3826
rect 4052 3823 4077 3826
rect 148 3813 213 3816
rect 306 3813 340 3816
rect 428 3813 437 3816
rect 484 3813 541 3816
rect 546 3813 588 3816
rect 642 3813 668 3816
rect 698 3813 724 3816
rect 762 3813 796 3816
rect 826 3813 844 3816
rect 890 3813 900 3816
rect 938 3813 980 3816
rect 1068 3813 1093 3816
rect 1228 3813 1245 3816
rect 1314 3813 1341 3816
rect 1378 3813 1404 3816
rect 1410 3813 1485 3816
rect 1636 3813 1661 3816
rect 1716 3813 1733 3816
rect 1772 3813 1797 3816
rect 1842 3813 1884 3816
rect 2084 3813 2093 3816
rect 2132 3813 2157 3816
rect 2196 3813 2205 3816
rect 2276 3813 2285 3816
rect 2370 3813 2396 3816
rect 2442 3813 2452 3816
rect 2490 3813 2524 3816
rect 2556 3813 2565 3816
rect 2596 3813 2645 3816
rect 2812 3813 2821 3816
rect 2850 3813 2868 3816
rect 642 3806 645 3813
rect 116 3803 141 3806
rect 156 3803 173 3806
rect 218 3803 228 3806
rect 322 3803 332 3806
rect 364 3803 373 3806
rect 612 3803 645 3806
rect 778 3803 788 3806
rect 820 3803 845 3806
rect 868 3803 893 3806
rect 954 3803 972 3806
rect 996 3803 1013 3806
rect 1140 3803 1149 3806
rect 1194 3803 1212 3806
rect 1236 3803 1253 3806
rect 1258 3803 1284 3806
rect 1308 3803 1333 3806
rect 1338 3805 1341 3813
rect 1370 3803 1396 3806
rect 1466 3803 1492 3806
rect 1524 3803 1533 3806
rect 1658 3805 1661 3813
rect 2890 3806 2893 3823
rect 3012 3813 3037 3816
rect 3068 3813 3077 3816
rect 3148 3813 3165 3816
rect 3284 3813 3309 3816
rect 3380 3813 3397 3816
rect 3436 3813 3453 3816
rect 3506 3813 3540 3816
rect 3562 3813 3612 3816
rect 3700 3813 3725 3816
rect 3770 3813 3796 3816
rect 3834 3813 3876 3816
rect 3906 3813 3972 3816
rect 1948 3803 1989 3806
rect 2204 3803 2229 3806
rect 2284 3803 2381 3806
rect 2506 3803 2532 3806
rect 2554 3803 2588 3806
rect 2810 3803 2860 3806
rect 2890 3803 2932 3806
rect 2956 3803 2973 3806
rect 3074 3805 3077 3813
rect 3098 3803 3124 3806
rect 3156 3803 3189 3806
rect 3306 3805 3309 3813
rect 3490 3803 3532 3806
rect 3620 3803 3661 3806
rect 3820 3803 3861 3806
rect 3980 3803 4021 3806
rect 4042 3803 4045 3814
rect 4058 3813 4092 3816
rect 4188 3813 4213 3816
rect 4308 3813 4317 3816
rect 4354 3813 4388 3816
rect 4434 3813 4533 3816
rect 4636 3813 4645 3816
rect 4122 3803 4164 3806
rect 4314 3805 4317 3813
rect 4330 3803 4380 3806
rect 4450 3803 4468 3806
rect 4642 3805 4645 3813
rect 2746 3793 2796 3796
rect 38 3767 4829 3773
rect 962 3743 996 3746
rect 1026 3743 1060 3746
rect 2818 3743 2828 3746
rect 290 3733 300 3736
rect 476 3733 509 3736
rect 532 3733 597 3736
rect 1068 3733 1077 3736
rect 1154 3733 1204 3736
rect 1228 3733 1253 3736
rect 1258 3733 1276 3736
rect 164 3723 173 3726
rect 268 3723 285 3726
rect 388 3723 413 3726
rect 458 3723 468 3726
rect 498 3723 508 3726
rect 540 3723 549 3726
rect 764 3723 773 3726
rect 1076 3723 1093 3726
rect 1106 3723 1132 3726
rect 1154 3716 1157 3733
rect 1258 3726 1261 3733
rect 1290 3726 1293 3735
rect 1500 3733 1533 3736
rect 1572 3733 1613 3736
rect 1932 3733 1965 3736
rect 1980 3733 1997 3736
rect 2020 3733 2037 3736
rect 2066 3733 2076 3736
rect 2034 3726 2037 3733
rect 1220 3723 1261 3726
rect 1284 3723 1293 3726
rect 1492 3723 1517 3726
rect 1636 3723 1653 3726
rect 1716 3723 1733 3726
rect 1906 3723 1924 3726
rect 1972 3723 1989 3726
rect 2034 3723 2068 3726
rect 2098 3725 2101 3736
rect 2130 3733 2140 3736
rect 2244 3733 2300 3736
rect 2332 3733 2372 3736
rect 2402 3733 2428 3736
rect 2524 3733 2597 3736
rect 2602 3733 2612 3736
rect 2628 3733 2645 3736
rect 2668 3733 2677 3736
rect 2682 3733 2692 3736
rect 2842 3733 2885 3736
rect 2916 3733 2940 3736
rect 2954 3733 3004 3736
rect 3028 3733 3077 3736
rect 3082 3733 3100 3736
rect 2106 3723 2148 3726
rect 2210 3723 2220 3726
rect 2282 3723 2308 3726
rect 2338 3723 2364 3726
rect 2396 3723 2429 3726
rect 2436 3723 2445 3726
rect 2458 3723 2500 3726
rect 2532 3723 2565 3726
rect 2586 3723 2604 3726
rect 2700 3723 2717 3726
rect 2754 3723 2780 3726
rect 2842 3725 2845 3733
rect 3274 3726 3277 3735
rect 3474 3733 3500 3736
rect 3516 3733 3565 3736
rect 3604 3733 3621 3736
rect 3676 3733 3717 3736
rect 4082 3726 4085 3735
rect 2908 3723 2925 3726
rect 2948 3723 3005 3726
rect 3124 3723 3149 3726
rect 3252 3723 3277 3726
rect 3340 3723 3365 3726
rect 3410 3723 3492 3726
rect 3554 3723 3580 3726
rect 3610 3723 3668 3726
rect 3732 3723 3781 3726
rect 3812 3723 3837 3726
rect 3996 3723 4021 3726
rect 4052 3723 4085 3726
rect 4092 3723 4117 3726
rect 4154 3723 4188 3726
rect 4218 3725 4221 3736
rect 4226 3733 4268 3736
rect 4300 3733 4317 3736
rect 4332 3733 4365 3736
rect 4524 3733 4533 3736
rect 4634 3733 4668 3736
rect 4740 3733 4757 3736
rect 4772 3733 4781 3736
rect 4258 3723 4276 3726
rect 4306 3723 4324 3726
rect 4474 3723 4499 3726
rect 4628 3723 4637 3726
rect 4650 3723 4676 3726
rect 4706 3723 4732 3726
rect 4738 3723 4764 3726
rect 1148 3713 1157 3716
rect 1194 3713 1204 3716
rect 2866 3713 2900 3716
rect 2970 3713 3004 3716
rect 14 3667 4853 3673
rect 3252 3633 3261 3636
rect 978 3623 997 3626
rect 1044 3623 1069 3626
rect 1194 3623 1204 3626
rect 1242 3623 1276 3626
rect 1356 3623 1413 3626
rect 2724 3623 2733 3626
rect 3268 3623 3277 3626
rect 4170 3623 4188 3626
rect 4202 3623 4212 3626
rect 4610 3623 4629 3626
rect 116 3613 141 3616
rect 194 3613 212 3616
rect 244 3613 261 3616
rect 370 3613 404 3616
rect 436 3613 445 3616
rect 484 3613 509 3616
rect 586 3613 604 3616
rect 780 3613 829 3616
rect 842 3613 860 3616
rect 914 3613 932 3616
rect 1100 3613 1117 3616
rect 1220 3613 1277 3616
rect 1298 3613 1309 3616
rect 1314 3613 1348 3616
rect 1354 3613 1420 3616
rect 1458 3613 1476 3616
rect 1682 3613 1692 3616
rect 1820 3613 1829 3616
rect 1900 3613 1909 3616
rect 2140 3613 2157 3616
rect 2196 3613 2205 3616
rect 2250 3613 2284 3616
rect 2548 3613 2573 3616
rect 2612 3613 2621 3616
rect 2668 3613 2701 3616
rect 1306 3606 1309 3613
rect 188 3603 213 3606
rect 372 3603 405 3606
rect 556 3603 605 3606
rect 666 3603 700 3606
rect 746 3603 764 3606
rect 788 3603 805 3606
rect 844 3603 861 3606
rect 906 3603 940 3606
rect 956 3603 1020 3606
rect 1148 3603 1181 3606
rect 1194 3603 1204 3606
rect 1250 3603 1276 3606
rect 1306 3603 1340 3606
rect 1740 3603 1789 3606
rect 1962 3603 1972 3606
rect 2210 3603 2220 3606
rect 2364 3603 2381 3606
rect 2386 3603 2428 3606
rect 2514 3603 2540 3606
rect 2698 3605 2701 3613
rect 2770 3606 2773 3614
rect 2860 3613 2909 3616
rect 2988 3613 3013 3616
rect 3044 3613 3053 3616
rect 3116 3613 3149 3616
rect 3274 3613 3341 3616
rect 3388 3613 3421 3616
rect 3570 3613 3580 3616
rect 3746 3613 3780 3616
rect 3812 3613 3837 3616
rect 3890 3613 3924 3616
rect 4012 3613 4037 3616
rect 4068 3613 4101 3616
rect 4108 3613 4117 3616
rect 4258 3613 4268 3616
rect 4298 3613 4372 3616
rect 4418 3613 4444 3616
rect 4490 3613 4499 3616
rect 4530 3613 4564 3616
rect 4626 3613 4637 3616
rect 2724 3603 2733 3606
rect 2770 3603 2797 3606
rect 2810 3603 2844 3606
rect 2868 3603 2901 3606
rect 2906 3605 2909 3613
rect 3050 3605 3053 3613
rect 3066 3603 3092 3606
rect 3130 3603 3172 3606
rect 3204 3603 3237 3606
rect 3426 3603 3452 3606
rect 3484 3603 3572 3606
rect 3604 3603 3621 3606
rect 3810 3603 3860 3606
rect 3892 3603 3909 3606
rect 3932 3603 3949 3606
rect 4098 3605 4101 3613
rect 4626 3606 4629 3613
rect 4226 3603 4260 3606
rect 4292 3603 4317 3606
rect 4322 3603 4364 3606
rect 4396 3603 4437 3606
rect 4468 3603 4485 3606
rect 4508 3603 4541 3606
rect 4572 3603 4629 3606
rect 2746 3593 2756 3596
rect 38 3567 4829 3573
rect 180 3533 205 3536
rect 228 3533 268 3536
rect 306 3526 309 3556
rect 3458 3553 3525 3556
rect 690 3543 732 3546
rect 826 3543 876 3546
rect 1026 3543 1044 3546
rect 2642 3543 2676 3546
rect 2690 3543 2716 3546
rect 2834 3543 2868 3546
rect 444 3533 469 3536
rect 530 3533 548 3536
rect 618 3533 629 3536
rect 684 3533 725 3536
rect 730 3533 740 3536
rect 778 3533 788 3536
rect 850 3533 884 3536
rect 1052 3533 1069 3536
rect 626 3526 629 3533
rect 1218 3526 1221 3534
rect 1250 3533 1276 3536
rect 108 3523 133 3526
rect 194 3523 204 3526
rect 292 3523 309 3526
rect 356 3523 381 3526
rect 418 3523 436 3526
rect 442 3523 468 3526
rect 524 3523 549 3526
rect 626 3523 636 3526
rect 754 3523 796 3526
rect 948 3523 957 3526
rect 1004 3523 1013 3526
rect 1060 3523 1077 3526
rect 1180 3523 1221 3526
rect 1298 3526 1301 3536
rect 1338 3533 1380 3536
rect 1418 3533 1508 3536
rect 1540 3533 1549 3536
rect 1596 3533 1613 3536
rect 1626 3533 1636 3536
rect 1812 3533 1821 3536
rect 2090 3533 2156 3536
rect 2234 3533 2300 3536
rect 2332 3533 2349 3536
rect 2570 3533 2612 3536
rect 2628 3533 2677 3536
rect 2684 3533 2717 3536
rect 2738 3533 2772 3536
rect 2828 3533 2845 3536
rect 2876 3533 2885 3536
rect 2890 3533 2916 3536
rect 1418 3526 1421 3533
rect 1818 3526 1821 3533
rect 2338 3526 2341 3533
rect 2938 3526 2941 3534
rect 3052 3533 3069 3536
rect 3108 3533 3156 3536
rect 3258 3533 3284 3536
rect 3322 3533 3332 3536
rect 3066 3526 3069 3533
rect 3322 3526 3325 3533
rect 3410 3526 3413 3536
rect 3436 3533 3453 3536
rect 3458 3526 3461 3553
rect 3482 3533 3532 3536
rect 3690 3533 3708 3536
rect 3788 3533 3805 3536
rect 4066 3526 4069 3534
rect 4146 3533 4164 3536
rect 4186 3533 4228 3536
rect 4244 3533 4285 3536
rect 4450 3533 4468 3536
rect 4636 3533 4669 3536
rect 4770 3526 4773 3534
rect 1298 3523 1324 3526
rect 1404 3523 1421 3526
rect 1532 3523 1565 3526
rect 1700 3523 1725 3526
rect 1770 3523 1788 3526
rect 1818 3523 1828 3526
rect 1866 3523 1884 3526
rect 2036 3523 2045 3526
rect 2202 3523 2212 3526
rect 2274 3523 2308 3526
rect 2338 3523 2380 3526
rect 2474 3523 2492 3526
rect 2522 3523 2532 3526
rect 2562 3523 2604 3526
rect 2692 3523 2701 3526
rect 2794 3523 2812 3526
rect 2938 3523 3021 3526
rect 3066 3523 3084 3526
rect 3180 3523 3205 3526
rect 3308 3523 3325 3526
rect 3362 3525 3413 3526
rect 3362 3523 3412 3525
rect 3444 3523 3461 3526
rect 3556 3523 3573 3526
rect 3626 3523 3652 3526
rect 3754 3523 3764 3526
rect 4036 3523 4069 3526
rect 4194 3523 4220 3526
rect 4338 3523 4364 3526
rect 4458 3523 4476 3526
rect 4538 3523 4564 3526
rect 4764 3523 4773 3526
rect 1244 3513 1261 3516
rect 2828 3513 2837 3516
rect 2898 3513 2916 3516
rect 3194 3513 3212 3516
rect 3236 3513 3285 3516
rect 4082 3513 4116 3516
rect 4140 3513 4157 3516
rect 14 3467 4853 3473
rect 4074 3433 4093 3436
rect 4140 3433 4157 3436
rect 1308 3423 1317 3426
rect 2884 3423 2901 3426
rect 3538 3416 3541 3426
rect 4050 3423 4060 3426
rect 164 3413 189 3416
rect 226 3413 236 3416
rect 258 3413 268 3416
rect 300 3413 317 3416
rect 578 3413 612 3416
rect 1004 3413 1013 3416
rect 1258 3413 1292 3416
rect 1436 3413 1461 3416
rect 1540 3413 1565 3416
rect 1596 3413 1621 3416
rect 1684 3413 1693 3416
rect 1740 3413 1749 3416
rect 1770 3413 1820 3416
rect 1866 3413 1908 3416
rect 1914 3413 1948 3416
rect 1980 3413 2013 3416
rect 2034 3413 2076 3416
rect 2308 3413 2333 3416
rect 2364 3413 2373 3416
rect 2378 3413 2388 3416
rect 2444 3413 2453 3416
rect 2484 3413 2509 3416
rect 2548 3413 2565 3416
rect 2834 3413 2868 3416
rect 3124 3413 3149 3416
rect 3236 3413 3245 3416
rect 3404 3413 3429 3416
rect 3514 3413 3572 3416
rect 3682 3413 3796 3416
rect 3826 3413 3852 3416
rect 3988 3413 4013 3416
rect 4074 3415 4077 3433
rect 4090 3426 4093 3433
rect 4090 3423 4132 3426
rect 4156 3423 4197 3426
rect 4162 3413 4204 3416
rect 4282 3413 4300 3416
rect 4324 3413 4389 3416
rect 4402 3413 4412 3416
rect 4444 3413 4468 3416
rect 4490 3413 4500 3416
rect 4644 3413 4653 3416
rect 4674 3413 4764 3416
rect 244 3403 269 3406
rect 292 3403 325 3406
rect 458 3403 468 3406
rect 636 3403 645 3406
rect 666 3403 700 3406
rect 996 3403 1045 3406
rect 1250 3403 1284 3406
rect 1308 3403 1325 3406
rect 1444 3403 1493 3406
rect 1618 3405 1621 3413
rect 1916 3403 1949 3406
rect 1978 3403 2084 3406
rect 2540 3403 2565 3406
rect 2666 3403 2724 3406
rect 2842 3403 2860 3406
rect 2884 3403 2909 3406
rect 2916 3403 2973 3406
rect 3426 3405 3429 3413
rect 3580 3403 3597 3406
rect 3706 3403 3788 3406
rect 3860 3403 3893 3406
rect 4010 3405 4013 3413
rect 4228 3403 4293 3406
rect 4370 3403 4420 3406
rect 4524 3403 4533 3406
rect 4650 3405 4653 3413
rect 818 3393 988 3396
rect 2890 3393 2908 3396
rect 38 3367 4829 3373
rect 2802 3343 2828 3346
rect 4514 3336 4517 3346
rect 188 3333 205 3336
rect 218 3333 236 3336
rect 268 3333 308 3336
rect 324 3333 349 3336
rect 402 3333 452 3336
rect 468 3333 517 3336
rect 540 3333 573 3336
rect 682 3333 764 3336
rect 906 3333 916 3336
rect 946 3333 1084 3336
rect 1154 3333 1212 3336
rect 1308 3333 1317 3336
rect 116 3323 141 3326
rect 404 3323 437 3326
rect 482 3323 516 3326
rect 780 3323 797 3326
rect 844 3323 861 3326
rect 914 3323 924 3326
rect 1042 3323 1076 3326
rect 1154 3323 1157 3333
rect 1466 3326 1469 3335
rect 1674 3333 1716 3336
rect 1772 3333 1797 3336
rect 2290 3333 2316 3336
rect 2346 3333 2364 3336
rect 2506 3333 2532 3336
rect 2658 3333 2676 3336
rect 2842 3333 2940 3336
rect 2970 3333 2996 3336
rect 3020 3333 3053 3336
rect 3172 3333 3181 3336
rect 3210 3333 3220 3336
rect 3252 3333 3269 3336
rect 3428 3333 3477 3336
rect 3684 3333 3693 3336
rect 3730 3326 3733 3336
rect 3756 3333 3781 3336
rect 3970 3326 3973 3334
rect 4202 3326 4205 3334
rect 4378 3333 4388 3336
rect 4476 3333 4517 3336
rect 4642 3333 4661 3336
rect 4772 3333 4789 3336
rect 1186 3323 1213 3326
rect 1388 3323 1413 3326
rect 1444 3323 1469 3326
rect 1476 3323 1485 3326
rect 1660 3323 1685 3326
rect 1732 3323 1749 3326
rect 1812 3323 1829 3326
rect 1866 3323 1892 3326
rect 1980 3323 1989 3326
rect 2076 3323 2085 3326
rect 2172 3323 2189 3326
rect 2234 3323 2244 3326
rect 2340 3323 2357 3326
rect 2362 3323 2372 3326
rect 2386 3323 2412 3326
rect 2450 3323 2468 3326
rect 2540 3323 2557 3326
rect 2594 3323 2620 3326
rect 2844 3323 2909 3326
rect 2956 3323 2997 3326
rect 3034 3323 3060 3326
rect 3090 3323 3116 3326
rect 3154 3323 3164 3326
rect 3258 3323 3284 3326
rect 3378 3323 3404 3326
rect 3436 3323 3461 3326
rect 3508 3323 3525 3326
rect 3564 3323 3589 3326
rect 3620 3323 3629 3326
rect 3676 3323 3685 3326
rect 3690 3325 3733 3326
rect 3690 3323 3732 3325
rect 3764 3323 3781 3326
rect 3900 3323 3925 3326
rect 3956 3323 3973 3326
rect 4042 3323 4052 3326
rect 4132 3323 4157 3326
rect 4188 3323 4205 3326
rect 4434 3323 4452 3326
rect 4514 3323 4548 3326
rect 4578 3323 4612 3326
rect 4642 3325 4645 3333
rect 1308 3313 1325 3316
rect 2970 3313 2996 3316
rect 3356 3313 3397 3316
rect 14 3267 4853 3273
rect 2306 3243 2317 3246
rect 1108 3223 1133 3226
rect 1322 3223 1356 3226
rect 1394 3216 1397 3226
rect 1426 3223 1445 3226
rect 84 3213 117 3216
rect 220 3213 237 3216
rect 292 3213 317 3216
rect 354 3213 364 3216
rect 370 3213 404 3216
rect 436 3213 445 3216
rect 700 3213 725 3216
rect 730 3213 756 3216
rect 786 3206 789 3214
rect 802 3213 876 3216
rect 908 3213 917 3216
rect 988 3213 1037 3216
rect 1044 3213 1061 3216
rect 1066 3213 1085 3216
rect 1172 3213 1189 3216
rect 1394 3213 1453 3216
rect 1490 3213 1572 3216
rect 1722 3213 1756 3216
rect 1802 3213 1828 3216
rect 2036 3213 2069 3216
rect 2140 3213 2148 3216
rect 2186 3213 2196 3216
rect 2284 3213 2309 3216
rect 2314 3213 2317 3243
rect 3426 3233 3469 3236
rect 3484 3233 3493 3236
rect 2820 3223 2861 3226
rect 2938 3223 2972 3226
rect 3354 3223 3364 3226
rect 2426 3213 2460 3216
rect 2492 3213 2517 3216
rect 2564 3213 2573 3216
rect 2626 3213 2660 3216
rect 2692 3213 2701 3216
rect 2732 3213 2741 3216
rect 2858 3213 2876 3216
rect 2994 3213 3069 3216
rect 3100 3213 3117 3216
rect 3194 3213 3220 3216
rect 3250 3213 3276 3216
rect 3426 3215 3429 3233
rect 3450 3223 3476 3226
rect 3538 3223 3556 3226
rect 3580 3223 3605 3226
rect 3620 3213 3637 3216
rect 3684 3213 3717 3216
rect 3756 3213 3773 3216
rect 3786 3213 3796 3216
rect 3954 3213 4085 3216
rect 4252 3213 4277 3216
rect 4308 3213 4317 3216
rect 4324 3213 4373 3216
rect 4434 3213 4444 3216
rect 4482 3213 4492 3216
rect 4652 3213 4661 3216
rect 4706 3213 4716 3216
rect 92 3203 117 3206
rect 372 3203 405 3206
rect 428 3203 469 3206
rect 570 3203 596 3206
rect 786 3203 805 3206
rect 810 3203 884 3206
rect 980 3203 1013 3206
rect 1052 3203 1077 3206
rect 1082 3205 1085 3213
rect 1114 3203 1133 3206
rect 1164 3203 1173 3206
rect 1178 3203 1356 3206
rect 1380 3203 1445 3206
rect 1450 3205 1453 3213
rect 1484 3203 1525 3206
rect 1554 3203 1564 3206
rect 1596 3203 1676 3206
rect 1708 3203 1749 3206
rect 1906 3203 1949 3206
rect 1954 3203 1980 3206
rect 2042 3203 2084 3206
rect 2194 3203 2204 3206
rect 2290 3203 2332 3206
rect 2348 3203 2396 3206
rect 2484 3203 2525 3206
rect 2626 3203 2668 3206
rect 2690 3203 2724 3206
rect 2738 3203 2796 3206
rect 2820 3203 2845 3206
rect 2858 3203 2861 3213
rect 2892 3203 2909 3206
rect 2930 3203 2972 3206
rect 2994 3205 2997 3213
rect 3634 3206 3637 3213
rect 3028 3203 3037 3206
rect 3122 3203 3156 3206
rect 3634 3203 3660 3206
rect 3682 3203 3732 3206
rect 3748 3203 3765 3206
rect 3770 3203 3804 3206
rect 3820 3203 3845 3206
rect 3890 3203 3916 3206
rect 3948 3203 3989 3206
rect 3994 3203 4012 3206
rect 4082 3203 4085 3213
rect 4314 3205 4317 3213
rect 4330 3203 4372 3206
rect 4404 3203 4429 3206
rect 4698 3203 4708 3206
rect 802 3196 805 3203
rect 802 3193 861 3196
rect 922 3193 972 3196
rect 994 3193 1021 3196
rect 38 3167 4829 3173
rect 842 3143 892 3146
rect 2882 3143 2940 3146
rect 546 3133 556 3136
rect 642 3133 652 3136
rect 124 3123 149 3126
rect 180 3123 197 3126
rect 340 3123 365 3126
rect 396 3123 421 3126
rect 484 3123 509 3126
rect 618 3123 660 3126
rect 786 3125 789 3136
rect 812 3133 829 3136
rect 836 3133 877 3136
rect 914 3133 956 3136
rect 844 3123 885 3126
rect 908 3123 917 3126
rect 954 3123 964 3126
rect 978 3123 987 3126
rect 1018 3125 1021 3136
rect 1138 3133 1164 3136
rect 1186 3133 1252 3136
rect 1276 3133 1293 3136
rect 1298 3133 1324 3136
rect 1348 3133 1389 3136
rect 1138 3126 1141 3133
rect 1506 3126 1509 3135
rect 1522 3133 1564 3136
rect 1596 3133 1645 3136
rect 1708 3133 1749 3136
rect 1852 3133 1933 3136
rect 1938 3133 1948 3136
rect 1964 3133 2044 3136
rect 2076 3133 2093 3136
rect 2148 3133 2157 3136
rect 2170 3133 2188 3136
rect 2260 3133 2269 3136
rect 2426 3133 2452 3136
rect 2466 3133 2508 3136
rect 2530 3133 2564 3136
rect 2578 3133 2628 3136
rect 2650 3133 2684 3136
rect 2850 3126 2853 3135
rect 2876 3133 2925 3136
rect 2948 3133 2981 3136
rect 2986 3133 3004 3136
rect 3034 3133 3076 3136
rect 1116 3123 1149 3126
rect 1188 3123 1253 3126
rect 1268 3123 1293 3126
rect 1340 3123 1373 3126
rect 1428 3123 1445 3126
rect 1484 3123 1509 3126
rect 1516 3123 1557 3126
rect 1588 3123 1597 3126
rect 1722 3123 1756 3126
rect 1866 3123 1940 3126
rect 2122 3123 2132 3126
rect 2178 3123 2196 3126
rect 2202 3123 2236 3126
rect 2378 3123 2396 3126
rect 2466 3123 2500 3126
rect 2532 3123 2549 3126
rect 2578 3123 2620 3126
rect 2652 3123 2661 3126
rect 2692 3123 2709 3126
rect 2804 3123 2853 3126
rect 3098 3126 3101 3135
rect 3140 3133 3181 3136
rect 3220 3133 3293 3136
rect 3356 3133 3365 3136
rect 3610 3126 3613 3135
rect 3626 3133 3660 3136
rect 3698 3133 3732 3136
rect 3882 3126 3885 3135
rect 4042 3133 4076 3136
rect 4108 3133 4125 3136
rect 4164 3133 4181 3136
rect 4276 3133 4317 3136
rect 4356 3133 4373 3136
rect 4468 3133 4493 3136
rect 4524 3133 4533 3136
rect 4636 3133 4653 3136
rect 4490 3126 4493 3133
rect 3098 3123 3181 3126
rect 3212 3123 3245 3126
rect 3282 3123 3348 3126
rect 3404 3123 3413 3126
rect 3460 3123 3493 3126
rect 3532 3123 3557 3126
rect 3588 3123 3613 3126
rect 3620 3123 3637 3126
rect 3706 3123 3740 3126
rect 3876 3123 3885 3126
rect 4114 3123 4148 3126
rect 4170 3123 4196 3126
rect 4226 3123 4268 3126
rect 4274 3123 4332 3126
rect 4362 3123 4396 3126
rect 4418 3123 4444 3126
rect 4490 3123 4516 3126
rect 4586 3123 4661 3126
rect 3242 3116 3245 3123
rect 1314 3113 1324 3116
rect 2876 3113 2933 3116
rect 2970 3113 3004 3116
rect 3034 3113 3076 3116
rect 3242 3113 3301 3116
rect 14 3067 4853 3073
rect 1026 3053 1045 3056
rect 916 3023 973 3026
rect 1180 3023 1189 3026
rect 2908 3023 2989 3026
rect 178 3013 188 3016
rect 180 3003 189 3006
rect 250 3003 260 3006
rect 290 3005 293 3016
rect 362 3013 396 3016
rect 402 3013 444 3016
rect 476 3013 517 3016
rect 404 3003 413 3006
rect 418 3003 452 3006
rect 468 3003 485 3006
rect 522 3003 525 3014
rect 556 3013 565 3016
rect 740 3013 749 3016
rect 796 3013 821 3016
rect 914 3013 980 3016
rect 1012 3013 1021 3016
rect 1092 3013 1157 3016
rect 818 3006 821 3013
rect 1186 3006 1189 3023
rect 1260 3013 1293 3016
rect 1356 3013 1381 3016
rect 1412 3013 1437 3016
rect 1532 3013 1557 3016
rect 1644 3013 1669 3016
rect 1700 3013 1733 3016
rect 1740 3013 1749 3016
rect 1754 3013 1764 3016
rect 594 3003 628 3006
rect 660 3003 669 3006
rect 818 3003 892 3006
rect 916 3003 925 3006
rect 930 3003 988 3006
rect 1004 3003 1077 3006
rect 1084 3003 1117 3006
rect 1146 3003 1156 3006
rect 1186 3003 1244 3006
rect 1268 3003 1317 3006
rect 1434 3005 1437 3013
rect 1540 3003 1597 3006
rect 1730 3005 1733 3013
rect 1842 3006 1845 3016
rect 1884 3013 1901 3016
rect 2188 3013 2221 3016
rect 2266 3013 2308 3016
rect 2340 3013 2381 3016
rect 2386 3013 2404 3016
rect 2532 3013 2541 3016
rect 2588 3013 2605 3016
rect 2652 3013 2661 3016
rect 2692 3013 2701 3016
rect 2866 3013 2892 3016
rect 3034 3013 3124 3016
rect 2386 3006 2389 3013
rect 1842 3003 1876 3006
rect 2084 3003 2101 3006
rect 2154 3003 2164 3006
rect 2180 3003 2229 3006
rect 2332 3003 2389 3006
rect 2650 3003 2684 3006
rect 2836 3003 2845 3006
rect 2858 3003 2884 3006
rect 2908 3003 2957 3006
rect 3132 3003 3141 3006
rect 3226 3003 3276 3006
rect 3458 3003 3461 3014
rect 3538 3013 3588 3016
rect 3738 3013 3764 3016
rect 3988 3013 4013 3016
rect 4018 3013 4060 3016
rect 4170 3013 4188 3016
rect 4524 3013 4549 3016
rect 4626 3013 4652 3016
rect 3484 3003 3493 3006
rect 3554 3003 3580 3006
rect 4026 3003 4052 3006
rect 4162 3003 4180 3006
rect 4610 3003 4644 3006
rect 4676 3003 4693 3006
rect 1026 2993 1076 2996
rect 1098 2993 1149 2996
rect 2098 2993 2149 2996
rect 2226 2993 2285 2996
rect 2090 2983 2117 2986
rect 38 2967 4829 2973
rect 1402 2953 1429 2956
rect 754 2943 828 2946
rect 874 2943 909 2946
rect 946 2943 1132 2946
rect 2874 2943 2908 2946
rect 2922 2943 2965 2946
rect 906 2936 909 2943
rect 2922 2936 2925 2943
rect 162 2933 196 2936
rect 218 2933 252 2936
rect 412 2933 461 2936
rect 490 2933 525 2936
rect 538 2933 548 2936
rect 836 2933 901 2936
rect 906 2933 916 2936
rect 940 2933 949 2936
rect 1122 2933 1140 2936
rect 1178 2933 1196 2936
rect 1220 2933 1229 2936
rect 1322 2933 1364 2936
rect 178 2923 188 2926
rect 220 2923 237 2926
rect 340 2923 365 2926
rect 442 2923 460 2926
rect 490 2925 493 2933
rect 1386 2926 1389 2935
rect 1460 2933 1469 2936
rect 1506 2933 1524 2936
rect 1556 2933 1581 2936
rect 1938 2933 1948 2936
rect 1980 2933 2005 2936
rect 2100 2933 2141 2936
rect 514 2923 556 2926
rect 580 2923 605 2926
rect 740 2923 749 2926
rect 844 2923 917 2926
rect 1148 2923 1197 2926
rect 1386 2923 1461 2926
rect 1548 2923 1557 2926
rect 1578 2923 1588 2926
rect 1618 2923 1644 2926
rect 1722 2923 1756 2926
rect 1802 2923 1836 2926
rect 1868 2923 1877 2926
rect 1906 2923 1956 2926
rect 2092 2923 2125 2926
rect 2146 2925 2149 2936
rect 2178 2933 2221 2936
rect 2330 2933 2356 2936
rect 2402 2933 2428 2936
rect 2548 2933 2581 2936
rect 2626 2933 2668 2936
rect 2684 2933 2717 2936
rect 2818 2933 2836 2936
rect 2860 2933 2909 2936
rect 2916 2933 2925 2936
rect 2930 2933 2972 2936
rect 2996 2933 3037 2936
rect 3076 2933 3085 2936
rect 3300 2933 3325 2936
rect 3362 2933 3516 2936
rect 3548 2933 3557 2936
rect 3620 2933 3661 2936
rect 3692 2933 3709 2936
rect 3714 2933 3740 2936
rect 3756 2933 3837 2936
rect 3898 2933 3940 2936
rect 3972 2933 3981 2936
rect 4010 2933 4028 2936
rect 4074 2933 4092 2936
rect 4124 2933 4133 2936
rect 4202 2933 4252 2936
rect 4268 2933 4301 2936
rect 4332 2933 4349 2936
rect 4354 2933 4364 2936
rect 2178 2925 2181 2933
rect 3714 2926 3717 2933
rect 2186 2923 2228 2926
rect 2266 2923 2284 2926
rect 2474 2923 2500 2926
rect 2562 2923 2580 2926
rect 2618 2923 2660 2926
rect 2834 2923 2844 2926
rect 2988 2923 3013 2926
rect 3170 2923 3196 2926
rect 3292 2923 3301 2926
rect 3514 2923 3524 2926
rect 3602 2923 3612 2926
rect 3650 2923 3717 2926
rect 3722 2923 3732 2926
rect 3764 2923 3829 2926
rect 3834 2923 3837 2933
rect 4298 2926 4301 2933
rect 3890 2923 3948 2926
rect 4018 2923 4036 2926
rect 4116 2923 4172 2926
rect 4218 2923 4244 2926
rect 4276 2923 4285 2926
rect 4298 2923 4357 2926
rect 4394 2923 4397 2935
rect 4402 2933 4445 2936
rect 4468 2933 4509 2936
rect 4532 2933 4565 2936
rect 4570 2933 4580 2936
rect 4756 2933 4765 2936
rect 4442 2925 4445 2933
rect 4506 2926 4509 2933
rect 4476 2923 4485 2926
rect 4506 2923 4573 2926
rect 4604 2923 4621 2926
rect 4666 2923 4748 2926
rect 940 2913 957 2916
rect 1250 2913 1276 2916
rect 1354 2913 1364 2916
rect 2860 2913 2893 2916
rect 3770 2913 3844 2916
rect 3868 2913 3925 2916
rect 2050 2893 2085 2896
rect 14 2867 4853 2873
rect 3284 2833 3301 2836
rect 3428 2833 3453 2836
rect 794 2823 805 2826
rect 956 2823 1013 2826
rect 2820 2823 2861 2826
rect 2892 2823 2925 2826
rect 2970 2823 2996 2826
rect 3266 2823 3276 2826
rect 3300 2823 3333 2826
rect 3386 2823 3420 2826
rect 3444 2823 3477 2826
rect 802 2816 805 2823
rect 92 2813 157 2816
rect 252 2813 261 2816
rect 380 2813 389 2816
rect 492 2813 517 2816
rect 562 2814 572 2816
rect 562 2813 573 2814
rect 604 2813 629 2816
rect 788 2813 797 2816
rect 802 2813 812 2816
rect 962 2813 1020 2816
rect 1058 2813 1140 2816
rect 1252 2813 1277 2816
rect 1308 2813 1325 2816
rect 1372 2813 1389 2816
rect 1682 2813 1692 2816
rect 1802 2813 1828 2816
rect 1884 2813 1901 2816
rect 2260 2813 2269 2816
rect 2330 2813 2364 2816
rect 2396 2813 2413 2816
rect 2444 2813 2453 2816
rect 2490 2813 2516 2816
rect 2554 2813 2596 2816
rect 2628 2813 2645 2816
rect 2692 2813 2717 2816
rect 2732 2813 2757 2816
rect 2778 2813 2804 2816
rect 2842 2813 2876 2816
rect 3034 2813 3060 2816
rect 3212 2813 3253 2816
rect 3354 2813 3364 2816
rect 3508 2813 3517 2816
rect 3666 2813 3684 2816
rect 3778 2813 3820 2816
rect 3850 2813 3884 2816
rect 3914 2813 3940 2816
rect 3986 2813 4012 2816
rect 4172 2813 4197 2816
rect 4268 2813 4277 2816
rect 4324 2813 4333 2816
rect 4346 2813 4372 2816
rect 4402 2813 4428 2816
rect 4466 2813 4476 2816
rect 4570 2813 4580 2816
rect 4610 2813 4636 2816
rect 258 2806 261 2813
rect 100 2803 157 2806
rect 258 2803 276 2806
rect 292 2803 333 2806
rect 570 2803 573 2813
rect 794 2806 797 2813
rect 596 2803 693 2806
rect 794 2803 820 2806
rect 882 2803 932 2806
rect 956 2803 965 2806
rect 1044 2803 1093 2806
rect 1106 2803 1148 2806
rect 1164 2803 1173 2806
rect 1338 2803 1356 2806
rect 1380 2803 1461 2806
rect 1506 2803 1588 2806
rect 1620 2803 1677 2806
rect 1836 2803 1845 2806
rect 1946 2803 1964 2806
rect 1986 2803 2004 2806
rect 2338 2803 2372 2806
rect 2402 2803 2436 2806
rect 2586 2803 2604 2806
rect 2620 2803 2629 2806
rect 2634 2803 2684 2806
rect 2698 2803 2724 2806
rect 2746 2803 2796 2806
rect 2820 2803 2845 2806
rect 2892 2803 2933 2806
rect 2940 2803 2949 2806
rect 2954 2803 2996 2806
rect 3020 2803 3045 2806
rect 3084 2803 3109 2806
rect 3250 2805 3253 2813
rect 3516 2803 3525 2806
rect 3692 2803 3701 2806
rect 3714 2803 3812 2806
rect 3844 2803 3876 2806
rect 3970 2803 4020 2806
rect 4036 2803 4077 2806
rect 4194 2805 4197 2813
rect 4330 2805 4333 2813
rect 4492 2803 4541 2806
rect 4780 2803 4789 2806
rect 2906 2793 2932 2796
rect 38 2767 4829 2773
rect 826 2736 829 2746
rect 834 2743 860 2746
rect 2802 2743 2828 2746
rect 196 2733 221 2736
rect 404 2733 413 2736
rect 436 2733 500 2736
rect 690 2733 700 2736
rect 124 2723 149 2726
rect 202 2723 220 2726
rect 386 2723 396 2726
rect 722 2725 725 2736
rect 804 2733 829 2736
rect 868 2733 973 2736
rect 1130 2733 1140 2736
rect 1292 2733 1325 2736
rect 1388 2733 1461 2736
rect 1500 2733 1533 2736
rect 970 2726 973 2733
rect 1658 2726 1661 2735
rect 1682 2733 1708 2736
rect 1804 2733 1829 2736
rect 1826 2726 1829 2733
rect 1890 2733 1901 2736
rect 1924 2733 1941 2736
rect 2082 2733 2124 2736
rect 2140 2733 2157 2736
rect 2234 2733 2244 2736
rect 1890 2726 1893 2733
rect 2266 2726 2269 2736
rect 2338 2733 2372 2736
rect 2618 2733 2652 2736
rect 2858 2733 2876 2736
rect 2900 2733 2909 2736
rect 2914 2733 2940 2736
rect 2970 2733 2996 2736
rect 3020 2733 3061 2736
rect 3100 2733 3132 2736
rect 3164 2733 3181 2736
rect 3202 2733 3212 2736
rect 3434 2733 3492 2736
rect 3514 2733 3581 2736
rect 3914 2726 3917 2735
rect 4242 2726 4245 2735
rect 4322 2733 4348 2736
rect 4506 2733 4525 2736
rect 4548 2733 4581 2736
rect 4610 2733 4644 2736
rect 4676 2733 4693 2736
rect 730 2723 796 2726
rect 876 2723 965 2726
rect 970 2723 1028 2726
rect 1060 2723 1069 2726
rect 1148 2723 1157 2726
rect 1210 2723 1228 2726
rect 1274 2723 1293 2726
rect 1380 2723 1389 2726
rect 1588 2723 1597 2726
rect 1644 2723 1661 2726
rect 1724 2723 1740 2726
rect 1826 2723 1837 2726
rect 1844 2723 1893 2726
rect 1932 2723 1941 2726
rect 2074 2723 2116 2726
rect 2148 2723 2245 2726
rect 2252 2723 2269 2726
rect 2324 2723 2365 2726
rect 2442 2723 2452 2726
rect 2482 2723 2508 2726
rect 2554 2723 2580 2726
rect 2612 2723 2645 2726
rect 2660 2723 2693 2726
rect 2732 2723 2741 2726
rect 2788 2723 2813 2726
rect 2866 2723 2884 2726
rect 2922 2723 2941 2726
rect 3034 2723 3076 2726
rect 3210 2723 3220 2726
rect 1298 2713 1364 2716
rect 2900 2713 2933 2716
rect 2938 2715 2941 2723
rect 2970 2713 2996 2716
rect 3402 2706 3405 2725
rect 3474 2723 3484 2726
rect 3420 2713 3469 2716
rect 3386 2703 3405 2706
rect 3754 2706 3757 2725
rect 3884 2723 3917 2726
rect 4156 2723 4181 2726
rect 4212 2723 4245 2726
rect 4308 2723 4341 2726
rect 4386 2723 4396 2726
rect 4426 2723 4452 2726
rect 4522 2725 4525 2733
rect 4570 2723 4621 2726
rect 4626 2723 4652 2726
rect 3764 2713 3789 2716
rect 3930 2713 3972 2716
rect 3996 2713 4029 2716
rect 4074 2713 4084 2716
rect 3754 2703 3789 2706
rect 4068 2703 4077 2706
rect 14 2667 4853 2673
rect 1218 2653 1253 2656
rect 4058 2633 4085 2636
rect 780 2623 829 2626
rect 1100 2623 1157 2626
rect 108 2613 133 2616
rect 178 2613 188 2616
rect 180 2603 189 2606
rect 218 2603 221 2614
rect 324 2613 349 2616
rect 388 2613 413 2616
rect 444 2613 461 2616
rect 514 2613 548 2616
rect 666 2613 708 2616
rect 906 2606 909 2614
rect 940 2613 949 2616
rect 1020 2613 1061 2616
rect 1066 2613 1084 2616
rect 1098 2613 1125 2616
rect 1170 2613 1173 2625
rect 1218 2623 1284 2626
rect 2828 2623 2845 2626
rect 3370 2623 3404 2626
rect 3428 2623 3461 2626
rect 4066 2623 4076 2626
rect 1188 2613 1285 2616
rect 1300 2613 1389 2616
rect 1460 2613 1485 2616
rect 1516 2613 1541 2616
rect 1548 2613 1557 2616
rect 1562 2613 1661 2616
rect 1772 2613 1781 2616
rect 1874 2613 1900 2616
rect 1938 2613 1980 2616
rect 2140 2613 2213 2616
rect 2274 2614 2332 2616
rect 2274 2613 2333 2614
rect 2364 2613 2413 2616
rect 2530 2613 2573 2616
rect 2778 2613 2812 2616
rect 2884 2613 2909 2616
rect 2940 2613 2957 2616
rect 3012 2613 3037 2616
rect 3068 2613 3101 2616
rect 3244 2613 3253 2616
rect 3292 2613 3301 2616
rect 3348 2613 3357 2616
rect 3364 2613 3397 2616
rect 3666 2613 3692 2616
rect 3810 2613 3860 2616
rect 3890 2613 3916 2616
rect 3946 2613 3964 2616
rect 3994 2613 4020 2616
rect 4082 2615 4085 2633
rect 4100 2623 4125 2626
rect 4148 2613 4172 2616
rect 4194 2613 4228 2616
rect 4266 2613 4284 2616
rect 4514 2613 4532 2616
rect 4612 2613 4668 2616
rect 4698 2613 4708 2616
rect 236 2603 268 2606
rect 450 2603 476 2606
rect 492 2603 540 2606
rect 628 2603 677 2606
rect 690 2603 700 2606
rect 722 2603 756 2606
rect 780 2603 837 2606
rect 844 2603 909 2606
rect 932 2603 949 2606
rect 1042 2603 1076 2606
rect 1106 2603 1172 2606
rect 1196 2603 1229 2606
rect 1234 2603 1284 2606
rect 1308 2603 1349 2606
rect 1538 2605 1541 2613
rect 1620 2603 1629 2606
rect 1650 2603 1668 2606
rect 1700 2603 1717 2606
rect 1852 2603 1901 2606
rect 1994 2603 2028 2606
rect 2060 2603 2117 2606
rect 2122 2603 2132 2606
rect 2162 2603 2228 2606
rect 2244 2603 2309 2606
rect 2330 2603 2333 2613
rect 2356 2603 2444 2606
rect 2882 2603 2924 2606
rect 2948 2603 2973 2606
rect 3098 2605 3101 2613
rect 3354 2605 3357 2613
rect 3442 2603 3476 2606
rect 3508 2603 3525 2606
rect 3716 2603 3765 2606
rect 3804 2603 3853 2606
rect 3868 2603 3901 2606
rect 3940 2603 3957 2606
rect 4106 2603 4132 2606
rect 4188 2603 4205 2606
rect 4258 2603 4292 2606
rect 4476 2603 4485 2606
rect 4556 2603 4589 2606
rect 4618 2603 4660 2606
rect 4732 2603 4781 2606
rect 1226 2596 1229 2603
rect 794 2593 836 2596
rect 954 2593 1004 2596
rect 1226 2593 1277 2596
rect 2834 2593 2868 2596
rect 38 2567 4829 2573
rect 858 2543 908 2546
rect 132 2533 165 2536
rect 188 2533 213 2536
rect 284 2533 317 2536
rect 340 2533 357 2536
rect 380 2533 429 2536
rect 114 2523 124 2526
rect 154 2523 164 2526
rect 196 2523 245 2526
rect 258 2523 276 2526
rect 378 2523 436 2526
rect 442 2523 445 2534
rect 730 2533 772 2536
rect 788 2533 829 2536
rect 834 2533 844 2536
rect 916 2533 957 2536
rect 1010 2533 1069 2536
rect 1092 2533 1109 2536
rect 450 2523 476 2526
rect 746 2523 764 2526
rect 852 2523 885 2526
rect 924 2523 965 2526
rect 1066 2525 1069 2533
rect 1130 2523 1188 2526
rect 1218 2525 1221 2536
rect 1530 2534 1580 2536
rect 1370 2526 1373 2534
rect 1530 2533 1581 2534
rect 1842 2533 1876 2536
rect 1906 2533 1916 2536
rect 1250 2523 1284 2526
rect 1338 2523 1364 2526
rect 1370 2523 1420 2526
rect 1516 2523 1549 2526
rect 1578 2523 1581 2533
rect 1588 2523 1597 2526
rect 1626 2523 1636 2526
rect 1682 2523 1692 2526
rect 1780 2523 1805 2526
rect 1842 2523 1884 2526
rect 1898 2523 1924 2526
rect 1964 2523 1981 2526
rect 2076 2523 2085 2526
rect 2098 2523 2124 2526
rect 2154 2523 2164 2526
rect 2210 2523 2220 2526
rect 996 2513 1061 2516
rect 1346 2513 1356 2516
rect 2274 2483 2277 2546
rect 2770 2543 2821 2546
rect 2874 2543 2900 2546
rect 2386 2533 2428 2536
rect 2570 2533 2612 2536
rect 2324 2523 2333 2526
rect 2402 2523 2436 2526
rect 2466 2523 2540 2526
rect 2572 2523 2613 2526
rect 2620 2523 2653 2526
rect 2770 2525 2773 2543
rect 2852 2533 2893 2536
rect 2908 2533 2917 2536
rect 2922 2533 2964 2536
rect 2988 2533 3037 2536
rect 3076 2533 3109 2536
rect 3226 2526 3229 2535
rect 3324 2533 3341 2536
rect 3372 2533 3381 2536
rect 3444 2533 3461 2536
rect 3466 2533 3492 2536
rect 3634 2533 3660 2536
rect 3338 2526 3341 2533
rect 3466 2526 3469 2533
rect 3890 2526 3893 2535
rect 4122 2533 4140 2536
rect 4346 2533 4364 2536
rect 4428 2533 4445 2536
rect 4482 2533 4517 2536
rect 4540 2533 4557 2536
rect 2778 2523 2836 2526
rect 3212 2523 3229 2526
rect 3236 2523 3245 2526
rect 3290 2523 3308 2526
rect 3338 2523 3356 2526
rect 3378 2523 3404 2526
rect 3458 2523 3469 2526
rect 3482 2523 3500 2526
rect 3530 2523 3620 2526
rect 3674 2523 3700 2526
rect 3876 2523 3893 2526
rect 4010 2523 4028 2526
rect 4164 2523 4197 2526
rect 2852 2513 2893 2516
rect 2930 2513 2964 2516
rect 4186 2513 4220 2516
rect 4234 2506 4237 2525
rect 4332 2523 4372 2526
rect 4402 2523 4420 2526
rect 4514 2525 4517 2533
rect 4668 2523 4685 2526
rect 4250 2513 4276 2516
rect 4434 2513 4452 2516
rect 4250 2506 4253 2513
rect 4234 2503 4253 2506
rect 4450 2503 4468 2506
rect 14 2467 4853 2473
rect 3322 2433 3349 2436
rect 3386 2433 3405 2436
rect 788 2423 829 2426
rect 946 2423 973 2426
rect 1242 2423 1316 2426
rect 1858 2423 1909 2426
rect 3290 2423 3308 2426
rect 946 2416 949 2423
rect 108 2413 117 2416
rect 172 2413 181 2416
rect 252 2413 261 2416
rect 308 2413 325 2416
rect 364 2413 373 2416
rect 420 2413 429 2416
rect 474 2413 500 2416
rect 530 2413 572 2416
rect 626 2413 636 2416
rect 642 2413 684 2416
rect 754 2413 772 2416
rect 868 2413 885 2416
rect 924 2413 949 2416
rect 954 2413 980 2416
rect 1082 2413 1092 2416
rect 1124 2413 1189 2416
rect 1228 2413 1237 2416
rect 1332 2413 1341 2416
rect 1420 2413 1445 2416
rect 1476 2413 1509 2416
rect 1722 2413 1732 2416
rect 1844 2413 1901 2416
rect 1956 2413 2029 2416
rect 2076 2413 2093 2416
rect 2274 2413 2300 2416
rect 426 2406 429 2413
rect 180 2403 189 2406
rect 426 2403 444 2406
rect 482 2403 492 2406
rect 524 2403 533 2406
rect 596 2403 605 2406
rect 610 2403 628 2406
rect 642 2403 692 2406
rect 722 2403 764 2406
rect 788 2403 797 2406
rect 1004 2403 1013 2406
rect 1034 2403 1100 2406
rect 1116 2403 1133 2406
rect 1154 2403 1212 2406
rect 1236 2403 1301 2406
rect 1306 2403 1316 2406
rect 1340 2403 1373 2406
rect 1506 2405 1509 2413
rect 2378 2406 2381 2416
rect 2516 2413 2557 2416
rect 2578 2413 2628 2416
rect 2732 2413 2749 2416
rect 3042 2413 3052 2416
rect 3084 2413 3148 2416
rect 3188 2413 3220 2416
rect 3322 2415 3325 2433
rect 3332 2423 3365 2426
rect 3386 2415 3389 2433
rect 3402 2426 3405 2433
rect 3402 2423 3436 2426
rect 3460 2423 3501 2426
rect 4476 2423 4509 2426
rect 3474 2413 3508 2416
rect 3578 2413 3596 2416
rect 3626 2413 3652 2416
rect 3658 2413 3700 2416
rect 3730 2413 3756 2416
rect 3794 2413 3820 2416
rect 3842 2413 3860 2416
rect 3898 2413 3940 2416
rect 3970 2413 3988 2416
rect 1578 2403 1588 2406
rect 1620 2403 1669 2406
rect 1836 2403 1932 2406
rect 2068 2403 2085 2406
rect 2114 2403 2164 2406
rect 2180 2403 2189 2406
rect 2324 2403 2381 2406
rect 2450 2403 2508 2406
rect 2580 2403 2636 2406
rect 2652 2403 2709 2406
rect 2714 2403 2724 2406
rect 3034 2403 3044 2406
rect 3106 2403 3140 2406
rect 3242 2403 3268 2406
rect 3506 2403 3516 2406
rect 3554 2403 3588 2406
rect 3620 2403 3645 2406
rect 3658 2405 3661 2413
rect 3858 2403 3868 2406
rect 3884 2403 3925 2406
rect 3964 2403 3981 2406
rect 3994 2405 3997 2416
rect 4050 2413 4076 2416
rect 4178 2413 4204 2416
rect 4324 2413 4333 2416
rect 4340 2413 4365 2416
rect 4370 2413 4380 2416
rect 4514 2413 4524 2416
rect 4570 2413 4588 2416
rect 4618 2413 4644 2416
rect 4330 2405 4333 2413
rect 4362 2406 4365 2413
rect 4362 2403 4388 2406
rect 4404 2403 4421 2406
rect 4506 2403 4516 2406
rect 4548 2403 4581 2406
rect 1034 2393 1037 2403
rect 1306 2396 1309 2403
rect 1274 2393 1309 2396
rect 1850 2393 1885 2396
rect 2858 2393 2876 2396
rect 1994 2383 2021 2386
rect 2354 2383 2477 2386
rect 38 2367 4829 2373
rect 858 2343 900 2346
rect 428 2333 437 2336
rect 620 2333 637 2336
rect 634 2326 637 2333
rect 826 2326 829 2334
rect 852 2333 885 2336
rect 908 2333 989 2336
rect 1012 2333 1053 2336
rect 1098 2333 1124 2336
rect 1228 2333 1285 2336
rect 1324 2333 1349 2336
rect 108 2323 133 2326
rect 244 2323 269 2326
rect 356 2323 381 2326
rect 468 2323 476 2326
rect 548 2323 589 2326
rect 634 2323 644 2326
rect 674 2323 700 2326
rect 778 2323 829 2326
rect 916 2323 925 2326
rect 986 2325 989 2333
rect 1554 2326 1557 2334
rect 1740 2333 1757 2336
rect 1804 2333 1821 2336
rect 1876 2333 1901 2336
rect 2034 2333 2084 2336
rect 2172 2333 2197 2336
rect 2210 2333 2244 2336
rect 2324 2333 2373 2336
rect 2434 2333 2468 2336
rect 2778 2333 2788 2336
rect 1148 2323 1157 2326
rect 1178 2323 1212 2326
rect 1298 2323 1316 2326
rect 1322 2323 1548 2326
rect 1554 2323 1580 2326
rect 1610 2323 1636 2326
rect 1706 2323 1732 2326
rect 1738 2323 1796 2326
rect 1884 2323 1909 2326
rect 1930 2323 1940 2326
rect 2122 2323 2132 2326
rect 2242 2323 2252 2326
rect 2370 2323 2373 2333
rect 2810 2326 2813 2334
rect 2818 2333 2868 2336
rect 2954 2326 2957 2334
rect 2980 2333 3037 2336
rect 3076 2333 3093 2336
rect 3106 2333 3116 2336
rect 3146 2333 3164 2336
rect 3212 2333 3229 2336
rect 3346 2326 3349 2334
rect 3362 2333 3404 2336
rect 3442 2333 3492 2336
rect 3674 2326 3677 2334
rect 3834 2333 3845 2336
rect 3868 2333 3917 2336
rect 4012 2333 4021 2336
rect 3842 2326 3845 2333
rect 4234 2326 4237 2334
rect 4258 2333 4276 2336
rect 4308 2333 4341 2336
rect 4362 2333 4380 2336
rect 4396 2333 4421 2336
rect 4532 2333 4541 2336
rect 4596 2333 4621 2336
rect 4660 2333 4677 2336
rect 4716 2333 4781 2336
rect 2378 2323 2396 2326
rect 2428 2323 2469 2326
rect 2476 2323 2501 2326
rect 2506 2323 2540 2326
rect 2570 2323 2596 2326
rect 2684 2323 2693 2326
rect 2786 2323 2796 2326
rect 2810 2323 2845 2326
rect 2866 2323 2876 2326
rect 2946 2323 2957 2326
rect 3068 2323 3085 2326
rect 3140 2323 3157 2326
rect 3276 2323 3301 2326
rect 3332 2323 3349 2326
rect 3428 2323 3500 2326
rect 3660 2323 3677 2326
rect 3826 2325 3845 2326
rect 3826 2323 3844 2325
rect 3876 2323 3925 2326
rect 3962 2323 4004 2326
rect 4212 2323 4237 2326
rect 4404 2323 4413 2326
rect 4482 2323 4508 2326
rect 4540 2323 4549 2326
rect 4602 2323 4636 2326
rect 4666 2323 4708 2326
rect 2946 2316 2949 2323
rect 2812 2313 2861 2316
rect 2892 2313 2949 2316
rect 4410 2313 4452 2316
rect 4426 2303 4468 2306
rect 14 2267 4853 2273
rect 930 2243 957 2246
rect 2554 2243 2589 2246
rect 3282 2243 3325 2246
rect 3522 2243 3581 2246
rect 3714 2233 3741 2236
rect 1172 2223 1245 2226
rect 1250 2223 1260 2226
rect 2890 2223 2908 2226
rect 4476 2223 4501 2226
rect 108 2213 133 2216
rect 178 2213 188 2216
rect 180 2203 189 2206
rect 218 2203 221 2214
rect 260 2213 277 2216
rect 316 2213 325 2216
rect 396 2213 421 2216
rect 436 2213 469 2216
rect 538 2213 564 2216
rect 602 2213 612 2216
rect 714 2213 740 2216
rect 908 2213 941 2216
rect 370 2203 380 2206
rect 402 2203 428 2206
rect 458 2203 468 2206
rect 634 2203 644 2206
rect 700 2203 733 2206
rect 764 2203 781 2206
rect 962 2203 965 2214
rect 996 2213 1021 2216
rect 1060 2213 1141 2216
rect 1242 2206 1245 2223
rect 1276 2213 1309 2216
rect 1500 2213 1517 2216
rect 1594 2213 1612 2216
rect 1994 2213 2028 2216
rect 2122 2213 2148 2216
rect 2410 2206 2413 2214
rect 2426 2213 2452 2216
rect 2498 2213 2508 2216
rect 2546 2213 2596 2216
rect 2628 2213 2661 2216
rect 2924 2213 2933 2216
rect 3028 2213 3053 2216
rect 3204 2213 3221 2216
rect 3282 2213 3332 2216
rect 3436 2213 3477 2216
rect 3482 2206 3485 2214
rect 3516 2213 3533 2216
rect 3594 2213 3612 2216
rect 3626 2213 3684 2216
rect 3714 2213 3764 2216
rect 3812 2213 3837 2216
rect 3868 2213 3877 2216
rect 3970 2213 4044 2216
rect 4082 2213 4140 2216
rect 4226 2213 4252 2216
rect 4290 2213 4316 2216
rect 4338 2213 4381 2216
rect 4418 2213 4436 2216
rect 4482 2213 4516 2216
rect 4554 2213 4564 2216
rect 988 2203 997 2206
rect 1002 2203 1052 2206
rect 1058 2203 1148 2206
rect 1172 2203 1181 2206
rect 1242 2203 1260 2206
rect 1284 2203 1301 2206
rect 1466 2203 1476 2206
rect 1508 2203 1533 2206
rect 1690 2203 1700 2206
rect 1732 2203 1893 2206
rect 1898 2203 1924 2206
rect 2036 2203 2053 2206
rect 2410 2203 2429 2206
rect 2586 2203 2604 2206
rect 2626 2203 2684 2206
rect 2836 2203 2845 2206
rect 2858 2203 2908 2206
rect 2932 2203 2989 2206
rect 3314 2203 3340 2206
rect 3370 2203 3412 2206
rect 3458 2203 3485 2206
rect 3620 2203 3637 2206
rect 3642 2203 3676 2206
rect 3874 2205 3877 2213
rect 3906 2203 3932 2206
rect 3964 2203 4013 2206
rect 4068 2203 4125 2206
rect 4324 2203 4373 2206
rect 4378 2205 4381 2213
rect 4546 2203 4556 2206
rect 4588 2203 4597 2206
rect 4618 2203 4628 2206
rect 4772 2203 4781 2206
rect 666 2193 692 2196
rect 1010 2193 1044 2196
rect 2426 2193 2429 2203
rect 2818 2193 2828 2196
rect 38 2167 4829 2173
rect 1442 2143 1461 2146
rect 2706 2143 2756 2146
rect 2922 2143 2964 2146
rect 1458 2136 1461 2143
rect 188 2133 197 2136
rect 284 2133 317 2136
rect 412 2133 437 2136
rect 458 2133 468 2136
rect 484 2133 525 2136
rect 636 2133 645 2136
rect 892 2133 965 2136
rect 988 2133 1061 2136
rect 1082 2133 1116 2136
rect 116 2123 141 2126
rect 282 2123 316 2126
rect 348 2123 388 2126
rect 420 2123 429 2126
rect 492 2123 517 2126
rect 522 2123 525 2133
rect 570 2123 612 2126
rect 660 2123 669 2126
rect 850 2123 884 2126
rect 898 2123 964 2126
rect 996 2123 1021 2126
rect 1138 2123 1141 2134
rect 1346 2133 1364 2136
rect 1388 2133 1453 2136
rect 1458 2133 1468 2136
rect 1500 2133 1517 2136
rect 1708 2133 1741 2136
rect 1962 2133 2044 2136
rect 2226 2133 2252 2136
rect 1250 2123 1317 2126
rect 1380 2123 1389 2126
rect 1458 2123 1476 2126
rect 1506 2123 1548 2126
rect 1628 2123 1645 2126
rect 1682 2123 1692 2126
rect 1786 2123 1812 2126
rect 1970 2123 2036 2126
rect 2146 2123 2164 2126
rect 2282 2123 2285 2134
rect 2426 2126 2429 2134
rect 2570 2133 2620 2136
rect 2642 2133 2692 2136
rect 2764 2133 2781 2136
rect 2786 2133 2812 2136
rect 2836 2133 2885 2136
rect 2890 2126 2893 2134
rect 2978 2133 2988 2136
rect 3068 2133 3085 2136
rect 3114 2133 3124 2136
rect 3298 2126 3301 2134
rect 3354 2133 3372 2136
rect 3522 2133 3572 2136
rect 3604 2133 3645 2136
rect 3762 2133 3796 2136
rect 3828 2133 3845 2136
rect 3858 2133 3876 2136
rect 3906 2133 3924 2136
rect 4082 2126 4085 2134
rect 4106 2133 4124 2136
rect 4156 2133 4173 2136
rect 4188 2133 4197 2136
rect 4236 2133 4245 2136
rect 4284 2133 4293 2136
rect 4666 2126 4669 2134
rect 2298 2123 2348 2126
rect 2402 2123 2429 2126
rect 2554 2123 2612 2126
rect 2644 2123 2661 2126
rect 2700 2123 2749 2126
rect 2772 2123 2797 2126
rect 2802 2123 2820 2126
rect 2882 2123 2893 2126
rect 2908 2123 2933 2126
rect 3018 2123 3060 2126
rect 3284 2123 3301 2126
rect 3396 2123 3485 2126
rect 3596 2123 3629 2126
rect 3634 2123 3660 2126
rect 3690 2123 3716 2126
rect 3762 2123 3804 2126
rect 3834 2123 3884 2126
rect 3890 2123 3932 2126
rect 4076 2123 4085 2126
rect 4162 2123 4180 2126
rect 4186 2123 4228 2126
rect 4234 2123 4260 2126
rect 4466 2123 4492 2126
rect 4652 2123 4669 2126
rect 1314 2116 1317 2123
rect 2882 2116 2885 2123
rect 1140 2113 1309 2116
rect 1314 2113 1364 2116
rect 2836 2113 2885 2116
rect 3330 2113 3365 2116
rect 3402 2113 3492 2116
rect 3516 2113 3565 2116
rect 14 2067 4853 2073
rect 2314 2033 2341 2036
rect 3210 2033 3229 2036
rect 1268 2023 1349 2026
rect 1354 2016 1357 2025
rect 2796 2023 2885 2026
rect 3154 2023 3196 2026
rect 2882 2016 2885 2023
rect 116 2013 141 2016
rect 236 2013 253 2016
rect 332 2013 341 2016
rect 556 2013 604 2016
rect 634 2013 652 2016
rect 754 2013 804 2016
rect 908 2013 1037 2016
rect 1052 2013 1237 2016
rect 1338 2013 1357 2016
rect 1372 2013 1429 2016
rect 1492 2013 1517 2016
rect 1564 2013 1573 2016
rect 1714 2013 1724 2016
rect 1868 2013 1909 2016
rect 1914 2013 1932 2016
rect 1964 2013 1973 2016
rect 2044 2013 2053 2016
rect 2100 2013 2141 2016
rect 2186 2013 2276 2016
rect 1570 2006 1573 2013
rect 2138 2006 2141 2013
rect 188 2003 205 2006
rect 570 2003 596 2006
rect 676 2003 685 2006
rect 714 2003 724 2006
rect 740 2003 765 2006
rect 802 2003 812 2006
rect 828 2003 861 2006
rect 1018 2003 1044 2006
rect 1058 2003 1244 2006
rect 1268 2003 1277 2006
rect 1306 2003 1356 2006
rect 1380 2003 1461 2006
rect 1570 2003 1612 2006
rect 1876 2003 1933 2006
rect 1956 2003 1965 2006
rect 2138 2003 2156 2006
rect 2274 2003 2284 2006
rect 2306 2003 2309 2014
rect 2314 2013 2396 2016
rect 2516 2013 2557 2016
rect 2578 2013 2588 2016
rect 2740 2013 2773 2016
rect 2882 2013 2893 2016
rect 2420 2003 2437 2006
rect 2570 2003 2596 2006
rect 2612 2003 2645 2006
rect 2770 2005 2773 2013
rect 2890 2005 2893 2013
rect 2914 2013 3029 2016
rect 3060 2013 3085 2016
rect 3210 2015 3213 2033
rect 3226 2026 3229 2033
rect 3330 2033 3349 2036
rect 3226 2023 3252 2026
rect 3276 2023 3309 2026
rect 3330 2015 3333 2033
rect 3346 2026 3349 2033
rect 3346 2023 3436 2026
rect 3460 2023 3485 2026
rect 3498 2013 3508 2016
rect 3668 2013 3701 2016
rect 3740 2013 3765 2016
rect 3796 2013 3861 2016
rect 3962 2013 3972 2016
rect 4002 2013 4028 2016
rect 2914 2005 2917 2013
rect 2954 2003 2980 2006
rect 3010 2003 3036 2006
rect 3074 2003 3116 2006
rect 3148 2003 3189 2006
rect 3498 2005 3501 2013
rect 3602 2003 3644 2006
rect 4066 2003 4069 2014
rect 4106 2013 4132 2016
rect 4242 2013 4252 2016
rect 4282 2013 4308 2016
rect 4378 2013 4404 2016
rect 4092 2003 4117 2006
rect 842 1993 892 1996
rect 906 1993 1036 1996
rect 38 1967 4829 1973
rect 642 1943 676 1946
rect 978 1936 981 1946
rect 2778 1943 2836 1946
rect 204 1933 213 1936
rect 242 1926 245 1936
rect 298 1933 308 1936
rect 372 1933 413 1936
rect 564 1933 581 1936
rect 636 1933 669 1936
rect 684 1933 717 1936
rect 852 1933 885 1936
rect 948 1933 965 1936
rect 978 1933 1116 1936
rect 1324 1933 1373 1936
rect 1530 1933 1540 1936
rect 1628 1933 1645 1936
rect 1698 1933 1724 1936
rect 1852 1933 1869 1936
rect 2044 1933 2061 1936
rect 2084 1933 2165 1936
rect 2402 1933 2421 1936
rect 2602 1933 2652 1936
rect 2834 1933 2844 1936
rect 2866 1933 2900 1936
rect 2924 1933 2949 1936
rect 3306 1933 3324 1936
rect 3410 1933 3420 1936
rect 3508 1933 3557 1936
rect 3578 1933 3612 1936
rect 3722 1933 3772 1936
rect 3788 1933 3821 1936
rect 3860 1933 3901 1936
rect 3956 1933 3965 1936
rect 4332 1933 4349 1936
rect 4428 1933 4437 1936
rect 4452 1933 4461 1936
rect 4508 1933 4517 1936
rect 4522 1933 4548 1936
rect 4604 1933 4612 1936
rect 4644 1933 4661 1936
rect 4772 1933 4789 1936
rect 116 1923 141 1926
rect 178 1923 196 1926
rect 202 1923 212 1926
rect 242 1925 261 1926
rect 244 1923 261 1925
rect 266 1923 276 1926
rect 324 1923 333 1926
rect 338 1923 364 1926
rect 570 1923 612 1926
rect 692 1923 725 1926
rect 764 1923 781 1926
rect 820 1923 829 1926
rect 898 1923 924 1926
rect 1124 1923 1157 1926
rect 1282 1923 1300 1926
rect 1330 1923 1380 1926
rect 1490 1923 1500 1926
rect 1530 1923 1533 1933
rect 2418 1926 2421 1933
rect 3554 1926 3557 1933
rect 1556 1923 1612 1926
rect 1714 1923 1732 1926
rect 1812 1923 1821 1926
rect 1826 1923 1836 1926
rect 1970 1923 2020 1926
rect 2050 1923 2076 1926
rect 2252 1923 2269 1926
rect 2306 1923 2332 1926
rect 2396 1923 2413 1926
rect 2418 1923 2428 1926
rect 2458 1923 2484 1926
rect 2596 1923 2637 1926
rect 2660 1923 2677 1926
rect 2772 1923 2797 1926
rect 2852 1923 2861 1926
rect 3100 1923 3125 1926
rect 3242 1923 3268 1926
rect 3300 1923 3317 1926
rect 3444 1923 3477 1926
rect 3554 1923 3605 1926
rect 3636 1923 3692 1926
rect 3730 1923 3764 1926
rect 3874 1923 3916 1926
rect 4068 1923 4093 1926
rect 4170 1923 4188 1926
rect 4258 1923 4284 1926
rect 4324 1923 4341 1926
rect 4394 1923 4404 1926
rect 4434 1923 4444 1926
rect 4458 1923 4468 1926
rect 4586 1923 4596 1926
rect 1330 1916 1333 1923
rect 1322 1913 1333 1916
rect 2050 1913 2069 1916
rect 2866 1913 2900 1916
rect 3162 1913 3212 1916
rect 3236 1913 3253 1916
rect 3338 1913 3364 1916
rect 3388 1913 3421 1916
rect 14 1867 4853 1873
rect 3234 1833 3284 1836
rect 3298 1833 3324 1836
rect 2836 1823 2845 1826
rect 2874 1816 2877 1825
rect 2898 1823 2917 1826
rect 3002 1823 3044 1826
rect 3250 1823 3268 1826
rect 3298 1823 3308 1826
rect 3332 1823 3341 1826
rect 3372 1823 3389 1826
rect 2898 1816 2901 1823
rect 3002 1816 3005 1823
rect 124 1813 149 1816
rect 308 1813 333 1816
rect 370 1813 380 1816
rect 428 1813 453 1816
rect 196 1803 221 1806
rect 226 1803 252 1806
rect 458 1803 461 1814
rect 490 1803 493 1814
rect 564 1813 589 1816
rect 602 1813 612 1816
rect 642 1813 676 1816
rect 754 1813 780 1816
rect 858 1813 876 1816
rect 1012 1813 1061 1816
rect 1108 1813 1117 1816
rect 1164 1813 1173 1816
rect 1266 1813 1364 1816
rect 1434 1813 1460 1816
rect 1466 1813 1516 1816
rect 1546 1813 1620 1816
rect 1642 1813 1716 1816
rect 1754 1813 1764 1816
rect 1858 1813 1925 1816
rect 1962 1813 1988 1816
rect 858 1806 861 1813
rect 1170 1806 1173 1813
rect 1754 1806 1757 1813
rect 2034 1806 2037 1816
rect 2092 1813 2117 1816
rect 2122 1806 2125 1816
rect 2146 1813 2164 1816
rect 2332 1813 2349 1816
rect 2500 1813 2525 1816
rect 2570 1813 2604 1816
rect 2660 1813 2693 1816
rect 2732 1813 2741 1816
rect 2802 1813 2820 1816
rect 2834 1813 2861 1816
rect 2874 1813 2885 1816
rect 2892 1813 2901 1816
rect 2906 1813 2924 1816
rect 2994 1813 3005 1816
rect 3060 1813 3084 1816
rect 3180 1813 3189 1816
rect 3228 1813 3261 1816
rect 3412 1813 3437 1816
rect 3508 1813 3517 1816
rect 3668 1813 3693 1816
rect 3724 1813 3733 1816
rect 3762 1813 3772 1816
rect 3802 1813 3828 1816
rect 3908 1813 3917 1816
rect 3964 1813 3981 1816
rect 3996 1813 4036 1816
rect 4172 1813 4228 1816
rect 4308 1813 4325 1816
rect 4364 1813 4413 1816
rect 4420 1813 4429 1816
rect 4546 1813 4580 1816
rect 4610 1813 4636 1816
rect 498 1803 540 1806
rect 636 1803 645 1806
rect 650 1803 668 1806
rect 700 1803 717 1806
rect 740 1803 765 1806
rect 788 1803 821 1806
rect 852 1803 861 1806
rect 892 1803 901 1806
rect 978 1803 988 1806
rect 1004 1803 1053 1806
rect 1170 1803 1236 1806
rect 1268 1803 1325 1806
rect 1410 1803 1452 1806
rect 1540 1803 1565 1806
rect 1636 1803 1653 1806
rect 1666 1803 1708 1806
rect 1740 1803 1757 1806
rect 1908 1803 1933 1806
rect 2012 1803 2069 1806
rect 2122 1803 2141 1806
rect 2178 1803 2196 1806
rect 2226 1803 2252 1806
rect 2258 1803 2308 1806
rect 2338 1803 2356 1806
rect 2450 1803 2476 1806
rect 2530 1803 2540 1806
rect 2578 1803 2612 1806
rect 2634 1803 2652 1806
rect 2794 1803 2812 1806
rect 2834 1805 2837 1813
rect 2842 1803 2860 1806
rect 2874 1803 2884 1806
rect 2932 1803 2972 1806
rect 2994 1805 2997 1813
rect 3148 1803 3157 1806
rect 3178 1803 3220 1806
rect 3378 1803 3396 1806
rect 3490 1803 3500 1806
rect 3730 1805 3733 1813
rect 4004 1803 4021 1806
rect 4060 1803 4148 1806
rect 4428 1803 4445 1806
rect 218 1793 221 1803
rect 706 1793 732 1796
rect 3154 1793 3164 1796
rect 38 1767 4829 1773
rect 858 1743 892 1746
rect 1010 1743 1076 1746
rect 178 1733 212 1736
rect 276 1733 309 1736
rect 178 1723 204 1726
rect 242 1723 268 1726
rect 346 1723 349 1734
rect 386 1733 420 1736
rect 500 1733 509 1736
rect 532 1733 557 1736
rect 794 1733 836 1736
rect 900 1733 933 1736
rect 1002 1733 1084 1736
rect 1122 1733 1140 1736
rect 1322 1733 1404 1736
rect 1426 1733 1469 1736
rect 1636 1733 1701 1736
rect 1754 1733 1812 1736
rect 1828 1733 1845 1736
rect 1916 1733 1948 1736
rect 2180 1733 2205 1736
rect 2242 1733 2252 1736
rect 2266 1733 2284 1736
rect 2306 1733 2316 1736
rect 492 1723 501 1726
rect 540 1723 557 1726
rect 908 1723 957 1726
rect 1004 1723 1021 1726
rect 1092 1723 1101 1726
rect 1114 1723 1148 1726
rect 1178 1723 1204 1726
rect 1250 1723 1292 1726
rect 1426 1725 1429 1733
rect 1842 1726 1845 1733
rect 1434 1723 1612 1726
rect 1690 1723 1708 1726
rect 1842 1723 1892 1726
rect 1978 1723 2012 1726
rect 2042 1723 2084 1726
rect 2202 1725 2205 1733
rect 2474 1726 2477 1745
rect 2820 1743 2845 1746
rect 3010 1743 3020 1746
rect 3090 1743 3116 1746
rect 2602 1733 2628 1736
rect 2786 1726 2789 1734
rect 3042 1733 3076 1736
rect 3114 1726 3117 1736
rect 3124 1733 3157 1736
rect 2452 1723 2477 1726
rect 2610 1723 2669 1726
rect 2610 1716 2613 1723
rect 1314 1713 1341 1716
rect 2506 1713 2524 1716
rect 2554 1713 2572 1716
rect 2596 1713 2613 1716
rect 2666 1716 2669 1723
rect 2778 1723 2789 1726
rect 2890 1723 2916 1726
rect 2922 1723 2948 1726
rect 2978 1723 2996 1726
rect 3042 1723 3117 1726
rect 3362 1723 3380 1726
rect 3394 1723 3397 1734
rect 3434 1723 3452 1726
rect 3458 1723 3468 1726
rect 3474 1723 3477 1734
rect 3642 1726 3645 1734
rect 3666 1733 3684 1736
rect 3756 1733 3765 1736
rect 3812 1733 3829 1736
rect 3850 1733 3860 1736
rect 4340 1733 4389 1736
rect 4434 1733 4452 1736
rect 4532 1733 4541 1736
rect 4604 1733 4613 1736
rect 4626 1733 4636 1736
rect 4668 1733 4765 1736
rect 3818 1726 3821 1733
rect 4610 1726 4613 1733
rect 3572 1723 3597 1726
rect 3628 1723 3645 1726
rect 3652 1723 3692 1726
rect 3738 1723 3788 1726
rect 3818 1723 3844 1726
rect 3858 1723 3868 1726
rect 3898 1723 3908 1726
rect 3938 1723 3972 1726
rect 4108 1723 4117 1726
rect 4244 1723 4253 1726
rect 4346 1723 4412 1726
rect 4514 1723 4524 1726
rect 4530 1723 4580 1726
rect 4610 1723 4644 1726
rect 2778 1716 2781 1723
rect 2666 1713 2684 1716
rect 2714 1713 2748 1716
rect 2772 1713 2781 1716
rect 2826 1713 2860 1716
rect 2884 1713 2901 1716
rect 3138 1713 3164 1716
rect 3210 1713 3228 1716
rect 3322 1713 3332 1716
rect 3356 1713 3373 1716
rect 2642 1703 2700 1706
rect 2722 1703 2764 1706
rect 2868 1703 2909 1706
rect 3258 1703 3348 1706
rect 14 1667 4853 1673
rect 2698 1653 2733 1656
rect 2866 1633 2916 1636
rect 3234 1633 3268 1636
rect 2882 1623 2900 1626
rect 2924 1623 3012 1626
rect 2882 1616 2885 1623
rect 114 1613 124 1616
rect 146 1613 164 1616
rect 236 1613 245 1616
rect 292 1613 301 1616
rect 306 1613 316 1616
rect 348 1614 357 1616
rect 346 1613 357 1614
rect 604 1613 621 1616
rect 626 1613 676 1616
rect 948 1613 1013 1616
rect 1028 1613 1093 1616
rect 1132 1613 1181 1616
rect 1252 1613 1261 1616
rect 1378 1613 1436 1616
rect 1530 1613 1556 1616
rect 1706 1613 1716 1616
rect 132 1603 165 1606
rect 346 1603 349 1613
rect 610 1603 668 1606
rect 706 1603 812 1606
rect 828 1603 861 1606
rect 940 1603 965 1606
rect 1020 1603 1037 1606
rect 1098 1603 1108 1606
rect 1124 1603 1165 1606
rect 1260 1603 1301 1606
rect 1322 1603 1348 1606
rect 1378 1605 1381 1613
rect 1530 1603 1548 1606
rect 1714 1603 1724 1606
rect 1746 1603 1749 1614
rect 1754 1613 1788 1616
rect 1954 1613 1980 1616
rect 2036 1613 2060 1616
rect 2130 1613 2156 1616
rect 2234 1613 2260 1616
rect 2410 1613 2420 1616
rect 2466 1613 2476 1616
rect 2802 1613 2828 1616
rect 2842 1613 2885 1616
rect 3084 1613 3101 1616
rect 3212 1613 3237 1616
rect 3298 1613 3332 1616
rect 3356 1613 3365 1616
rect 3370 1613 3388 1616
rect 3444 1613 3453 1616
rect 1890 1603 1916 1606
rect 2010 1603 2020 1606
rect 2522 1603 2532 1606
rect 2714 1603 2836 1606
rect 842 1593 932 1596
rect 954 1593 1012 1596
rect 2842 1595 2845 1613
rect 3042 1603 3076 1606
rect 3220 1603 3245 1606
rect 3330 1595 3333 1606
rect 3370 1603 3373 1613
rect 3570 1607 3573 1616
rect 3578 1607 3581 1616
rect 3588 1613 3605 1616
rect 3636 1613 3709 1616
rect 3746 1613 3788 1616
rect 3898 1613 3916 1616
rect 3922 1613 3948 1616
rect 3978 1613 4012 1616
rect 4116 1613 4149 1616
rect 4258 1613 4292 1616
rect 4322 1613 4372 1616
rect 4418 1613 4436 1616
rect 4532 1613 4588 1616
rect 4716 1613 4733 1616
rect 3706 1607 3709 1613
rect 4146 1607 4149 1613
rect 3660 1603 3677 1606
rect 3754 1603 3780 1606
rect 3818 1603 3844 1606
rect 3924 1603 3933 1606
rect 3972 1603 3997 1606
rect 4042 1603 4052 1606
rect 4180 1603 4220 1606
rect 4330 1603 4364 1606
rect 4460 1603 4508 1606
rect 4540 1603 4565 1606
rect 4612 1603 4677 1606
rect 3402 1593 3420 1596
rect 4674 1593 4677 1603
rect 38 1567 4829 1573
rect 308 1533 317 1536
rect 108 1523 133 1526
rect 164 1523 197 1526
rect 236 1523 261 1526
rect 306 1523 316 1526
rect 346 1525 349 1536
rect 354 1533 388 1536
rect 506 1526 509 1546
rect 1098 1536 1101 1556
rect 3204 1543 3213 1546
rect 514 1533 524 1536
rect 540 1533 549 1536
rect 682 1533 708 1536
rect 740 1533 757 1536
rect 812 1533 821 1536
rect 850 1526 853 1536
rect 892 1533 901 1536
rect 1068 1533 1077 1536
rect 1098 1533 1148 1536
rect 1226 1533 1260 1536
rect 1434 1533 1476 1536
rect 1660 1533 1733 1536
rect 1778 1533 1836 1536
rect 1874 1533 1884 1536
rect 1930 1533 1956 1536
rect 1978 1533 1997 1536
rect 2332 1533 2341 1536
rect 3050 1533 3092 1536
rect 3106 1533 3124 1536
rect 3202 1533 3228 1536
rect 3242 1533 3276 1536
rect 3330 1533 3348 1536
rect 3380 1533 3405 1536
rect 3572 1533 3581 1536
rect 3690 1533 3708 1536
rect 3740 1533 3749 1536
rect 3754 1533 3788 1536
rect 3812 1533 3837 1536
rect 3922 1533 3964 1536
rect 3988 1533 4013 1536
rect 4028 1533 4061 1536
rect 4122 1533 4140 1536
rect 4188 1533 4221 1536
rect 4252 1533 4277 1536
rect 4322 1533 4340 1536
rect 4394 1533 4428 1536
rect 4458 1533 4484 1536
rect 4508 1533 4517 1536
rect 412 1523 421 1526
rect 426 1523 460 1526
rect 484 1523 493 1526
rect 506 1523 516 1526
rect 548 1523 557 1526
rect 676 1523 701 1526
rect 706 1523 716 1526
rect 746 1523 788 1526
rect 820 1523 837 1526
rect 850 1523 876 1526
rect 972 1523 997 1526
rect 1034 1523 1060 1526
rect 1082 1523 1140 1526
rect 1172 1523 1252 1526
rect 1298 1523 1340 1526
rect 1442 1523 1468 1526
rect 1580 1523 1605 1526
rect 1642 1523 1652 1526
rect 1706 1523 1740 1526
rect 1772 1523 1837 1526
rect 1850 1523 1876 1526
rect 1922 1523 1948 1526
rect 1978 1525 1981 1533
rect 1986 1523 2068 1526
rect 2164 1523 2173 1526
rect 2266 1523 2316 1526
rect 2338 1523 2388 1526
rect 2458 1523 2484 1526
rect 2644 1523 2700 1526
rect 2922 1523 2925 1533
rect 3050 1526 3053 1533
rect 3028 1523 3053 1526
rect 3108 1523 3117 1526
rect 3122 1523 3132 1526
rect 3170 1523 3180 1526
rect 3210 1523 3236 1526
rect 3306 1523 3356 1526
rect 3620 1523 3629 1526
rect 3682 1523 3716 1526
rect 3882 1523 3900 1526
rect 3954 1523 3972 1526
rect 3170 1516 3173 1523
rect 2260 1513 2277 1516
rect 2924 1513 2933 1516
rect 3148 1513 3173 1516
rect 3244 1513 3269 1516
rect 4010 1515 4013 1533
rect 4066 1523 4084 1526
rect 4114 1523 4117 1533
rect 4162 1526 4165 1533
rect 4162 1523 4173 1526
rect 4186 1523 4228 1526
rect 4234 1523 4244 1526
rect 4250 1523 4253 1533
rect 4450 1526 4453 1533
rect 4522 1526 4525 1536
rect 4530 1533 4556 1536
rect 4586 1533 4644 1536
rect 4676 1533 4685 1536
rect 4748 1533 4765 1536
rect 4356 1523 4373 1526
rect 4450 1523 4477 1526
rect 4500 1523 4525 1526
rect 4578 1523 4581 1533
rect 4682 1526 4685 1533
rect 4762 1526 4765 1533
rect 4626 1523 4652 1526
rect 4682 1523 4724 1526
rect 4762 1523 4780 1526
rect 4170 1515 4173 1523
rect 4186 1513 4220 1516
rect 4322 1513 4340 1516
rect 4394 1513 4428 1516
rect 4458 1513 4484 1516
rect 4522 1513 4556 1516
rect 1914 1503 1933 1506
rect 2226 1503 2252 1506
rect 3300 1503 3325 1506
rect 14 1467 4853 1473
rect 738 1423 757 1426
rect 738 1416 741 1423
rect 818 1416 821 1426
rect 3244 1423 3253 1426
rect 3908 1423 3917 1426
rect 4106 1423 4148 1426
rect 260 1413 269 1416
rect 434 1413 444 1416
rect 450 1413 508 1416
rect 540 1413 565 1416
rect 676 1413 701 1416
rect 732 1413 741 1416
rect 746 1413 764 1416
rect 794 1413 828 1416
rect 948 1413 1005 1416
rect 1020 1413 1037 1416
rect 1148 1413 1157 1416
rect 1196 1413 1221 1416
rect 1258 1413 1292 1416
rect 1506 1413 1556 1416
rect 1604 1413 1629 1416
rect 1844 1413 1869 1416
rect 1900 1413 1909 1416
rect 2010 1413 2020 1416
rect 2050 1413 2068 1416
rect 2106 1413 2124 1416
rect 2212 1413 2229 1416
rect 2268 1413 2325 1416
rect 2588 1413 2629 1416
rect 2658 1413 2668 1416
rect 2762 1413 2780 1416
rect 3010 1413 3052 1416
rect 3076 1413 3085 1416
rect 3242 1413 3260 1416
rect 3266 1413 3300 1416
rect 3324 1413 3397 1416
rect 3402 1413 3412 1416
rect 3436 1413 3541 1416
rect 3716 1413 3725 1416
rect 3772 1413 3781 1416
rect 3786 1413 3796 1416
rect 3818 1413 3844 1416
rect 3858 1413 3892 1416
rect 3972 1413 3981 1416
rect 4028 1413 4037 1416
rect 4042 1413 4100 1416
rect 4164 1413 4205 1416
rect 4244 1413 4269 1416
rect 4300 1413 4317 1416
rect 4396 1413 4437 1416
rect 4596 1413 4621 1416
rect 4660 1413 4677 1416
rect 4314 1407 4317 1413
rect 186 1403 196 1406
rect 212 1403 221 1406
rect 378 1403 396 1406
rect 452 1403 485 1406
rect 490 1403 516 1406
rect 546 1403 572 1406
rect 772 1403 805 1406
rect 818 1403 836 1406
rect 914 1403 940 1406
rect 994 1403 1012 1406
rect 1266 1403 1284 1406
rect 1434 1403 1476 1406
rect 1676 1403 1733 1406
rect 2596 1403 2605 1406
rect 2762 1403 2772 1406
rect 3004 1403 3053 1406
rect 3130 1403 3228 1406
rect 3268 1403 3293 1406
rect 490 1396 493 1403
rect 474 1393 493 1396
rect 866 1393 932 1396
rect 954 1393 1004 1396
rect 3076 1393 3093 1396
rect 3298 1395 3301 1406
rect 3316 1403 3349 1406
rect 3812 1403 3821 1406
rect 3852 1403 3877 1406
rect 4108 1403 4141 1406
rect 4172 1403 4181 1406
rect 4354 1403 4372 1406
rect 4404 1403 4421 1406
rect 3330 1393 3412 1396
rect 38 1367 4829 1373
rect 858 1343 892 1346
rect 906 1343 964 1346
rect 2554 1336 2557 1344
rect 3108 1343 3117 1346
rect 3322 1343 3348 1346
rect 148 1333 181 1336
rect 298 1333 317 1336
rect 340 1333 365 1336
rect 106 1323 140 1326
rect 220 1323 229 1326
rect 276 1323 285 1326
rect 292 1323 309 1326
rect 314 1325 317 1333
rect 404 1323 429 1326
rect 466 1325 469 1336
rect 514 1333 540 1336
rect 570 1333 596 1336
rect 628 1333 661 1336
rect 780 1333 805 1336
rect 818 1333 828 1336
rect 844 1333 869 1336
rect 900 1333 933 1336
rect 972 1333 981 1336
rect 506 1323 532 1326
rect 578 1323 604 1326
rect 700 1323 725 1326
rect 762 1323 772 1326
rect 794 1323 820 1326
rect 908 1323 965 1326
rect 980 1323 1037 1326
rect 1068 1323 1093 1326
rect 1122 1325 1125 1336
rect 1148 1333 1157 1336
rect 1162 1333 1244 1336
rect 1266 1333 1316 1336
rect 1354 1333 1364 1336
rect 1436 1333 1477 1336
rect 1156 1323 1165 1326
rect 1218 1323 1236 1326
rect 1466 1323 1476 1326
rect 1506 1325 1509 1336
rect 1522 1333 1540 1336
rect 1572 1333 1581 1336
rect 1628 1333 1653 1336
rect 1658 1333 1684 1336
rect 1716 1333 1749 1336
rect 1772 1333 1781 1336
rect 1786 1333 1804 1336
rect 2452 1333 2469 1336
rect 2498 1333 2540 1336
rect 2554 1333 2573 1336
rect 2596 1333 2605 1336
rect 2674 1333 2692 1336
rect 2850 1333 2860 1336
rect 3082 1333 3092 1336
rect 3146 1333 3164 1336
rect 3188 1333 3213 1336
rect 3266 1333 3284 1336
rect 3300 1333 3317 1336
rect 3370 1333 3396 1336
rect 3508 1333 3517 1336
rect 3540 1333 3565 1336
rect 3674 1333 3708 1336
rect 3844 1333 3957 1336
rect 3996 1333 4029 1336
rect 4282 1333 4316 1336
rect 4348 1333 4357 1336
rect 4388 1333 4397 1336
rect 4498 1333 4508 1336
rect 4538 1333 4564 1336
rect 4602 1333 4613 1336
rect 4652 1333 4693 1336
rect 4772 1333 4789 1336
rect 2570 1326 2573 1333
rect 3266 1326 3269 1333
rect 1564 1323 1604 1326
rect 1634 1323 1692 1326
rect 1738 1323 1748 1326
rect 1780 1323 1805 1326
rect 1812 1323 1821 1326
rect 1858 1323 1884 1326
rect 1930 1323 1996 1326
rect 2034 1323 2052 1326
rect 1962 1313 1965 1323
rect 2114 1306 2117 1325
rect 2204 1323 2213 1326
rect 2274 1323 2284 1326
rect 2426 1323 2444 1326
rect 2474 1323 2532 1326
rect 2570 1323 2588 1326
rect 2666 1323 2684 1326
rect 2716 1323 2748 1326
rect 2842 1323 2868 1326
rect 2988 1323 3037 1326
rect 3180 1323 3269 1326
rect 3314 1323 3348 1326
rect 3372 1323 3404 1326
rect 3514 1323 3524 1326
rect 3562 1323 3565 1333
rect 3570 1323 3573 1333
rect 3610 1323 3668 1326
rect 3706 1323 3709 1333
rect 4162 1326 4165 1333
rect 4602 1326 4605 1333
rect 3746 1323 3788 1326
rect 3794 1323 3836 1326
rect 3988 1323 4029 1326
rect 4068 1323 4156 1326
rect 4162 1323 4188 1326
rect 4226 1323 4244 1326
rect 4354 1323 4380 1326
rect 4524 1323 4557 1326
rect 4580 1323 4605 1326
rect 4610 1323 4628 1326
rect 4666 1323 4708 1326
rect 4738 1323 4764 1326
rect 2426 1316 2429 1323
rect 2124 1313 2165 1316
rect 2412 1313 2429 1316
rect 2996 1313 3037 1316
rect 3154 1313 3164 1316
rect 3818 1313 3828 1316
rect 2114 1303 2133 1306
rect 3052 1303 3077 1306
rect 14 1267 4853 1273
rect 2124 1233 2141 1236
rect 3092 1233 3109 1236
rect 2042 1223 2116 1226
rect 2130 1223 2140 1226
rect 2346 1223 2380 1226
rect 3050 1223 3084 1226
rect 3108 1223 3117 1226
rect 3884 1223 3909 1226
rect 2346 1216 2349 1223
rect 108 1213 133 1216
rect 178 1213 188 1216
rect 218 1206 221 1214
rect 226 1213 260 1216
rect 266 1213 276 1216
rect 308 1213 349 1216
rect 418 1213 428 1216
rect 434 1213 460 1216
rect 492 1213 501 1216
rect 682 1213 716 1216
rect 746 1213 772 1216
rect 858 1213 884 1216
rect 972 1213 997 1216
rect 1052 1213 1077 1216
rect 1108 1213 1157 1216
rect 1162 1213 1204 1216
rect 1540 1213 1557 1216
rect 1564 1213 1573 1216
rect 1610 1213 1636 1216
rect 1770 1213 1788 1216
rect 1890 1213 1940 1216
rect 1972 1213 2013 1216
rect 1154 1206 1157 1213
rect 1770 1206 1773 1213
rect 180 1203 189 1206
rect 218 1203 253 1206
rect 268 1203 277 1206
rect 300 1203 348 1206
rect 436 1203 461 1206
rect 626 1203 644 1206
rect 676 1203 685 1206
rect 698 1203 708 1206
rect 740 1203 757 1206
rect 780 1203 797 1206
rect 802 1203 812 1206
rect 828 1203 837 1206
rect 842 1203 892 1206
rect 964 1203 973 1206
rect 1154 1203 1212 1206
rect 1234 1203 1316 1206
rect 1348 1203 1373 1206
rect 1490 1203 1516 1206
rect 1546 1203 1556 1206
rect 1756 1203 1773 1206
rect 1970 1203 2028 1206
rect 2130 1203 2133 1214
rect 2252 1213 2277 1216
rect 2308 1213 2317 1216
rect 2324 1213 2349 1216
rect 2522 1213 2532 1216
rect 2538 1213 2581 1216
rect 2634 1213 2653 1216
rect 3028 1213 3077 1216
rect 3172 1213 3229 1216
rect 2314 1207 2317 1213
rect 2522 1206 2525 1213
rect 2650 1207 2653 1213
rect 2180 1203 2205 1206
rect 2346 1203 2380 1206
rect 2404 1203 2413 1206
rect 2506 1203 2525 1206
rect 2540 1203 2581 1206
rect 2586 1203 2604 1206
rect 2754 1203 2764 1206
rect 2882 1203 2900 1206
rect 3122 1203 3156 1206
rect 3180 1203 3189 1206
rect 3210 1203 3228 1206
rect 3242 1203 3245 1214
rect 3276 1213 3309 1216
rect 3340 1213 3349 1216
rect 3716 1213 3741 1216
rect 3772 1213 3781 1216
rect 3802 1213 3820 1216
rect 3850 1213 3876 1216
rect 4026 1213 4044 1216
rect 4050 1207 4053 1216
rect 4220 1213 4237 1216
rect 4276 1213 4301 1216
rect 4308 1213 4325 1216
rect 4388 1213 4469 1216
rect 4580 1213 4589 1216
rect 4594 1213 4628 1216
rect 3268 1203 3301 1206
rect 922 1193 956 1196
rect 970 1193 996 1196
rect 2506 1195 2509 1203
rect 2586 1196 2589 1203
rect 2570 1193 2589 1196
rect 3314 1195 3317 1206
rect 3636 1203 3677 1206
rect 3794 1203 3812 1206
rect 4330 1203 4364 1206
rect 4460 1203 4493 1206
rect 4532 1203 4541 1206
rect 4546 1203 4564 1206
rect 4588 1203 4605 1206
rect 38 1167 4829 1173
rect 906 1143 932 1146
rect 946 1143 1060 1146
rect 3146 1143 3164 1146
rect 570 1133 580 1136
rect 892 1133 901 1136
rect 1068 1133 1109 1136
rect 1148 1133 1221 1136
rect 1404 1133 1437 1136
rect 1460 1133 1469 1136
rect 1724 1133 1749 1136
rect 1772 1133 1829 1136
rect 1986 1133 2028 1136
rect 2410 1133 2420 1136
rect 2532 1133 2541 1136
rect 2730 1133 2748 1136
rect 2866 1133 2892 1136
rect 3010 1133 3020 1136
rect 3066 1133 3084 1136
rect 3132 1133 3141 1136
rect 3252 1133 3261 1136
rect 3282 1133 3308 1136
rect 3330 1133 3348 1136
rect 3578 1133 3588 1136
rect 3666 1133 3676 1136
rect 3772 1133 3781 1136
rect 3794 1133 3900 1136
rect 3980 1133 4021 1136
rect 4140 1133 4165 1136
rect 4194 1133 4220 1136
rect 4252 1133 4285 1136
rect 4298 1133 4308 1136
rect 4420 1133 4453 1136
rect 4466 1133 4476 1136
rect 4538 1133 4556 1136
rect 4626 1133 4636 1136
rect 4674 1133 4684 1136
rect 4764 1133 4781 1136
rect 3330 1126 3333 1133
rect 164 1123 173 1126
rect 228 1123 237 1126
rect 284 1123 309 1126
rect 508 1123 533 1126
rect 610 1123 628 1126
rect 762 1123 772 1126
rect 818 1123 828 1126
rect 866 1123 884 1126
rect 948 1123 1061 1126
rect 1082 1123 1140 1126
rect 1316 1123 1341 1126
rect 1386 1123 1396 1126
rect 1418 1123 1436 1126
rect 1482 1123 1492 1126
rect 1530 1123 1548 1126
rect 1628 1123 1653 1126
rect 1690 1123 1716 1126
rect 1722 1123 1748 1126
rect 1850 1123 1892 1126
rect 2010 1123 2020 1126
rect 2058 1123 2076 1126
rect 2170 1113 2204 1116
rect 2210 1106 2213 1125
rect 2234 1123 2284 1126
rect 2330 1123 2340 1126
rect 2586 1123 2596 1126
rect 2730 1123 2756 1126
rect 2874 1123 2900 1126
rect 3028 1123 3085 1126
rect 3092 1123 3109 1126
rect 3130 1123 3164 1126
rect 3194 1123 3228 1126
rect 3260 1123 3309 1126
rect 3316 1123 3333 1126
rect 3372 1123 3389 1126
rect 3532 1123 3541 1126
rect 3548 1123 3589 1126
rect 3730 1123 3805 1126
rect 3938 1123 3972 1126
rect 4068 1123 4132 1126
rect 4258 1123 4316 1126
rect 4354 1123 4396 1126
rect 4426 1123 4484 1126
rect 4594 1123 4644 1126
rect 4674 1123 4692 1126
rect 4722 1123 4756 1126
rect 2228 1113 2277 1116
rect 3098 1113 3108 1116
rect 2194 1103 2213 1106
rect 14 1067 4853 1073
rect 3074 1033 3093 1036
rect 2322 1016 2325 1025
rect 2354 1023 2364 1026
rect 2386 1016 2389 1025
rect 3028 1023 3037 1026
rect 3074 1016 3077 1033
rect 124 1013 149 1016
rect 154 1013 164 1016
rect 196 1013 229 1016
rect 234 1013 244 1016
rect 250 1013 284 1016
rect 428 1013 445 1016
rect 540 1013 549 1016
rect 634 1013 676 1016
rect 722 1013 748 1016
rect 842 1013 860 1016
rect 866 1013 892 1016
rect 1012 1013 1125 1016
rect 1140 1013 1197 1016
rect 1228 1013 1237 1016
rect 1330 1013 1364 1016
rect 1452 1013 1509 1016
rect 1524 1013 1533 1016
rect 1580 1013 1589 1016
rect 1594 1013 1620 1016
rect 1674 1013 1740 1016
rect 1786 1013 1797 1016
rect 1802 1013 1820 1016
rect 1858 1013 1884 1016
rect 1978 1013 1996 1016
rect 2010 1013 2020 1016
rect 2058 1013 2084 1016
rect 2114 1013 2172 1016
rect 2194 1013 2228 1016
rect 2268 1013 2301 1016
rect 2308 1013 2325 1016
rect 2340 1013 2349 1016
rect 2372 1013 2389 1016
rect 2410 1013 2452 1016
rect 2476 1013 2509 1016
rect 2540 1013 2549 1016
rect 2572 1013 2620 1016
rect 2652 1013 2677 1016
rect 2690 1013 2716 1016
rect 2818 1013 2836 1016
rect 3020 1013 3045 1016
rect 3052 1013 3077 1016
rect 3090 1015 3093 1033
rect 3114 1023 3164 1026
rect 3834 1023 3844 1026
rect 4306 1023 4372 1026
rect 4442 1023 4524 1026
rect 4610 1023 4636 1026
rect 3180 1013 3212 1016
rect 3250 1013 3268 1016
rect 3300 1013 3404 1016
rect 3594 1013 3668 1016
rect 3706 1013 3796 1016
rect 3826 1013 3852 1016
rect 4026 1013 4076 1016
rect 634 1006 637 1013
rect 722 1006 725 1013
rect 1794 1006 1797 1013
rect 2410 1007 2413 1013
rect 2546 1007 2549 1013
rect 4226 1007 4229 1016
rect 4388 1013 4405 1016
rect 4428 1013 4517 1016
rect 4540 1013 4549 1016
rect 116 1003 133 1006
rect 252 1003 285 1006
rect 308 1003 348 1006
rect 628 1003 637 1006
rect 642 1003 668 1006
rect 700 1003 725 1006
rect 868 1003 885 1006
rect 986 1003 1004 1006
rect 1114 1003 1132 1006
rect 1154 1003 1204 1006
rect 1236 1003 1253 1006
rect 1372 1003 1421 1006
rect 1490 1003 1516 1006
rect 1764 1003 1789 1006
rect 1794 1003 1828 1006
rect 2004 1003 2021 1006
rect 2044 1003 2069 1006
rect 2180 1003 2221 1006
rect 2236 1003 2253 1006
rect 2274 1003 2300 1006
rect 2314 1003 2324 1006
rect 2348 1003 2365 1006
rect 930 993 996 996
rect 1010 993 1124 996
rect 2450 995 2453 1006
rect 2596 1003 2605 1006
rect 2610 1003 2628 1006
rect 2810 1003 2828 1006
rect 2946 1003 3012 1006
rect 3026 1003 3044 1006
rect 3154 1003 3164 1006
rect 3188 1003 3197 1006
rect 3234 1003 3276 1006
rect 3298 1003 3396 1006
rect 3692 1003 3733 1006
rect 3738 1003 3788 1006
rect 3860 1003 3901 1006
rect 3940 1003 3965 1006
rect 3970 1003 3988 1006
rect 4100 1003 4148 1006
rect 4266 1003 4372 1006
rect 4396 1003 4405 1006
rect 4436 1003 4445 1006
rect 4450 1003 4524 1006
rect 4596 1003 4621 1006
rect 4660 1003 4677 1006
rect 38 967 4829 973
rect 2482 936 2485 944
rect 130 933 164 936
rect 284 933 309 936
rect 346 933 356 936
rect 452 933 461 936
rect 564 933 573 936
rect 754 933 780 936
rect 812 933 821 936
rect 852 933 885 936
rect 1068 933 1125 936
rect 1244 933 1269 936
rect 1370 933 1388 936
rect 1426 933 1484 936
rect 1506 926 1509 936
rect 1748 933 1765 936
rect 2042 933 2052 936
rect 2130 933 2172 936
rect 2482 933 2493 936
rect 2610 933 2628 936
rect 2994 933 3020 936
rect 3172 933 3181 936
rect 3218 933 3284 936
rect 3300 933 3309 936
rect 154 923 172 926
rect 212 923 237 926
rect 298 923 308 926
rect 354 923 364 926
rect 394 923 428 926
rect 492 923 517 926
rect 546 923 556 926
rect 692 923 717 926
rect 748 923 781 926
rect 818 923 828 926
rect 972 923 997 926
rect 1034 923 1060 926
rect 1074 923 1124 926
rect 1156 923 1165 926
rect 1250 923 1276 926
rect 1412 923 1469 926
rect 1506 925 1525 926
rect 1508 923 1525 925
rect 1650 923 1676 926
rect 1708 923 1725 926
rect 1740 923 1757 926
rect 1834 923 1860 926
rect 2130 916 2133 933
rect 2490 926 2493 933
rect 2154 923 2197 926
rect 2236 923 2261 926
rect 2306 923 2324 926
rect 2450 923 2460 926
rect 2490 923 2524 926
rect 2564 923 2620 926
rect 2754 923 2772 926
rect 3028 923 3077 926
rect 2082 913 2100 916
rect 2124 913 2133 916
rect 2332 913 2357 916
rect 3036 913 3053 916
rect 3074 906 3077 923
rect 3090 906 3093 925
rect 3114 923 3156 926
rect 3218 923 3221 933
rect 3338 926 3341 936
rect 3482 933 3508 936
rect 3628 933 3645 936
rect 3676 933 3693 936
rect 3740 933 3757 936
rect 3778 933 3788 936
rect 3812 933 3837 936
rect 3922 933 3932 936
rect 4020 933 4061 936
rect 4186 933 4220 936
rect 4250 933 4308 936
rect 4338 933 4412 936
rect 4450 933 4476 936
rect 4500 933 4517 936
rect 3954 926 3957 933
rect 4154 926 4157 933
rect 3226 923 3276 926
rect 3308 923 3317 926
rect 3322 923 3348 926
rect 3380 923 3461 926
rect 3490 923 3516 926
rect 3548 923 3573 926
rect 3698 923 3732 926
rect 3810 923 3868 926
rect 3914 923 3940 926
rect 3954 923 3965 926
rect 3970 923 4012 926
rect 4098 923 4140 926
rect 4146 923 4157 926
rect 4178 926 4181 933
rect 4178 923 4205 926
rect 4428 923 4469 926
rect 4492 923 4557 926
rect 3962 916 3965 923
rect 3108 913 3141 916
rect 3562 913 3580 916
rect 3634 913 3652 916
rect 3682 913 3724 916
rect 3812 913 3853 916
rect 3876 913 3893 916
rect 3962 913 4004 916
rect 4026 913 4068 916
rect 4146 915 4149 923
rect 4354 913 4412 916
rect 4450 913 4476 916
rect 3074 903 3093 906
rect 14 867 4853 873
rect 2154 833 2180 836
rect 2106 823 2124 826
rect 3028 823 3037 826
rect 3050 823 3068 826
rect 3948 823 3997 826
rect 4074 823 4084 826
rect 3050 816 3053 823
rect 3994 816 3997 823
rect 108 813 117 816
rect 300 813 317 816
rect 364 813 389 816
rect 420 813 453 816
rect 492 814 532 816
rect 450 806 453 813
rect 490 813 532 814
rect 628 813 637 816
rect 666 813 684 816
rect 714 813 724 816
rect 450 803 468 806
rect 490 803 493 813
rect 666 806 669 813
rect 842 806 845 816
rect 866 813 876 816
rect 914 813 940 816
rect 1004 813 1045 816
rect 1068 813 1093 816
rect 1108 813 1117 816
rect 1156 813 1181 816
rect 1258 813 1276 816
rect 1290 813 1324 816
rect 1362 813 1372 816
rect 1530 813 1548 816
rect 1666 813 1684 816
rect 1714 813 1740 816
rect 1778 813 1796 816
rect 556 803 565 806
rect 594 803 604 806
rect 660 803 669 806
rect 708 803 717 806
rect 732 803 741 806
rect 786 803 804 806
rect 820 803 837 806
rect 842 803 868 806
rect 978 803 996 806
rect 1050 803 1060 806
rect 1100 803 1109 806
rect 1218 803 1228 806
rect 1298 803 1332 806
rect 1354 803 1364 806
rect 1522 803 1540 806
rect 1612 803 1637 806
rect 1708 803 1733 806
rect 1748 803 1773 806
rect 1802 803 1812 806
rect 1834 803 1837 814
rect 1874 813 1900 816
rect 1972 813 2029 816
rect 2194 813 2236 816
rect 2260 813 2285 816
rect 2338 807 2341 816
rect 2490 813 2524 816
rect 2530 813 2548 816
rect 2580 813 2620 816
rect 2730 813 2740 816
rect 2850 813 2884 816
rect 3020 813 3053 816
rect 3130 813 3172 816
rect 3186 813 3212 816
rect 3298 813 3324 816
rect 3356 813 3365 816
rect 3548 813 3597 816
rect 3620 813 3645 816
rect 3762 813 3868 816
rect 3898 813 3940 816
rect 3994 813 4005 816
rect 4026 813 4092 816
rect 4162 813 4172 816
rect 4234 813 4284 816
rect 4346 813 4356 816
rect 4530 813 4556 816
rect 4658 813 4716 816
rect 4722 813 4773 816
rect 2490 806 2493 813
rect 3130 806 3133 813
rect 3594 807 3597 813
rect 4002 807 4005 813
rect 4658 807 4661 813
rect 4722 807 4725 813
rect 1938 803 1948 806
rect 1964 803 2037 806
rect 2290 803 2308 806
rect 2482 803 2493 806
rect 2532 803 2541 806
rect 2572 803 2589 806
rect 2714 803 2732 806
rect 2844 803 2869 806
rect 2994 803 3012 806
rect 3116 803 3133 806
rect 3236 803 3309 806
rect 3490 803 3524 806
rect 3626 803 3652 806
rect 3684 803 3724 806
rect 3850 803 3860 806
rect 3884 803 3893 806
rect 4100 803 4149 806
rect 4154 803 4164 806
rect 4314 803 4348 806
rect 4442 803 4476 806
rect 4580 803 4628 806
rect 978 793 988 796
rect 1002 793 1052 796
rect 1074 793 1092 796
rect 2482 795 2485 803
rect 3258 783 3293 786
rect 38 767 4829 773
rect 1010 743 1028 746
rect 180 733 189 736
rect 194 733 204 736
rect 260 733 293 736
rect 108 723 133 726
rect 178 723 196 726
rect 228 723 236 726
rect 268 723 308 726
rect 354 723 388 726
rect 418 725 421 736
rect 426 733 436 736
rect 810 733 820 736
rect 850 733 884 736
rect 1036 733 1069 736
rect 1178 733 1204 736
rect 1220 733 1268 736
rect 1300 733 1325 736
rect 1426 733 1460 736
rect 1490 733 1508 736
rect 1892 733 1909 736
rect 2460 733 2469 736
rect 2474 733 2532 736
rect 2538 733 2564 736
rect 2818 733 2828 736
rect 2994 733 3020 736
rect 3042 733 3068 736
rect 3220 733 3245 736
rect 3276 733 3317 736
rect 1906 726 1909 733
rect 2538 726 2541 733
rect 3466 726 3469 736
rect 3514 733 3532 736
rect 3562 733 3596 736
rect 3698 733 3724 736
rect 3828 733 3868 736
rect 3978 733 4020 736
rect 4124 733 4197 736
rect 4266 733 4276 736
rect 4476 733 4485 736
rect 4546 733 4580 736
rect 4684 733 4716 736
rect 444 723 453 726
rect 508 723 533 726
rect 570 723 580 726
rect 684 723 693 726
rect 892 723 909 726
rect 946 723 972 726
rect 1044 723 1077 726
rect 1116 723 1141 726
rect 1172 723 1189 726
rect 1292 723 1301 726
rect 1516 723 1533 726
rect 1570 723 1596 726
rect 1684 723 1709 726
rect 1740 723 1765 726
rect 1836 723 1861 726
rect 1906 723 1916 726
rect 1946 723 1972 726
rect 2066 723 2076 726
rect 2164 723 2189 726
rect 2226 723 2236 726
rect 2452 723 2525 726
rect 2538 725 2557 726
rect 2540 723 2557 725
rect 2588 723 2597 726
rect 2602 723 2676 726
rect 2770 723 2788 726
rect 2890 723 2900 726
rect 2980 723 3021 726
rect 3028 723 3069 726
rect 3076 723 3101 726
rect 3218 723 3252 726
rect 3284 723 3301 726
rect 3356 723 3381 726
rect 3444 723 3469 726
rect 3474 723 3492 726
rect 3514 723 3540 726
rect 3570 723 3604 726
rect 3642 723 3668 726
rect 3762 723 3804 726
rect 4018 723 4028 726
rect 4074 723 4100 726
rect 4130 723 4236 726
rect 4266 723 4284 726
rect 4322 723 4325 733
rect 4770 726 4773 733
rect 4338 723 4348 726
rect 4426 723 4452 726
rect 4490 723 4516 726
rect 4562 723 4588 726
rect 4690 723 4724 726
rect 4754 723 4764 726
rect 4770 723 4789 726
rect 2594 716 2597 723
rect 2594 713 2645 716
rect 3082 713 3116 716
rect 3140 713 3165 716
rect 3508 713 3525 716
rect 3620 713 3645 716
rect 14 667 4853 673
rect 2380 623 2413 626
rect 3060 623 3077 626
rect 3114 623 3124 626
rect 284 613 309 616
rect 340 613 365 616
rect 370 613 380 616
rect 514 613 540 616
rect 580 613 597 616
rect 690 613 700 616
rect 706 613 716 616
rect 746 613 764 616
rect 810 613 828 616
rect 866 613 876 616
rect 914 613 940 616
rect 1004 613 1021 616
rect 1044 613 1069 616
rect 1084 613 1093 616
rect 1098 613 1124 616
rect 1146 613 1196 616
rect 1306 613 1340 616
rect 1346 613 1380 616
rect 1426 613 1436 616
rect 1490 613 1500 616
rect 1554 613 1564 616
rect 1610 613 1620 616
rect 1682 613 1724 616
rect 1810 613 1828 616
rect 1930 613 1948 616
rect 2010 613 2020 616
rect 2058 613 2068 616
rect 2098 613 2124 616
rect 2162 613 2172 616
rect 2354 613 2372 616
rect 2450 613 2460 616
rect 2522 613 2549 616
rect 2580 613 2605 616
rect 2610 613 2620 616
rect 2754 613 2764 616
rect 1554 606 1557 613
rect 1682 606 1685 613
rect 116 603 173 606
rect 196 603 221 606
rect 354 603 372 606
rect 514 603 532 606
rect 586 603 620 606
rect 642 603 676 606
rect 738 603 756 606
rect 788 603 821 606
rect 858 603 868 606
rect 978 603 996 606
rect 1036 603 1061 606
rect 1076 603 1117 606
rect 1148 603 1189 606
rect 1194 603 1204 606
rect 1220 603 1276 606
rect 1308 603 1325 606
rect 1524 603 1557 606
rect 1676 603 1685 606
rect 1780 603 1820 606
rect 2306 603 2332 606
rect 2402 603 2420 606
rect 2500 603 2541 606
rect 2546 605 2549 613
rect 2602 606 2605 613
rect 2874 606 2877 616
rect 2900 613 2973 616
rect 2980 613 2997 616
rect 3066 613 3084 616
rect 3308 613 3333 616
rect 3428 613 3453 616
rect 3460 613 3477 616
rect 3484 613 3509 616
rect 3540 613 3565 616
rect 3586 613 3628 616
rect 3666 613 3724 616
rect 3868 613 3932 616
rect 4260 613 4285 616
rect 4316 613 4325 616
rect 4330 613 4348 616
rect 4386 613 4428 616
rect 4490 613 4500 616
rect 4538 613 4572 616
rect 2602 603 2628 606
rect 2858 605 2877 606
rect 2970 605 2973 613
rect 2858 603 2876 605
rect 3020 603 3029 606
rect 3106 603 3124 606
rect 3148 603 3173 606
rect 3450 605 3453 613
rect 3466 603 3476 606
rect 3490 603 3508 606
rect 3554 603 3564 606
rect 3594 603 3620 606
rect 3644 603 3717 606
rect 3796 603 3821 606
rect 3826 603 3844 606
rect 3956 603 4004 606
rect 4116 603 4157 606
rect 4372 603 4389 606
rect 4458 603 4492 606
rect 4596 603 4628 606
rect 978 593 988 596
rect 1002 593 1028 596
rect 1042 593 1068 596
rect 3162 593 3172 596
rect 38 567 4829 573
rect 938 543 972 546
rect 986 543 996 546
rect 1010 543 1036 546
rect 3050 543 3092 546
rect 3242 543 3252 546
rect 180 533 205 536
rect 364 533 389 536
rect 466 533 500 536
rect 514 533 564 536
rect 628 533 637 536
rect 788 533 836 536
rect 858 533 900 536
rect 932 533 941 536
rect 946 533 980 536
rect 1004 533 1029 536
rect 1044 533 1053 536
rect 1194 533 1212 536
rect 1228 533 1268 536
rect 1300 533 1309 536
rect 1322 533 1340 536
rect 1362 533 1396 536
rect 1434 533 1508 536
rect 1530 533 1572 536
rect 1676 533 1685 536
rect 1756 533 1780 536
rect 1802 533 1812 536
rect 1858 533 1892 536
rect 1914 533 1948 536
rect 1970 533 1996 536
rect 2426 533 2444 536
rect 3036 533 3077 536
rect 3186 533 3236 536
rect 3250 533 3260 536
rect 186 523 204 526
rect 236 523 245 526
rect 346 523 356 526
rect 378 523 388 526
rect 426 523 436 526
rect 468 523 477 526
rect 498 523 508 526
rect 530 523 572 526
rect 676 523 685 526
rect 738 523 764 526
rect 802 523 828 526
rect 866 523 908 526
rect 988 523 997 526
rect 1012 523 1037 526
rect 1092 523 1101 526
rect 1178 523 1204 526
rect 1292 523 1301 526
rect 1364 523 1397 526
rect 1404 523 1429 526
rect 1442 523 1500 526
rect 1532 523 1541 526
rect 1580 523 1613 526
rect 1714 523 1732 526
rect 1890 523 1900 526
rect 1922 523 1940 526
rect 2004 523 2013 526
rect 2090 523 2100 526
rect 2188 523 2197 526
rect 2300 523 2309 526
rect 2356 523 2365 526
rect 2370 523 2388 526
rect 2434 523 2468 526
rect 2514 523 2532 526
rect 2580 523 2605 526
rect 2916 523 2940 526
rect 2964 523 2973 526
rect 3012 524 3028 527
rect 3442 526 3445 534
rect 3458 533 3468 536
rect 3498 533 3516 536
rect 3586 533 3604 536
rect 3628 534 3660 536
rect 3628 533 3661 534
rect 3692 533 3717 536
rect 3114 523 3156 526
rect 3268 523 3277 526
rect 3380 523 3445 526
rect 3452 523 3461 526
rect 3476 523 3509 526
rect 3538 523 3564 526
rect 3602 523 3612 526
rect 3658 523 3661 533
rect 3762 523 3788 526
rect 3884 523 3932 526
rect 3938 523 3941 534
rect 3946 533 3980 536
rect 4028 533 4037 536
rect 4042 533 4076 536
rect 4162 526 4165 534
rect 4308 533 4317 536
rect 4338 533 4348 536
rect 4380 533 4420 536
rect 4458 533 4492 536
rect 4524 533 4564 536
rect 4668 533 4677 536
rect 4690 533 4700 536
rect 4772 533 4781 536
rect 4004 523 4020 526
rect 4100 523 4156 526
rect 4162 523 4180 526
rect 4210 523 4236 526
rect 4300 523 4356 526
rect 4516 523 4565 526
rect 4578 523 4604 526
rect 4634 523 4660 526
rect 4682 523 4708 526
rect 4738 523 4764 526
rect 3010 513 3020 516
rect 3460 513 3469 516
rect 3580 513 3597 516
rect 3004 503 3021 506
rect 14 467 4853 473
rect 2612 433 2629 436
rect 3052 433 3069 436
rect 3092 433 3117 436
rect 2628 423 2637 426
rect 3026 423 3044 426
rect 3068 423 3077 426
rect 3098 423 3108 426
rect 3570 423 3580 426
rect 3026 416 3029 423
rect 108 413 133 416
rect 164 413 197 416
rect 202 403 205 414
rect 290 413 316 416
rect 348 413 388 416
rect 420 413 437 416
rect 484 413 501 416
rect 562 413 580 416
rect 610 406 613 416
rect 618 413 644 416
rect 700 413 709 416
rect 852 413 861 416
rect 882 413 932 416
rect 1018 413 1044 416
rect 1100 413 1125 416
rect 1220 413 1229 416
rect 1234 413 1308 416
rect 1458 413 1500 416
rect 1642 413 1652 416
rect 1666 413 1684 416
rect 1858 413 1884 416
rect 1916 413 1925 416
rect 1970 413 1980 416
rect 2060 413 2069 416
rect 2106 413 2132 416
rect 2170 413 2180 416
rect 2226 413 2236 416
rect 2282 413 2292 416
rect 2410 406 2413 416
rect 2460 413 2469 416
rect 2516 413 2525 416
rect 2540 413 2557 416
rect 2684 413 2709 416
rect 2740 413 2749 416
rect 2892 413 2909 416
rect 2970 413 2980 416
rect 3020 413 3029 416
rect 3228 413 3237 416
rect 3284 413 3317 416
rect 3420 413 3437 416
rect 3484 413 3509 416
rect 3524 413 3541 416
rect 3588 413 3605 416
rect 3698 413 3724 416
rect 3730 413 3773 416
rect 3804 413 3829 416
rect 3868 413 3877 416
rect 3924 413 3941 416
rect 3980 413 3997 416
rect 4092 413 4124 416
rect 4186 413 4204 416
rect 4260 413 4285 416
rect 4372 413 4397 416
rect 4428 413 4437 416
rect 4500 413 4509 416
rect 3770 406 3773 413
rect 340 403 381 406
rect 418 403 436 406
rect 546 403 572 406
rect 610 403 652 406
rect 674 403 692 406
rect 962 403 972 406
rect 1092 403 1117 406
rect 1290 403 1316 406
rect 1508 403 1517 406
rect 1660 403 1685 406
rect 1914 403 1948 406
rect 1962 403 1988 406
rect 2010 403 2052 406
rect 2396 403 2413 406
rect 2522 403 2532 406
rect 2546 403 2564 406
rect 2994 403 3012 406
rect 3114 403 3148 406
rect 3426 403 3452 406
rect 3466 403 3476 406
rect 3692 403 3717 406
rect 3732 403 3741 406
rect 3746 403 3756 406
rect 3770 403 3780 406
rect 4100 403 4109 406
rect 4132 403 4141 406
rect 4434 405 4437 413
rect 3122 393 3140 396
rect 3122 383 3125 393
rect 38 367 4829 373
rect 1074 343 1092 346
rect 1114 343 1124 346
rect 1138 343 1148 346
rect 1162 343 1204 346
rect 3586 343 3597 346
rect 3586 336 3589 343
rect 188 333 221 336
rect 372 333 389 336
rect 594 333 628 336
rect 938 333 956 336
rect 1090 333 1100 336
rect 1156 333 1173 336
rect 1202 333 1212 336
rect 1284 333 1333 336
rect 1660 333 1669 336
rect 1708 333 1749 336
rect 1772 333 1797 336
rect 2002 333 2036 336
rect 2194 333 2220 336
rect 2570 333 2604 336
rect 2764 333 2788 336
rect 3042 333 3052 336
rect 3084 333 3101 336
rect 116 323 141 326
rect 276 323 301 326
rect 338 323 364 326
rect 370 323 388 326
rect 594 323 597 333
rect 1794 326 1797 333
rect 3402 326 3405 335
rect 3418 333 3428 336
rect 3442 333 3452 336
rect 3500 333 3509 336
rect 3516 333 3533 336
rect 3580 333 3589 336
rect 3594 333 3604 336
rect 3628 333 3637 336
rect 3866 326 3869 335
rect 3930 333 3956 336
rect 3978 333 3996 336
rect 4322 333 4348 336
rect 4380 333 4389 336
rect 4394 333 4412 336
rect 4434 333 4452 336
rect 4540 333 4549 336
rect 4554 333 4604 336
rect 3978 326 3981 333
rect 4386 326 4389 333
rect 4434 326 4437 333
rect 636 323 685 326
rect 858 323 868 326
rect 940 323 949 326
rect 964 323 973 326
rect 1010 323 1036 326
rect 1108 323 1125 326
rect 1140 323 1149 326
rect 1164 323 1205 326
rect 1234 323 1260 326
rect 1722 323 1748 326
rect 1794 323 1804 326
rect 1954 323 1964 326
rect 2018 323 2028 326
rect 2194 323 2228 326
rect 2242 323 2260 326
rect 2290 323 2316 326
rect 2410 323 2420 326
rect 2466 323 2476 326
rect 2586 323 2612 326
rect 2732 323 2756 326
rect 2844 323 2861 326
rect 2914 323 2948 326
rect 2986 323 3004 326
rect 3066 323 3076 326
rect 3082 323 3108 326
rect 3140 323 3157 326
rect 3252 323 3269 326
rect 3364 323 3405 326
rect 3418 323 3436 326
rect 3460 323 3485 326
rect 3492 323 3501 326
rect 3586 323 3612 326
rect 3788 323 3797 326
rect 3844 323 3869 326
rect 3964 323 3981 326
rect 4020 323 4036 326
rect 4146 323 4156 326
rect 4242 323 4268 326
rect 4316 323 4356 326
rect 4386 323 4437 326
rect 4476 323 4532 326
rect 4628 323 4645 326
rect 3418 315 3421 323
rect 3468 313 3484 316
rect 3580 313 3589 316
rect 3628 313 3645 316
rect 14 267 4853 273
rect 1762 223 1781 226
rect 2700 223 2708 226
rect 3468 223 3485 226
rect 1762 216 1765 223
rect 114 213 140 216
rect 226 213 236 216
rect 348 213 357 216
rect 420 213 437 216
rect 468 213 485 216
rect 570 213 580 216
rect 618 213 644 216
rect 682 213 692 216
rect 698 213 724 216
rect 754 213 804 216
rect 834 213 844 216
rect 914 213 940 216
rect 986 213 1012 216
rect 1076 213 1085 216
rect 1124 213 1133 216
rect 1138 213 1148 216
rect 1228 213 1237 216
rect 1338 213 1348 216
rect 1458 213 1484 216
rect 1564 213 1573 216
rect 1586 213 1604 216
rect 1668 213 1685 216
rect 1748 213 1765 216
rect 1770 213 1788 216
rect 1986 213 1996 216
rect 2010 213 2036 216
rect 2114 213 2132 216
rect 2170 213 2188 216
rect 2234 213 2244 216
rect 2410 213 2420 216
rect 2572 213 2581 216
rect 2586 213 2621 216
rect 2636 213 2653 216
rect 2660 213 2677 216
rect 2722 213 2740 216
rect 2746 213 2756 216
rect 2788 213 2797 216
rect 2802 213 2812 216
rect 2818 213 2852 216
rect 2890 213 2908 216
rect 2938 213 2972 216
rect 3052 213 3069 216
rect 3188 213 3197 216
rect 3292 213 3309 216
rect 3460 213 3477 216
rect 3530 213 3556 216
rect 3588 213 3597 216
rect 3612 213 3636 216
rect 3700 213 3724 216
rect 3772 213 3812 216
rect 4108 213 4141 216
rect 4228 213 4253 216
rect 4284 213 4293 216
rect 148 203 173 206
rect 196 203 213 206
rect 228 203 237 206
rect 340 203 373 206
rect 402 203 412 206
rect 522 203 532 206
rect 570 203 588 206
rect 604 203 645 206
rect 674 203 684 206
rect 706 203 716 206
rect 754 203 796 206
rect 868 203 877 206
rect 898 203 948 206
rect 970 203 1004 206
rect 1068 203 1077 206
rect 1116 203 1149 206
rect 1178 203 1188 206
rect 1276 203 1325 206
rect 1340 203 1349 206
rect 1378 203 1412 206
rect 1434 203 1444 206
rect 1466 203 1492 206
rect 1514 203 1556 206
rect 1578 203 1596 206
rect 1634 203 1644 206
rect 1682 203 1724 206
rect 1740 203 1749 206
rect 1754 203 1796 206
rect 1826 203 1852 206
rect 1866 203 1932 206
rect 1954 203 1988 206
rect 2002 203 2044 206
rect 2074 203 2100 206
rect 2578 203 2604 206
rect 2634 203 2652 206
rect 2674 205 2677 213
rect 2700 203 2709 206
rect 2746 205 2749 213
rect 3066 206 3069 213
rect 4394 206 4397 216
rect 4756 213 4765 216
rect 2820 203 2837 206
rect 2892 203 2901 206
rect 3026 203 3036 206
rect 3066 203 3076 206
rect 3410 203 3452 206
rect 3466 203 3484 206
rect 3660 203 3676 206
rect 3738 203 3748 206
rect 3826 203 3836 206
rect 3884 203 3917 206
rect 3930 203 3948 206
rect 3996 203 4005 206
rect 4116 203 4133 206
rect 4340 203 4357 206
rect 4362 203 4404 206
rect 4588 203 4596 206
rect 1018 193 1060 196
rect 38 167 4829 173
rect 850 133 884 136
rect 900 133 925 136
rect 2586 133 2596 136
rect 2810 126 2813 135
rect 2826 133 2844 136
rect 2850 133 2868 136
rect 2956 133 2973 136
rect 3194 126 3197 135
rect 4594 133 4628 136
rect 108 123 117 126
rect 204 123 221 126
rect 668 123 685 126
rect 746 123 756 126
rect 1324 123 1333 126
rect 1380 123 1389 126
rect 1450 123 1460 126
rect 1506 123 1524 126
rect 1570 123 1580 126
rect 1730 123 1740 126
rect 1882 123 1892 126
rect 2042 123 2052 126
rect 2492 123 2517 126
rect 2548 123 2581 126
rect 2610 123 2620 126
rect 2650 123 2676 126
rect 2748 123 2773 126
rect 2804 123 2813 126
rect 2820 123 2837 126
rect 2852 123 2861 126
rect 2938 123 2948 126
rect 2954 123 2972 126
rect 3004 123 3052 126
rect 3082 123 3108 126
rect 3146 123 3188 126
rect 3194 123 3204 126
rect 3298 123 3308 126
rect 3548 123 3573 126
rect 3652 123 3677 126
rect 3708 123 3717 126
rect 3756 123 3765 126
rect 3812 123 3821 126
rect 4084 123 4093 126
rect 4300 123 4309 126
rect 4412 123 4421 126
rect 4516 123 4541 126
rect 4580 123 4605 126
rect 14 67 4853 73
rect 38 37 4829 57
rect 14 13 4853 33
<< metal2 >>
rect 14 13 34 4727
rect 38 37 58 4703
rect 90 4593 93 4606
rect 114 4546 117 4616
rect 98 4543 117 4546
rect 90 4513 93 4536
rect 98 4523 101 4543
rect 106 4533 117 4536
rect 138 4533 141 4546
rect 114 4413 117 4526
rect 130 4503 133 4526
rect 146 4513 149 4526
rect 170 4446 173 4616
rect 242 4613 245 4626
rect 282 4613 285 4626
rect 234 4573 237 4606
rect 258 4593 261 4606
rect 170 4443 181 4446
rect 90 4383 93 4406
rect 178 4403 181 4443
rect 194 4436 197 4546
rect 202 4483 205 4526
rect 210 4523 213 4536
rect 218 4523 221 4536
rect 226 4496 229 4536
rect 234 4533 237 4546
rect 226 4493 237 4496
rect 186 4433 197 4436
rect 186 4406 189 4433
rect 194 4413 197 4426
rect 186 4403 197 4406
rect 194 4386 197 4403
rect 186 4383 197 4386
rect 82 3686 85 4216
rect 114 4123 117 4216
rect 154 4123 157 4136
rect 162 4133 165 4326
rect 186 4266 189 4383
rect 186 4263 197 4266
rect 186 4226 189 4246
rect 178 4223 189 4226
rect 178 4146 181 4223
rect 178 4143 189 4146
rect 186 4126 189 4143
rect 194 4133 197 4263
rect 162 4113 165 4126
rect 170 4123 181 4126
rect 186 4123 197 4126
rect 130 4013 133 4026
rect 162 4013 165 4036
rect 170 4013 173 4026
rect 130 3913 133 3926
rect 162 3903 165 3926
rect 170 3913 173 3926
rect 106 3723 109 3816
rect 138 3793 141 3806
rect 170 3803 173 3826
rect 82 3683 93 3686
rect 90 3603 93 3683
rect 154 3656 157 3746
rect 170 3723 173 3786
rect 186 3743 189 4123
rect 194 3883 197 4016
rect 202 4013 205 4126
rect 210 4123 213 4416
rect 218 4393 221 4406
rect 218 4333 221 4356
rect 226 4313 229 4416
rect 234 4403 237 4493
rect 242 4456 245 4526
rect 250 4493 253 4526
rect 258 4506 261 4526
rect 266 4523 269 4576
rect 258 4503 265 4506
rect 242 4453 249 4456
rect 234 4206 237 4386
rect 246 4356 249 4453
rect 262 4446 265 4503
rect 258 4443 265 4446
rect 246 4353 253 4356
rect 242 4306 245 4336
rect 250 4323 253 4353
rect 258 4333 261 4443
rect 274 4383 277 4596
rect 306 4533 309 4546
rect 338 4543 341 4616
rect 386 4613 389 4626
rect 378 4593 381 4606
rect 402 4603 405 4616
rect 426 4613 429 4626
rect 346 4543 365 4546
rect 346 4533 349 4543
rect 282 4503 285 4526
rect 306 4413 309 4526
rect 322 4503 325 4526
rect 354 4413 357 4536
rect 362 4523 365 4543
rect 370 4533 373 4556
rect 378 4523 381 4566
rect 386 4473 389 4526
rect 402 4523 405 4596
rect 418 4503 421 4526
rect 434 4456 437 4566
rect 482 4533 485 4616
rect 506 4576 509 4606
rect 502 4573 509 4576
rect 490 4513 493 4536
rect 502 4456 505 4573
rect 530 4546 533 4616
rect 514 4543 533 4546
rect 514 4523 517 4543
rect 434 4453 445 4456
rect 502 4453 509 4456
rect 402 4413 413 4416
rect 346 4343 365 4346
rect 242 4303 253 4306
rect 250 4236 253 4303
rect 282 4256 285 4316
rect 282 4253 289 4256
rect 242 4233 253 4236
rect 242 4213 245 4233
rect 234 4203 245 4206
rect 202 3996 205 4006
rect 210 4003 213 4036
rect 218 3996 221 4016
rect 202 3993 221 3996
rect 202 3943 221 3946
rect 202 3933 205 3943
rect 210 3903 213 3936
rect 218 3923 221 3943
rect 202 3763 205 3866
rect 154 3653 161 3656
rect 138 3613 141 3626
rect 158 3576 161 3653
rect 170 3593 173 3616
rect 178 3613 181 3626
rect 154 3573 161 3576
rect 82 3533 85 3556
rect 130 3513 133 3526
rect 154 3443 157 3573
rect 186 3553 189 3736
rect 210 3723 213 3816
rect 218 3813 221 3846
rect 218 3786 221 3806
rect 226 3803 229 4146
rect 242 4133 245 4203
rect 286 4176 289 4253
rect 298 4206 301 4336
rect 306 4213 309 4326
rect 322 4323 325 4336
rect 346 4333 349 4343
rect 354 4323 357 4336
rect 362 4323 365 4343
rect 370 4333 373 4346
rect 378 4243 381 4376
rect 298 4203 309 4206
rect 282 4173 289 4176
rect 234 4013 237 4026
rect 242 3863 245 4126
rect 282 4106 285 4173
rect 306 4166 309 4203
rect 330 4193 333 4206
rect 362 4203 365 4216
rect 386 4166 389 4196
rect 306 4163 313 4166
rect 290 4113 293 4126
rect 282 4103 293 4106
rect 266 4003 269 4036
rect 282 4003 285 4086
rect 258 3933 261 3966
rect 290 3956 293 4103
rect 310 4086 313 4163
rect 378 4163 389 4166
rect 306 4083 313 4086
rect 290 3953 301 3956
rect 234 3793 237 3816
rect 218 3783 225 3786
rect 242 3783 245 3806
rect 250 3786 253 3886
rect 258 3813 261 3846
rect 266 3803 269 3946
rect 274 3943 293 3946
rect 274 3923 277 3943
rect 282 3903 285 3936
rect 290 3933 293 3943
rect 274 3813 277 3826
rect 290 3813 293 3926
rect 298 3906 301 3953
rect 306 3923 309 4083
rect 322 4003 325 4126
rect 330 4113 333 4126
rect 330 3906 333 4026
rect 346 4013 349 4136
rect 378 4116 381 4163
rect 394 4123 397 4216
rect 410 4213 413 4386
rect 442 4376 445 4453
rect 458 4413 461 4426
rect 434 4373 445 4376
rect 434 4346 437 4373
rect 434 4343 445 4346
rect 442 4296 445 4343
rect 458 4313 461 4326
rect 434 4293 445 4296
rect 378 4113 389 4116
rect 362 4013 365 4066
rect 354 3943 357 4006
rect 362 3913 365 3926
rect 298 3903 309 3906
rect 330 3903 341 3906
rect 306 3836 309 3903
rect 298 3833 309 3836
rect 274 3786 277 3806
rect 250 3783 261 3786
rect 222 3716 225 3783
rect 218 3713 225 3716
rect 162 3523 165 3546
rect 170 3513 173 3526
rect 194 3523 197 3676
rect 210 3596 213 3606
rect 218 3603 221 3713
rect 234 3686 237 3766
rect 234 3683 245 3686
rect 226 3596 229 3616
rect 210 3593 229 3596
rect 234 3593 237 3606
rect 202 3543 221 3546
rect 202 3533 205 3543
rect 210 3523 213 3536
rect 218 3523 221 3543
rect 226 3533 229 3546
rect 234 3503 237 3526
rect 210 3426 213 3446
rect 242 3436 245 3683
rect 250 3536 253 3626
rect 258 3603 261 3783
rect 270 3783 277 3786
rect 270 3716 273 3783
rect 282 3723 285 3806
rect 298 3803 301 3833
rect 290 3733 293 3786
rect 270 3713 277 3716
rect 274 3623 277 3713
rect 306 3636 309 3816
rect 322 3803 325 3896
rect 338 3836 341 3903
rect 330 3833 341 3836
rect 314 3733 317 3756
rect 306 3633 313 3636
rect 274 3603 277 3616
rect 298 3613 301 3626
rect 250 3533 261 3536
rect 238 3433 245 3436
rect 186 3413 189 3426
rect 206 3423 213 3426
rect 138 3336 141 3406
rect 206 3356 209 3423
rect 206 3353 213 3356
rect 90 3286 93 3336
rect 130 3333 141 3336
rect 90 3283 101 3286
rect 98 3056 101 3283
rect 130 3276 133 3333
rect 138 3313 141 3326
rect 170 3323 173 3346
rect 178 3313 181 3326
rect 202 3313 205 3336
rect 130 3273 141 3276
rect 114 3213 117 3226
rect 114 3193 117 3206
rect 82 3053 101 3056
rect 138 3056 141 3273
rect 162 3213 165 3226
rect 210 3216 213 3353
rect 218 3333 221 3416
rect 226 3413 229 3426
rect 206 3213 213 3216
rect 206 3156 209 3213
rect 226 3206 229 3376
rect 238 3346 241 3433
rect 258 3426 261 3533
rect 250 3423 261 3426
rect 250 3346 253 3423
rect 258 3353 261 3416
rect 266 3403 269 3426
rect 274 3413 277 3556
rect 282 3533 293 3536
rect 298 3533 301 3596
rect 310 3576 313 3633
rect 306 3573 313 3576
rect 306 3553 309 3573
rect 322 3553 325 3776
rect 330 3756 333 3833
rect 338 3803 349 3806
rect 354 3773 357 3816
rect 370 3803 373 3926
rect 386 3886 389 4113
rect 434 4036 437 4293
rect 458 4123 461 4206
rect 482 4156 485 4436
rect 506 4433 509 4453
rect 498 4413 501 4426
rect 490 4303 493 4326
rect 498 4313 501 4326
rect 514 4216 517 4506
rect 522 4473 525 4526
rect 530 4286 533 4536
rect 562 4533 565 4546
rect 570 4533 573 4556
rect 586 4543 589 4616
rect 658 4613 661 4626
rect 610 4593 613 4606
rect 538 4513 541 4526
rect 538 4413 541 4496
rect 562 4426 565 4526
rect 578 4476 581 4526
rect 586 4523 589 4536
rect 602 4533 605 4546
rect 594 4493 597 4526
rect 578 4473 589 4476
rect 546 4396 549 4406
rect 554 4403 557 4426
rect 562 4423 581 4426
rect 562 4396 565 4416
rect 570 4403 573 4416
rect 578 4413 581 4423
rect 546 4393 565 4396
rect 546 4343 565 4346
rect 546 4333 549 4343
rect 554 4303 557 4336
rect 562 4323 565 4343
rect 530 4283 541 4286
rect 482 4153 493 4156
rect 466 4143 485 4146
rect 466 4133 469 4143
rect 466 4046 469 4126
rect 474 4123 477 4136
rect 482 4123 485 4143
rect 426 4033 437 4036
rect 426 3946 429 4033
rect 434 4013 437 4026
rect 458 3956 461 4046
rect 466 4043 485 4046
rect 490 4043 493 4153
rect 498 4133 501 4216
rect 510 4213 517 4216
rect 510 4156 513 4213
rect 510 4153 517 4156
rect 498 4103 501 4126
rect 506 4123 509 4136
rect 514 4113 517 4153
rect 522 4093 525 4206
rect 530 4183 533 4216
rect 538 4203 541 4283
rect 570 4243 573 4336
rect 546 4196 549 4216
rect 554 4203 557 4216
rect 570 4213 573 4236
rect 586 4216 589 4473
rect 578 4213 589 4216
rect 562 4196 565 4206
rect 546 4193 565 4196
rect 546 4143 565 4146
rect 530 4096 533 4126
rect 546 4123 549 4143
rect 554 4103 557 4136
rect 562 4133 565 4143
rect 562 4113 565 4126
rect 530 4093 549 4096
rect 466 4013 469 4036
rect 474 4013 477 4026
rect 418 3943 429 3946
rect 450 3953 461 3956
rect 402 3913 405 3926
rect 386 3883 405 3886
rect 330 3753 341 3756
rect 330 3733 333 3746
rect 290 3493 293 3533
rect 282 3413 285 3426
rect 274 3383 277 3406
rect 282 3403 293 3406
rect 282 3373 285 3403
rect 238 3343 245 3346
rect 250 3343 261 3346
rect 218 3203 229 3206
rect 206 3153 213 3156
rect 146 3113 149 3126
rect 138 3053 149 3056
rect 82 2743 85 3053
rect 146 3036 149 3053
rect 146 3033 153 3036
rect 98 2913 101 2936
rect 106 2923 109 3016
rect 122 2746 125 3006
rect 150 2976 153 3033
rect 146 2973 153 2976
rect 146 2856 149 2973
rect 162 2933 165 3016
rect 170 3013 173 3116
rect 178 2876 181 3036
rect 186 2996 189 3006
rect 194 3003 197 3126
rect 210 3106 213 3153
rect 218 3133 221 3203
rect 226 3123 229 3196
rect 210 3103 221 3106
rect 202 2996 205 3016
rect 186 2993 205 2996
rect 202 2913 205 2926
rect 210 2903 213 3006
rect 218 3003 221 3103
rect 234 3023 237 3216
rect 242 3163 245 3343
rect 250 3323 253 3336
rect 258 3236 261 3343
rect 266 3333 269 3346
rect 290 3316 293 3396
rect 298 3373 301 3526
rect 314 3333 317 3536
rect 330 3533 333 3576
rect 338 3563 341 3753
rect 362 3646 365 3746
rect 402 3743 405 3883
rect 418 3866 421 3943
rect 450 3933 453 3953
rect 418 3863 429 3866
rect 426 3766 429 3863
rect 434 3813 437 3896
rect 466 3893 469 3926
rect 426 3763 433 3766
rect 410 3713 413 3726
rect 430 3656 433 3763
rect 442 3703 445 3726
rect 458 3713 461 3726
rect 430 3653 437 3656
rect 346 3643 365 3646
rect 346 3573 349 3643
rect 354 3613 357 3636
rect 362 3613 365 3626
rect 370 3603 373 3616
rect 402 3596 405 3606
rect 410 3603 413 3636
rect 418 3596 421 3616
rect 426 3603 429 3646
rect 402 3593 421 3596
rect 378 3513 381 3526
rect 410 3523 413 3546
rect 418 3513 421 3526
rect 322 3393 325 3406
rect 338 3376 341 3406
rect 322 3373 341 3376
rect 298 3323 309 3326
rect 290 3313 301 3316
rect 250 3233 261 3236
rect 250 3186 253 3233
rect 250 3183 261 3186
rect 258 3136 261 3183
rect 266 3143 269 3256
rect 258 3133 269 3136
rect 242 3086 245 3126
rect 242 3083 253 3086
rect 250 3036 253 3083
rect 242 3033 253 3036
rect 218 2933 221 2946
rect 234 2883 237 2926
rect 242 2916 245 3033
rect 250 3003 253 3016
rect 266 2966 269 3133
rect 274 2983 277 3006
rect 258 2963 269 2966
rect 258 2923 261 2963
rect 266 2933 269 2956
rect 282 2946 285 3166
rect 298 3156 301 3313
rect 306 3293 309 3323
rect 314 3313 317 3326
rect 322 3253 325 3373
rect 330 3303 333 3336
rect 314 3213 317 3226
rect 294 3153 301 3156
rect 294 3106 297 3153
rect 338 3146 341 3366
rect 346 3333 349 3346
rect 354 3313 357 3336
rect 362 3323 365 3416
rect 378 3333 381 3406
rect 418 3403 421 3416
rect 394 3333 397 3346
rect 402 3333 405 3396
rect 434 3366 437 3653
rect 482 3646 485 4043
rect 498 3906 501 4016
rect 514 3996 517 4006
rect 522 4003 525 4036
rect 530 3996 533 4016
rect 546 4013 549 4093
rect 514 3993 533 3996
rect 530 3943 549 3946
rect 530 3933 533 3943
rect 498 3903 509 3906
rect 506 3766 509 3903
rect 530 3896 533 3916
rect 522 3893 533 3896
rect 522 3806 525 3893
rect 538 3813 541 3936
rect 546 3923 549 3943
rect 554 3826 557 4096
rect 562 3893 565 4016
rect 554 3823 565 3826
rect 522 3803 533 3806
rect 498 3763 509 3766
rect 482 3643 489 3646
rect 442 3523 445 3626
rect 458 3593 461 3616
rect 486 3576 489 3643
rect 482 3573 489 3576
rect 434 3363 445 3366
rect 346 3213 349 3236
rect 354 3213 357 3226
rect 370 3213 373 3326
rect 386 3313 389 3326
rect 294 3103 301 3106
rect 290 3013 293 3026
rect 274 2943 285 2946
rect 274 2923 277 2943
rect 242 2913 269 2916
rect 178 2873 213 2876
rect 146 2853 173 2856
rect 154 2813 157 2826
rect 154 2793 157 2806
rect 98 2656 101 2746
rect 122 2743 133 2746
rect 130 2696 133 2743
rect 146 2713 149 2726
rect 82 2653 101 2656
rect 122 2693 133 2696
rect 170 2693 173 2853
rect 194 2813 197 2826
rect 210 2806 213 2873
rect 202 2803 213 2806
rect 178 2703 181 2726
rect 186 2713 189 2726
rect 202 2723 205 2803
rect 218 2743 237 2746
rect 218 2733 221 2743
rect 218 2696 221 2726
rect 226 2703 229 2736
rect 234 2723 237 2743
rect 242 2716 245 2906
rect 266 2803 269 2913
rect 282 2826 285 2936
rect 298 2906 301 3103
rect 314 2933 317 3146
rect 338 3143 349 3146
rect 346 3096 349 3143
rect 338 3093 349 3096
rect 338 2946 341 3093
rect 362 3013 365 3126
rect 394 3056 397 3216
rect 402 3196 405 3206
rect 410 3203 413 3236
rect 418 3196 421 3216
rect 426 3203 429 3346
rect 434 3313 437 3326
rect 442 3213 445 3363
rect 450 3306 453 3556
rect 482 3553 485 3573
rect 466 3543 485 3546
rect 466 3533 469 3543
rect 474 3523 477 3536
rect 482 3523 485 3543
rect 490 3533 493 3546
rect 498 3503 501 3763
rect 506 3743 525 3746
rect 506 3733 509 3743
rect 514 3703 517 3736
rect 522 3723 525 3743
rect 530 3646 533 3803
rect 546 3723 549 3816
rect 562 3756 565 3823
rect 554 3753 565 3756
rect 554 3733 557 3753
rect 522 3643 533 3646
rect 506 3613 509 3626
rect 506 3533 509 3596
rect 522 3513 525 3643
rect 530 3533 533 3636
rect 538 3613 541 3646
rect 546 3613 549 3626
rect 554 3586 557 3656
rect 578 3593 581 4213
rect 586 3923 589 3936
rect 594 3906 597 4246
rect 602 4233 605 4406
rect 610 4403 613 4536
rect 618 4513 621 4526
rect 642 4436 645 4496
rect 642 4433 653 4436
rect 626 4413 629 4426
rect 642 4413 645 4433
rect 634 4403 645 4406
rect 650 4403 653 4416
rect 658 4413 661 4426
rect 666 4356 669 4436
rect 674 4403 677 4446
rect 690 4413 693 4616
rect 698 4613 701 4626
rect 698 4523 701 4606
rect 706 4503 709 4536
rect 714 4523 717 4616
rect 810 4613 813 4626
rect 730 4533 733 4546
rect 706 4413 709 4436
rect 698 4383 701 4406
rect 714 4403 717 4416
rect 738 4403 741 4426
rect 754 4413 757 4526
rect 762 4513 765 4606
rect 842 4583 845 4616
rect 850 4613 853 4626
rect 850 4556 853 4606
rect 842 4553 853 4556
rect 858 4603 869 4606
rect 762 4413 765 4456
rect 666 4353 677 4356
rect 610 4333 613 4346
rect 634 4343 653 4346
rect 618 4293 621 4326
rect 634 4323 637 4343
rect 642 4303 645 4336
rect 650 4333 653 4343
rect 610 4213 613 4226
rect 618 4036 621 4116
rect 626 4043 629 4266
rect 650 4233 653 4326
rect 674 4266 677 4353
rect 698 4313 701 4326
rect 666 4263 677 4266
rect 714 4263 717 4336
rect 738 4313 741 4326
rect 666 4246 669 4263
rect 658 4243 669 4246
rect 650 4213 653 4226
rect 658 4166 661 4243
rect 698 4213 709 4216
rect 738 4203 741 4226
rect 746 4213 749 4336
rect 754 4223 757 4406
rect 770 4403 773 4506
rect 778 4413 781 4426
rect 794 4333 797 4416
rect 810 4403 813 4546
rect 818 4503 821 4536
rect 826 4473 829 4526
rect 842 4523 845 4553
rect 858 4533 861 4603
rect 938 4593 941 4616
rect 946 4603 965 4606
rect 834 4386 837 4516
rect 822 4383 837 4386
rect 794 4303 797 4326
rect 746 4193 749 4206
rect 654 4163 661 4166
rect 634 4113 637 4126
rect 642 4103 645 4126
rect 654 4086 657 4163
rect 674 4113 677 4126
rect 722 4086 725 4136
rect 770 4123 773 4276
rect 802 4273 805 4326
rect 810 4323 813 4336
rect 822 4316 825 4383
rect 818 4313 825 4316
rect 810 4226 813 4256
rect 786 4223 813 4226
rect 786 4213 789 4223
rect 778 4203 789 4206
rect 794 4203 797 4216
rect 786 4103 789 4136
rect 654 4083 661 4086
rect 722 4083 741 4086
rect 618 4033 629 4036
rect 610 3973 613 4016
rect 626 3966 629 4033
rect 610 3963 629 3966
rect 590 3903 597 3906
rect 590 3826 593 3903
rect 590 3823 597 3826
rect 594 3806 597 3823
rect 602 3813 605 3926
rect 610 3886 613 3963
rect 626 3933 629 3956
rect 642 3933 645 4006
rect 618 3913 621 3926
rect 610 3883 621 3886
rect 594 3803 613 3806
rect 538 3583 557 3586
rect 538 3473 541 3583
rect 546 3456 549 3526
rect 554 3523 557 3576
rect 562 3533 573 3536
rect 578 3533 581 3546
rect 570 3513 573 3526
rect 586 3486 589 3616
rect 594 3523 597 3736
rect 602 3596 605 3606
rect 610 3603 613 3803
rect 618 3796 621 3883
rect 618 3793 629 3796
rect 626 3656 629 3793
rect 626 3653 637 3656
rect 618 3596 621 3616
rect 626 3603 629 3646
rect 634 3613 637 3653
rect 602 3593 621 3596
rect 602 3523 605 3556
rect 610 3533 613 3566
rect 618 3533 621 3546
rect 610 3523 621 3526
rect 610 3503 613 3523
rect 626 3516 629 3596
rect 642 3573 645 3926
rect 658 3906 661 4083
rect 666 3923 669 3936
rect 698 3933 701 3976
rect 658 3903 669 3906
rect 666 3836 669 3903
rect 658 3833 669 3836
rect 658 3706 661 3833
rect 666 3793 669 3816
rect 698 3813 701 3926
rect 706 3923 709 4016
rect 714 3956 717 4046
rect 714 3953 725 3956
rect 722 3866 725 3953
rect 714 3863 725 3866
rect 738 3866 741 4083
rect 738 3863 749 3866
rect 658 3703 669 3706
rect 666 3626 669 3703
rect 682 3636 685 3746
rect 714 3736 717 3863
rect 746 3803 749 3863
rect 754 3843 757 4026
rect 770 3993 773 4006
rect 762 3923 765 3946
rect 770 3943 789 3946
rect 794 3943 797 4016
rect 802 4003 805 4136
rect 810 4123 813 4223
rect 818 4186 821 4313
rect 834 4223 837 4336
rect 842 4253 845 4326
rect 850 4303 853 4336
rect 858 4333 861 4526
rect 866 4523 869 4546
rect 898 4456 901 4536
rect 946 4523 949 4603
rect 954 4533 957 4546
rect 962 4513 965 4596
rect 978 4563 981 4626
rect 1042 4613 1045 4626
rect 1074 4613 1077 4636
rect 1082 4613 1085 4626
rect 898 4453 909 4456
rect 866 4323 869 4416
rect 906 4376 909 4453
rect 922 4393 925 4406
rect 898 4373 909 4376
rect 882 4293 885 4326
rect 898 4256 901 4373
rect 906 4343 925 4346
rect 906 4333 909 4343
rect 898 4253 905 4256
rect 834 4186 837 4206
rect 818 4183 837 4186
rect 834 4166 837 4183
rect 834 4163 845 4166
rect 818 4036 821 4136
rect 842 4036 845 4163
rect 866 4123 869 4216
rect 902 4176 905 4253
rect 898 4173 905 4176
rect 898 4136 901 4173
rect 898 4133 905 4136
rect 890 4063 893 4126
rect 902 4046 905 4133
rect 902 4043 909 4046
rect 810 4033 821 4036
rect 834 4033 845 4036
rect 834 3993 837 4033
rect 770 3933 773 3943
rect 770 3893 773 3926
rect 778 3903 781 3936
rect 786 3923 789 3943
rect 802 3893 805 3986
rect 850 3956 853 4016
rect 842 3953 853 3956
rect 842 3933 845 3953
rect 762 3813 765 3826
rect 778 3793 781 3806
rect 714 3733 725 3736
rect 682 3633 693 3636
rect 666 3623 677 3626
rect 666 3553 669 3606
rect 618 3513 629 3516
rect 642 3533 661 3536
rect 586 3483 597 3486
rect 546 3453 557 3456
rect 554 3436 557 3453
rect 554 3433 561 3436
rect 474 3413 477 3426
rect 514 3413 517 3426
rect 458 3323 461 3406
rect 474 3323 477 3356
rect 482 3313 485 3376
rect 450 3303 461 3306
rect 458 3246 461 3303
rect 490 3256 493 3406
rect 514 3333 517 3346
rect 522 3316 525 3396
rect 558 3376 561 3433
rect 554 3373 561 3376
rect 450 3243 461 3246
rect 482 3253 493 3256
rect 514 3313 525 3316
rect 402 3193 421 3196
rect 450 3186 453 3243
rect 442 3183 453 3186
rect 394 3053 405 3056
rect 402 3013 405 3053
rect 410 3003 413 3026
rect 418 3003 421 3156
rect 442 3036 445 3183
rect 442 3033 453 3036
rect 338 2943 349 2946
rect 298 2903 317 2906
rect 274 2823 285 2826
rect 274 2803 277 2823
rect 282 2793 285 2816
rect 298 2813 301 2886
rect 238 2713 245 2716
rect 250 2713 253 2726
rect 218 2693 229 2696
rect 66 2546 69 2586
rect 82 2566 85 2653
rect 82 2563 93 2566
rect 66 2543 77 2546
rect 74 2486 77 2543
rect 66 2483 77 2486
rect 66 1696 69 2483
rect 90 2466 93 2563
rect 122 2536 125 2693
rect 130 2613 133 2626
rect 162 2613 165 2636
rect 170 2613 173 2626
rect 178 2556 181 2616
rect 186 2596 189 2606
rect 194 2603 197 2636
rect 202 2596 205 2616
rect 186 2593 205 2596
rect 154 2553 181 2556
rect 122 2533 133 2536
rect 82 2463 93 2466
rect 82 2413 85 2463
rect 114 2413 117 2526
rect 130 2466 133 2533
rect 122 2463 133 2466
rect 82 2176 85 2406
rect 122 2396 125 2463
rect 154 2453 157 2553
rect 162 2543 181 2546
rect 162 2533 165 2543
rect 170 2466 173 2536
rect 178 2523 181 2543
rect 162 2463 173 2466
rect 154 2396 157 2416
rect 162 2413 165 2463
rect 114 2393 125 2396
rect 150 2393 157 2396
rect 114 2316 117 2393
rect 130 2323 133 2386
rect 150 2316 153 2393
rect 162 2323 165 2376
rect 114 2313 125 2316
rect 150 2313 157 2316
rect 82 2173 93 2176
rect 90 1993 93 2173
rect 90 1836 93 1936
rect 122 1846 125 2313
rect 130 2213 133 2226
rect 154 2126 157 2313
rect 170 2236 173 2456
rect 194 2416 197 2536
rect 210 2533 213 2606
rect 218 2533 221 2606
rect 226 2603 229 2693
rect 238 2626 241 2713
rect 258 2696 261 2736
rect 266 2723 269 2736
rect 282 2733 285 2746
rect 306 2723 309 2736
rect 314 2716 317 2903
rect 346 2896 349 2943
rect 362 2913 365 2926
rect 394 2903 397 2926
rect 402 2913 405 2926
rect 442 2923 445 3016
rect 338 2893 349 2896
rect 330 2723 333 2806
rect 338 2786 341 2893
rect 354 2793 357 2806
rect 338 2783 349 2786
rect 346 2746 349 2783
rect 346 2743 353 2746
rect 306 2713 317 2716
rect 234 2623 241 2626
rect 234 2593 237 2623
rect 242 2503 245 2526
rect 178 2383 181 2416
rect 194 2413 205 2416
rect 178 2333 181 2376
rect 186 2323 189 2406
rect 202 2366 205 2413
rect 226 2393 229 2406
rect 194 2363 205 2366
rect 194 2276 197 2363
rect 218 2333 221 2346
rect 250 2343 253 2696
rect 258 2693 277 2696
rect 258 2583 261 2646
rect 274 2613 277 2693
rect 282 2603 285 2626
rect 290 2613 293 2636
rect 298 2603 301 2616
rect 306 2573 309 2713
rect 350 2686 353 2743
rect 346 2683 353 2686
rect 314 2553 317 2606
rect 330 2576 333 2606
rect 346 2593 349 2683
rect 362 2623 365 2726
rect 386 2723 389 2816
rect 394 2706 397 2796
rect 410 2743 429 2746
rect 410 2733 413 2743
rect 390 2703 397 2706
rect 390 2636 393 2703
rect 390 2633 397 2636
rect 322 2573 333 2576
rect 314 2533 317 2546
rect 258 2413 261 2526
rect 314 2513 317 2526
rect 322 2413 325 2573
rect 330 2523 333 2546
rect 346 2493 349 2536
rect 354 2533 357 2546
rect 362 2406 365 2616
rect 394 2613 397 2633
rect 402 2543 405 2726
rect 410 2713 413 2726
rect 418 2723 421 2736
rect 426 2723 429 2743
rect 434 2733 437 2816
rect 442 2616 445 2806
rect 450 2766 453 3033
rect 458 3013 461 3026
rect 466 3003 469 3206
rect 474 3113 477 3136
rect 482 3106 485 3253
rect 514 3236 517 3313
rect 514 3233 525 3236
rect 506 3123 509 3216
rect 522 3116 525 3233
rect 530 3213 533 3326
rect 546 3176 549 3336
rect 538 3173 549 3176
rect 538 3126 541 3173
rect 546 3133 549 3146
rect 538 3123 549 3126
rect 522 3113 533 3116
rect 482 3103 493 3106
rect 458 2943 477 2946
rect 458 2933 461 2943
rect 466 2903 469 2936
rect 474 2923 477 2943
rect 482 2933 485 3006
rect 490 2996 493 3103
rect 514 3013 517 3026
rect 490 2993 501 2996
rect 498 2926 501 2993
rect 490 2923 501 2926
rect 490 2853 493 2923
rect 466 2793 469 2806
rect 450 2763 461 2766
rect 458 2666 461 2763
rect 490 2713 493 2816
rect 514 2813 517 2926
rect 522 2923 525 3006
rect 530 2856 533 3113
rect 546 3103 549 3123
rect 538 2933 541 3016
rect 530 2853 537 2856
rect 534 2766 537 2853
rect 546 2813 549 3006
rect 554 2806 557 3373
rect 570 3346 573 3416
rect 578 3413 581 3476
rect 594 3396 597 3483
rect 586 3393 597 3396
rect 586 3373 589 3393
rect 562 3343 573 3346
rect 562 3223 565 3343
rect 570 3313 573 3336
rect 586 3333 589 3356
rect 618 3336 621 3513
rect 642 3496 645 3533
rect 638 3493 645 3496
rect 638 3426 641 3493
rect 650 3433 653 3526
rect 666 3483 669 3526
rect 626 3413 629 3426
rect 638 3423 645 3426
rect 642 3403 645 3423
rect 618 3333 625 3336
rect 610 3286 613 3326
rect 602 3283 613 3286
rect 562 3143 565 3216
rect 570 3203 573 3216
rect 602 3213 605 3283
rect 622 3276 625 3333
rect 618 3273 625 3276
rect 610 3203 613 3226
rect 570 3133 573 3196
rect 562 3113 565 3126
rect 562 3013 565 3106
rect 578 3023 581 3126
rect 618 3123 621 3273
rect 626 3193 629 3206
rect 634 3123 637 3396
rect 666 3313 669 3406
rect 674 3393 677 3623
rect 690 3566 693 3633
rect 706 3613 709 3726
rect 722 3606 725 3733
rect 770 3706 773 3726
rect 762 3703 773 3706
rect 762 3646 765 3703
rect 786 3656 789 3846
rect 810 3813 813 3916
rect 818 3893 821 3926
rect 850 3886 853 3906
rect 842 3883 853 3886
rect 818 3806 821 3846
rect 826 3813 829 3856
rect 842 3836 845 3883
rect 858 3843 861 3996
rect 842 3833 853 3836
rect 802 3763 805 3806
rect 810 3803 821 3806
rect 810 3733 813 3803
rect 834 3733 837 3816
rect 786 3653 793 3656
rect 762 3643 773 3646
rect 682 3563 693 3566
rect 714 3603 725 3606
rect 682 3533 685 3563
rect 690 3493 693 3546
rect 682 3333 685 3486
rect 714 3483 717 3603
rect 722 3493 725 3536
rect 706 3413 709 3456
rect 722 3413 725 3476
rect 730 3413 733 3536
rect 746 3523 749 3606
rect 762 3603 765 3626
rect 770 3563 773 3643
rect 778 3533 781 3646
rect 790 3526 793 3653
rect 826 3613 829 3666
rect 834 3613 837 3726
rect 842 3703 845 3806
rect 850 3776 853 3833
rect 858 3793 861 3816
rect 850 3773 857 3776
rect 854 3686 857 3773
rect 854 3683 869 3686
rect 842 3613 845 3676
rect 802 3583 805 3606
rect 858 3596 861 3606
rect 866 3603 869 3683
rect 874 3643 877 3896
rect 882 3683 885 4006
rect 906 3986 909 4043
rect 902 3983 909 3986
rect 902 3926 905 3983
rect 914 3966 917 4336
rect 922 4323 925 4343
rect 930 4333 933 4416
rect 986 4413 989 4536
rect 994 4503 997 4606
rect 1090 4603 1093 4616
rect 1098 4596 1101 4606
rect 1106 4603 1109 4636
rect 1114 4596 1117 4616
rect 1122 4603 1125 4616
rect 1130 4613 1133 4646
rect 1130 4596 1133 4606
rect 1098 4593 1117 4596
rect 1122 4593 1133 4596
rect 1106 4536 1109 4556
rect 1002 4513 1005 4526
rect 1018 4503 1021 4536
rect 1090 4533 1109 4536
rect 1042 4413 1045 4426
rect 1050 4413 1053 4526
rect 970 4386 973 4406
rect 962 4383 973 4386
rect 978 4383 981 4396
rect 938 4323 941 4336
rect 962 4236 965 4383
rect 962 4233 973 4236
rect 922 4193 925 4226
rect 970 4216 973 4233
rect 946 4196 949 4216
rect 970 4213 977 4216
rect 946 4193 957 4196
rect 962 4193 965 4206
rect 954 4186 957 4193
rect 954 4183 965 4186
rect 938 4143 957 4146
rect 938 4133 941 4143
rect 946 4123 949 4136
rect 954 4123 957 4143
rect 962 4123 965 4183
rect 974 4156 977 4213
rect 970 4153 977 4156
rect 970 4106 973 4153
rect 986 4146 989 4406
rect 1018 4343 1021 4356
rect 994 4313 997 4326
rect 1010 4236 1013 4336
rect 1002 4233 1013 4236
rect 1002 4213 1005 4233
rect 1034 4216 1037 4336
rect 1050 4313 1053 4366
rect 1058 4356 1061 4416
rect 1082 4396 1085 4406
rect 1090 4403 1093 4533
rect 1098 4446 1101 4526
rect 1106 4483 1109 4526
rect 1122 4523 1125 4593
rect 1098 4443 1109 4446
rect 1098 4396 1101 4416
rect 1082 4393 1101 4396
rect 1058 4353 1065 4356
rect 1062 4286 1065 4353
rect 1082 4316 1085 4336
rect 1106 4333 1109 4443
rect 1138 4436 1141 4606
rect 1146 4513 1149 4686
rect 1154 4553 1157 4616
rect 1162 4476 1165 4546
rect 1170 4533 1173 4636
rect 1178 4613 1181 4626
rect 1186 4543 1189 4616
rect 1218 4613 1221 4626
rect 1266 4593 1269 4606
rect 1306 4593 1309 4606
rect 1354 4603 1357 4616
rect 1386 4586 1389 4616
rect 1378 4583 1389 4586
rect 1162 4473 1173 4476
rect 1130 4433 1141 4436
rect 1114 4393 1125 4396
rect 1122 4323 1125 4346
rect 1130 4333 1133 4433
rect 1154 4373 1157 4406
rect 1162 4403 1165 4416
rect 1170 4403 1173 4473
rect 1202 4423 1205 4536
rect 1210 4523 1213 4536
rect 1266 4533 1269 4556
rect 1274 4533 1277 4566
rect 1306 4533 1309 4546
rect 1226 4513 1229 4526
rect 1058 4283 1065 4286
rect 1058 4263 1061 4283
rect 1034 4213 1045 4216
rect 986 4143 993 4146
rect 962 4103 973 4106
rect 914 3963 925 3966
rect 890 3906 893 3926
rect 902 3923 909 3926
rect 890 3903 897 3906
rect 894 3836 897 3903
rect 890 3833 897 3836
rect 890 3813 893 3833
rect 906 3816 909 3923
rect 922 3903 925 3963
rect 930 3933 933 4016
rect 962 3976 965 4103
rect 978 4013 981 4136
rect 978 3993 981 4006
rect 990 3986 993 4143
rect 986 3983 993 3986
rect 962 3973 969 3976
rect 946 3943 949 3956
rect 898 3813 909 3816
rect 930 3813 933 3926
rect 890 3783 893 3806
rect 898 3736 901 3813
rect 906 3793 909 3806
rect 914 3793 917 3806
rect 898 3733 905 3736
rect 890 3676 893 3726
rect 882 3673 893 3676
rect 874 3596 877 3616
rect 858 3593 877 3596
rect 882 3583 885 3673
rect 890 3613 893 3646
rect 902 3636 905 3733
rect 898 3633 905 3636
rect 898 3596 901 3633
rect 906 3603 909 3616
rect 914 3613 917 3696
rect 898 3593 909 3596
rect 802 3533 805 3556
rect 818 3533 821 3566
rect 826 3533 829 3546
rect 714 3393 717 3406
rect 722 3403 733 3406
rect 738 3376 741 3496
rect 754 3436 757 3526
rect 786 3523 793 3526
rect 786 3466 789 3523
rect 778 3463 789 3466
rect 754 3433 765 3436
rect 722 3373 741 3376
rect 722 3266 725 3373
rect 722 3263 741 3266
rect 642 3203 645 3236
rect 690 3203 693 3226
rect 642 3133 645 3146
rect 666 3133 669 3146
rect 674 3136 677 3156
rect 674 3133 685 3136
rect 634 3013 637 3026
rect 570 2933 589 2936
rect 562 2906 565 2926
rect 562 2903 573 2906
rect 570 2836 573 2903
rect 562 2833 573 2836
rect 562 2813 565 2833
rect 586 2813 589 2933
rect 594 2903 597 3006
rect 642 2973 645 3006
rect 602 2913 605 2926
rect 530 2763 537 2766
rect 546 2803 557 2806
rect 530 2746 533 2763
rect 514 2733 517 2746
rect 522 2743 533 2746
rect 522 2733 525 2743
rect 450 2663 461 2666
rect 506 2666 509 2726
rect 522 2693 525 2726
rect 530 2703 533 2736
rect 506 2663 517 2666
rect 450 2643 453 2663
rect 410 2533 413 2616
rect 434 2613 445 2616
rect 458 2613 461 2626
rect 466 2613 469 2646
rect 370 2496 373 2526
rect 378 2513 381 2526
rect 426 2513 429 2536
rect 434 2496 437 2613
rect 450 2546 453 2606
rect 442 2543 453 2546
rect 442 2533 445 2543
rect 370 2493 381 2496
rect 378 2436 381 2493
rect 370 2433 381 2436
rect 426 2493 437 2496
rect 426 2436 429 2493
rect 426 2433 437 2436
rect 370 2413 373 2433
rect 434 2416 437 2433
rect 426 2413 437 2416
rect 338 2366 341 2406
rect 362 2403 373 2406
rect 330 2363 341 2366
rect 314 2333 317 2356
rect 202 2283 205 2326
rect 266 2313 269 2326
rect 298 2303 301 2326
rect 306 2313 309 2326
rect 194 2273 213 2276
rect 162 2213 165 2236
rect 170 2233 181 2236
rect 170 2213 173 2226
rect 178 2193 181 2233
rect 186 2196 189 2206
rect 194 2203 197 2236
rect 202 2196 205 2216
rect 186 2193 205 2196
rect 138 2113 141 2126
rect 154 2123 165 2126
rect 170 2123 173 2136
rect 138 2013 141 2026
rect 162 1936 165 2123
rect 178 2113 181 2126
rect 194 2113 197 2136
rect 202 2036 205 2126
rect 210 2046 213 2273
rect 330 2226 333 2363
rect 306 2223 333 2226
rect 218 2173 221 2206
rect 234 2203 237 2216
rect 218 2133 229 2136
rect 218 2113 221 2126
rect 226 2123 229 2133
rect 210 2043 229 2046
rect 170 2013 173 2036
rect 194 2033 205 2036
rect 178 2013 181 2026
rect 194 1936 197 2033
rect 202 2013 205 2026
rect 202 1996 205 2006
rect 210 2003 213 2036
rect 218 1996 221 2016
rect 226 2003 229 2043
rect 234 2023 237 2196
rect 242 2156 245 2176
rect 242 2153 253 2156
rect 250 2076 253 2153
rect 274 2123 277 2216
rect 282 2113 285 2126
rect 242 2073 253 2076
rect 202 1993 221 1996
rect 158 1933 165 1936
rect 190 1933 197 1936
rect 210 1943 229 1946
rect 210 1933 213 1943
rect 138 1913 141 1926
rect 158 1876 161 1933
rect 170 1903 173 1926
rect 178 1913 181 1926
rect 158 1873 165 1876
rect 122 1843 133 1846
rect 82 1833 93 1836
rect 82 1766 85 1833
rect 82 1763 93 1766
rect 98 1763 101 1806
rect 130 1796 133 1843
rect 146 1813 149 1826
rect 122 1793 133 1796
rect 66 1693 77 1696
rect 74 1586 77 1693
rect 66 1583 77 1586
rect 66 1423 69 1583
rect 90 1566 93 1763
rect 122 1736 125 1793
rect 162 1776 165 1873
rect 190 1846 193 1933
rect 202 1856 205 1926
rect 218 1903 221 1936
rect 226 1923 229 1943
rect 202 1853 209 1856
rect 190 1843 197 1846
rect 154 1773 165 1776
rect 154 1746 157 1773
rect 154 1743 161 1746
rect 122 1733 133 1736
rect 114 1613 117 1726
rect 130 1606 133 1733
rect 158 1686 161 1743
rect 178 1733 181 1816
rect 186 1813 189 1826
rect 194 1796 197 1843
rect 190 1793 197 1796
rect 154 1683 161 1686
rect 82 1563 93 1566
rect 122 1603 133 1606
rect 66 996 69 1416
rect 82 1403 85 1563
rect 82 1133 85 1396
rect 106 1323 109 1416
rect 74 1003 77 1026
rect 82 1013 85 1116
rect 106 1113 109 1126
rect 90 1013 93 1036
rect 122 1016 125 1603
rect 130 1513 133 1526
rect 146 1433 149 1616
rect 154 1576 157 1683
rect 162 1613 165 1626
rect 162 1596 165 1606
rect 170 1603 173 1726
rect 178 1623 181 1726
rect 190 1716 193 1793
rect 206 1786 209 1853
rect 218 1803 229 1806
rect 202 1783 209 1786
rect 202 1723 205 1783
rect 218 1723 221 1796
rect 234 1776 237 1936
rect 242 1933 245 2073
rect 250 2013 253 2056
rect 250 1916 253 1996
rect 246 1913 253 1916
rect 246 1826 249 1913
rect 258 1833 261 1926
rect 266 1906 269 2016
rect 282 1993 285 2006
rect 306 1983 309 2223
rect 322 2136 325 2216
rect 330 2213 333 2223
rect 314 2126 317 2136
rect 322 2133 333 2136
rect 314 2123 333 2126
rect 338 2043 341 2146
rect 370 2136 373 2403
rect 378 2313 381 2326
rect 410 2323 413 2366
rect 418 2313 421 2326
rect 362 2133 373 2136
rect 362 2066 365 2133
rect 362 2063 373 2066
rect 266 1903 277 1906
rect 274 1846 277 1903
rect 290 1853 293 1936
rect 298 1933 301 1946
rect 330 1923 333 1946
rect 338 1923 341 2016
rect 370 2003 373 2063
rect 266 1843 277 1846
rect 246 1823 253 1826
rect 226 1773 237 1776
rect 250 1776 253 1823
rect 266 1813 269 1843
rect 378 1836 381 2126
rect 394 2066 397 2156
rect 402 2123 405 2206
rect 418 2203 421 2216
rect 394 2063 405 2066
rect 386 2013 389 2026
rect 394 2013 397 2056
rect 402 2003 405 2063
rect 410 1933 413 2016
rect 418 1993 421 2026
rect 426 2013 429 2413
rect 442 2406 445 2526
rect 450 2523 453 2536
rect 482 2533 485 2616
rect 490 2603 493 2626
rect 498 2613 501 2636
rect 514 2613 517 2663
rect 498 2516 501 2596
rect 450 2413 453 2516
rect 490 2513 501 2516
rect 466 2413 469 2506
rect 490 2436 493 2513
rect 490 2433 501 2436
rect 434 2393 437 2406
rect 442 2403 461 2406
rect 434 2333 437 2346
rect 434 2173 437 2326
rect 442 2306 445 2403
rect 450 2323 453 2356
rect 442 2303 449 2306
rect 446 2176 449 2303
rect 458 2203 461 2336
rect 466 2243 469 2326
rect 474 2316 477 2416
rect 498 2413 501 2433
rect 482 2333 485 2406
rect 506 2383 509 2406
rect 490 2323 493 2346
rect 498 2323 501 2336
rect 474 2313 481 2316
rect 478 2236 481 2313
rect 474 2233 481 2236
rect 466 2213 469 2226
rect 474 2213 477 2233
rect 490 2213 493 2316
rect 506 2283 509 2326
rect 514 2313 517 2576
rect 530 2413 533 2616
rect 546 2596 549 2803
rect 562 2626 565 2696
rect 570 2673 573 2806
rect 578 2783 581 2806
rect 594 2636 597 2806
rect 618 2803 621 2936
rect 650 2933 653 3126
rect 666 3123 677 3126
rect 674 3023 677 3123
rect 682 3096 685 3126
rect 682 3093 689 3096
rect 686 3016 689 3093
rect 698 3066 701 3136
rect 722 3123 725 3216
rect 698 3063 717 3066
rect 682 3013 689 3016
rect 666 2963 669 3006
rect 682 2966 685 3013
rect 682 2963 689 2966
rect 642 2913 645 2926
rect 686 2896 689 2963
rect 682 2893 689 2896
rect 682 2876 685 2893
rect 674 2873 685 2876
rect 626 2793 629 2816
rect 674 2756 677 2873
rect 698 2836 701 2926
rect 714 2896 717 3063
rect 730 3043 733 3246
rect 738 3106 741 3263
rect 746 3123 749 3416
rect 762 3366 765 3433
rect 754 3363 765 3366
rect 754 3343 757 3363
rect 778 3336 781 3463
rect 762 3333 781 3336
rect 762 3246 765 3333
rect 794 3306 797 3456
rect 810 3443 813 3526
rect 850 3496 853 3536
rect 890 3523 893 3576
rect 906 3556 909 3593
rect 902 3553 909 3556
rect 902 3506 905 3553
rect 922 3543 925 3806
rect 938 3746 941 3816
rect 954 3783 957 3926
rect 966 3776 969 3973
rect 966 3773 973 3776
rect 934 3743 941 3746
rect 962 3743 965 3756
rect 934 3686 937 3743
rect 934 3683 941 3686
rect 938 3663 941 3683
rect 946 3613 949 3736
rect 902 3503 909 3506
rect 842 3493 853 3496
rect 810 3393 821 3396
rect 842 3376 845 3493
rect 906 3486 909 3503
rect 922 3493 925 3536
rect 946 3496 949 3546
rect 954 3523 957 3726
rect 962 3613 965 3646
rect 970 3596 973 3773
rect 978 3663 981 3936
rect 966 3593 973 3596
rect 938 3493 949 3496
rect 842 3373 849 3376
rect 754 3243 765 3246
rect 786 3303 797 3306
rect 786 3246 789 3303
rect 786 3243 797 3246
rect 754 3176 757 3243
rect 770 3213 773 3226
rect 762 3183 765 3206
rect 754 3173 765 3176
rect 762 3156 765 3173
rect 762 3153 769 3156
rect 738 3103 745 3106
rect 742 3036 745 3103
rect 766 3086 769 3153
rect 778 3123 781 3206
rect 786 3096 789 3206
rect 794 3173 797 3243
rect 802 3213 805 3306
rect 818 3303 821 3336
rect 846 3276 849 3373
rect 858 3313 861 3326
rect 842 3273 849 3276
rect 842 3216 845 3273
rect 842 3213 853 3216
rect 762 3083 769 3086
rect 778 3093 789 3096
rect 762 3056 765 3083
rect 738 3033 745 3036
rect 758 3053 765 3056
rect 730 2933 733 2966
rect 690 2833 701 2836
rect 706 2893 717 2896
rect 690 2803 693 2833
rect 706 2803 709 2893
rect 674 2753 685 2756
rect 594 2633 605 2636
rect 562 2623 589 2626
rect 562 2613 565 2623
rect 554 2603 565 2606
rect 570 2603 573 2616
rect 546 2593 557 2596
rect 530 2373 533 2406
rect 538 2313 541 2336
rect 522 2236 525 2246
rect 482 2193 485 2206
rect 498 2203 501 2236
rect 518 2233 525 2236
rect 442 2173 449 2176
rect 442 2153 445 2173
rect 434 2133 437 2146
rect 442 2113 445 2136
rect 458 2133 461 2156
rect 506 2143 509 2216
rect 518 2156 521 2233
rect 538 2213 541 2226
rect 514 2153 521 2156
rect 450 2076 453 2126
rect 458 2093 461 2126
rect 474 2113 477 2126
rect 514 2123 517 2153
rect 522 2133 533 2136
rect 538 2133 541 2156
rect 546 2133 549 2186
rect 554 2153 557 2593
rect 586 2586 589 2623
rect 578 2583 589 2586
rect 578 2536 581 2583
rect 602 2566 605 2633
rect 618 2613 621 2726
rect 674 2723 677 2736
rect 682 2706 685 2753
rect 690 2733 693 2786
rect 706 2733 717 2736
rect 722 2733 725 2796
rect 674 2703 685 2706
rect 674 2636 677 2703
rect 690 2643 693 2726
rect 674 2633 685 2636
rect 594 2563 605 2566
rect 594 2543 597 2563
rect 578 2533 589 2536
rect 642 2533 645 2546
rect 562 2393 565 2406
rect 578 2403 581 2476
rect 586 2413 589 2533
rect 666 2523 669 2616
rect 674 2603 677 2616
rect 682 2596 685 2633
rect 706 2613 709 2726
rect 714 2683 717 2733
rect 730 2723 733 2816
rect 738 2706 741 3033
rect 746 2923 749 3016
rect 758 2996 761 3053
rect 758 2993 765 2996
rect 762 2976 765 2993
rect 754 2943 757 2976
rect 762 2973 773 2976
rect 770 2926 773 2973
rect 762 2923 773 2926
rect 762 2866 765 2923
rect 762 2863 773 2866
rect 746 2766 749 2786
rect 770 2766 773 2863
rect 746 2763 757 2766
rect 730 2703 741 2706
rect 730 2626 733 2703
rect 754 2696 757 2763
rect 746 2693 757 2696
rect 766 2763 773 2766
rect 730 2623 737 2626
rect 678 2593 685 2596
rect 678 2516 681 2593
rect 674 2513 681 2516
rect 602 2403 605 2426
rect 610 2356 613 2406
rect 602 2353 613 2356
rect 602 2333 605 2353
rect 586 2303 589 2326
rect 594 2293 597 2326
rect 610 2313 613 2326
rect 626 2323 629 2426
rect 642 2413 645 2496
rect 642 2393 645 2406
rect 658 2366 661 2416
rect 674 2406 677 2513
rect 690 2486 693 2606
rect 722 2526 725 2606
rect 734 2556 737 2623
rect 734 2553 741 2556
rect 706 2523 725 2526
rect 706 2506 709 2523
rect 706 2503 713 2506
rect 690 2483 701 2486
rect 674 2403 681 2406
rect 650 2363 661 2366
rect 634 2333 637 2356
rect 650 2286 653 2363
rect 678 2346 681 2403
rect 678 2343 685 2346
rect 674 2303 677 2326
rect 650 2283 661 2286
rect 658 2243 661 2283
rect 586 2203 589 2216
rect 562 2133 565 2146
rect 450 2073 469 2076
rect 466 2013 469 2073
rect 378 1833 389 1836
rect 250 1773 261 1776
rect 190 1713 197 1716
rect 178 1596 181 1616
rect 162 1593 181 1596
rect 154 1573 161 1576
rect 158 1436 161 1573
rect 154 1433 161 1436
rect 146 1256 149 1426
rect 154 1393 157 1433
rect 162 1396 165 1416
rect 170 1413 173 1516
rect 186 1493 189 1646
rect 194 1613 197 1713
rect 226 1643 229 1773
rect 234 1703 237 1726
rect 194 1513 197 1526
rect 178 1403 181 1426
rect 186 1413 189 1436
rect 210 1426 213 1616
rect 242 1613 245 1726
rect 258 1666 261 1773
rect 254 1663 261 1666
rect 254 1606 257 1663
rect 282 1613 285 1816
rect 330 1813 333 1826
rect 306 1636 309 1736
rect 314 1713 317 1736
rect 330 1733 333 1766
rect 322 1723 333 1726
rect 338 1713 341 1726
rect 346 1676 349 1726
rect 338 1673 349 1676
rect 306 1633 333 1636
rect 250 1603 257 1606
rect 298 1603 301 1616
rect 306 1613 309 1626
rect 194 1423 213 1426
rect 186 1396 189 1406
rect 162 1393 189 1396
rect 178 1333 181 1366
rect 178 1306 181 1326
rect 170 1303 181 1306
rect 170 1256 173 1303
rect 146 1253 153 1256
rect 170 1253 181 1256
rect 130 1213 133 1226
rect 150 1196 153 1253
rect 162 1213 165 1236
rect 170 1213 173 1226
rect 150 1193 157 1196
rect 154 1086 157 1193
rect 170 1106 173 1126
rect 66 993 85 996
rect 82 506 85 993
rect 98 913 101 1006
rect 106 933 109 1016
rect 118 1013 125 1016
rect 146 1083 157 1086
rect 166 1103 173 1106
rect 118 946 121 1013
rect 118 943 125 946
rect 114 906 117 926
rect 110 903 117 906
rect 110 836 113 903
rect 110 833 117 836
rect 114 813 117 833
rect 122 626 125 943
rect 130 933 133 1006
rect 146 1003 149 1083
rect 166 1036 169 1103
rect 146 856 149 936
rect 154 923 157 1036
rect 166 1033 173 1036
rect 178 1033 181 1253
rect 194 1246 197 1423
rect 202 1363 205 1416
rect 210 1413 221 1416
rect 210 1373 213 1413
rect 218 1276 221 1406
rect 226 1333 229 1436
rect 234 1403 237 1526
rect 250 1503 253 1603
rect 258 1513 261 1526
rect 290 1523 293 1536
rect 298 1513 301 1526
rect 242 1413 245 1426
rect 250 1383 253 1496
rect 266 1413 269 1446
rect 234 1326 237 1346
rect 290 1343 293 1506
rect 306 1443 309 1526
rect 314 1513 317 1536
rect 322 1426 325 1616
rect 330 1613 333 1633
rect 338 1606 341 1673
rect 354 1613 357 1796
rect 362 1733 365 1816
rect 370 1813 373 1826
rect 370 1723 373 1806
rect 386 1786 389 1833
rect 418 1803 421 1826
rect 426 1813 429 2006
rect 442 1983 445 2006
rect 514 1936 517 2066
rect 522 2013 525 2126
rect 530 2003 533 2126
rect 538 2016 541 2126
rect 546 2063 549 2126
rect 538 2013 549 2016
rect 554 2013 557 2126
rect 570 2123 573 2136
rect 546 1983 549 2006
rect 562 2003 565 2026
rect 570 1993 573 2006
rect 514 1933 525 1936
rect 450 1813 453 1926
rect 474 1813 477 1826
rect 458 1793 461 1806
rect 386 1783 397 1786
rect 466 1783 469 1806
rect 330 1603 341 1606
rect 330 1533 341 1536
rect 330 1513 333 1526
rect 346 1516 349 1606
rect 354 1523 357 1536
rect 346 1513 357 1516
rect 362 1513 365 1616
rect 378 1613 381 1776
rect 386 1733 389 1756
rect 394 1726 397 1783
rect 482 1773 485 1886
rect 490 1813 493 1836
rect 426 1726 429 1756
rect 434 1733 445 1736
rect 450 1733 453 1746
rect 386 1723 397 1726
rect 386 1703 389 1723
rect 386 1556 389 1576
rect 378 1553 389 1556
rect 354 1456 357 1513
rect 354 1453 361 1456
rect 322 1423 333 1426
rect 282 1333 293 1336
rect 298 1333 301 1376
rect 314 1346 317 1416
rect 330 1356 333 1423
rect 358 1396 361 1453
rect 378 1436 381 1553
rect 402 1546 405 1726
rect 418 1723 429 1726
rect 442 1643 445 1726
rect 490 1706 493 1806
rect 498 1803 501 1906
rect 506 1783 509 1926
rect 522 1846 525 1933
rect 546 1923 549 1976
rect 578 1973 581 2156
rect 602 2146 605 2216
rect 626 2206 629 2226
rect 618 2203 629 2206
rect 634 2203 637 2216
rect 658 2213 661 2226
rect 594 2143 605 2146
rect 594 2096 597 2143
rect 610 2103 613 2136
rect 626 2103 629 2126
rect 594 2093 605 2096
rect 602 2046 605 2093
rect 598 2043 605 2046
rect 598 1996 601 2043
rect 618 2016 621 2096
rect 610 2013 621 2016
rect 610 2003 621 2006
rect 626 2003 629 2036
rect 634 2013 637 2046
rect 642 2013 645 2136
rect 650 2133 653 2206
rect 658 2193 669 2196
rect 658 2026 661 2156
rect 666 2113 669 2126
rect 654 2023 661 2026
rect 598 1993 605 1996
rect 602 1943 605 1993
rect 522 1843 533 1846
rect 530 1766 533 1843
rect 530 1763 541 1766
rect 506 1743 525 1746
rect 506 1733 509 1743
rect 498 1713 501 1726
rect 506 1706 509 1726
rect 490 1703 509 1706
rect 394 1543 405 1546
rect 418 1546 421 1616
rect 418 1543 429 1546
rect 378 1433 389 1436
rect 354 1393 361 1396
rect 354 1376 357 1393
rect 306 1343 317 1346
rect 322 1353 333 1356
rect 346 1373 357 1376
rect 186 1243 197 1246
rect 210 1273 221 1276
rect 186 1213 189 1243
rect 186 1196 189 1206
rect 194 1203 197 1236
rect 202 1196 205 1216
rect 186 1193 205 1196
rect 186 1096 189 1166
rect 186 1093 193 1096
rect 170 1003 173 1033
rect 190 1026 193 1093
rect 178 1013 181 1026
rect 186 1023 193 1026
rect 186 993 189 1023
rect 202 946 205 1186
rect 210 1163 213 1273
rect 226 1213 229 1326
rect 234 1323 241 1326
rect 282 1323 301 1326
rect 306 1323 309 1343
rect 238 1226 241 1323
rect 234 1223 241 1226
rect 234 1206 237 1223
rect 258 1213 269 1216
rect 258 1206 261 1213
rect 226 1203 237 1206
rect 250 1203 261 1206
rect 226 1096 229 1203
rect 274 1196 277 1206
rect 282 1203 285 1216
rect 290 1196 293 1216
rect 298 1203 301 1323
rect 274 1193 293 1196
rect 218 1093 229 1096
rect 202 943 213 946
rect 146 853 153 856
rect 150 796 153 853
rect 162 813 165 916
rect 170 906 173 926
rect 170 903 181 906
rect 186 903 189 936
rect 146 793 153 796
rect 146 773 149 793
rect 130 713 133 726
rect 162 723 165 746
rect 170 713 173 726
rect 178 636 181 903
rect 210 843 213 943
rect 202 813 205 826
rect 194 793 197 806
rect 218 783 221 1093
rect 226 1013 229 1026
rect 234 1013 237 1126
rect 306 1106 309 1126
rect 298 1103 309 1106
rect 250 1013 253 1026
rect 282 1013 285 1056
rect 298 1046 301 1103
rect 298 1043 309 1046
rect 282 996 285 1006
rect 290 1003 293 1026
rect 298 996 301 1016
rect 306 1003 309 1043
rect 282 993 301 996
rect 314 956 317 1216
rect 322 1196 325 1353
rect 330 1323 333 1336
rect 346 1213 349 1373
rect 370 1366 373 1416
rect 378 1393 381 1406
rect 386 1386 389 1433
rect 394 1426 397 1543
rect 402 1433 405 1536
rect 410 1533 421 1536
rect 394 1423 405 1426
rect 362 1363 373 1366
rect 378 1383 389 1386
rect 362 1333 365 1363
rect 354 1196 357 1216
rect 362 1203 365 1326
rect 378 1286 381 1383
rect 402 1346 405 1423
rect 418 1416 421 1526
rect 426 1523 429 1543
rect 418 1413 429 1416
rect 410 1393 413 1406
rect 418 1403 429 1406
rect 434 1396 437 1416
rect 426 1393 437 1396
rect 442 1396 445 1606
rect 466 1593 469 1616
rect 466 1523 469 1536
rect 474 1533 485 1536
rect 490 1523 493 1616
rect 450 1413 453 1446
rect 498 1426 501 1696
rect 506 1543 509 1626
rect 514 1536 517 1736
rect 522 1723 525 1743
rect 538 1626 541 1763
rect 546 1753 549 1826
rect 554 1803 557 1936
rect 570 1883 573 1926
rect 570 1783 573 1806
rect 578 1776 581 1936
rect 642 1933 645 1946
rect 586 1813 589 1836
rect 570 1773 581 1776
rect 554 1733 557 1746
rect 534 1623 541 1626
rect 534 1556 537 1623
rect 534 1553 541 1556
rect 506 1533 517 1536
rect 506 1516 509 1533
rect 506 1513 517 1516
rect 498 1423 509 1426
rect 442 1393 449 1396
rect 402 1343 413 1346
rect 410 1296 413 1343
rect 426 1323 429 1393
rect 402 1293 413 1296
rect 378 1283 397 1286
rect 370 1213 373 1226
rect 378 1203 381 1236
rect 394 1216 397 1283
rect 402 1276 405 1293
rect 446 1286 449 1393
rect 458 1313 461 1326
rect 466 1303 469 1376
rect 442 1283 449 1286
rect 402 1273 413 1276
rect 402 1223 405 1273
rect 394 1213 405 1216
rect 322 1193 333 1196
rect 298 953 317 956
rect 298 926 301 953
rect 306 943 325 946
rect 306 933 309 943
rect 234 913 237 926
rect 266 903 269 926
rect 274 913 277 926
rect 298 923 309 926
rect 242 813 245 826
rect 298 816 301 836
rect 290 813 301 816
rect 186 713 189 736
rect 194 733 197 746
rect 210 713 213 726
rect 170 633 181 636
rect 122 623 133 626
rect 106 523 109 616
rect 130 576 133 623
rect 122 573 133 576
rect 74 503 85 506
rect 74 446 77 503
rect 66 443 77 446
rect 66 376 69 443
rect 82 383 85 406
rect 66 373 93 376
rect 90 306 93 373
rect 82 303 93 306
rect 82 133 85 303
rect 122 233 125 573
rect 162 523 165 616
rect 170 613 173 633
rect 170 596 173 606
rect 178 603 181 616
rect 186 596 189 616
rect 170 593 189 596
rect 130 413 133 426
rect 170 423 173 526
rect 186 523 189 556
rect 194 486 197 606
rect 202 553 205 656
rect 218 603 221 776
rect 226 683 229 726
rect 242 723 245 736
rect 250 723 253 796
rect 258 766 261 786
rect 290 766 293 813
rect 258 763 269 766
rect 290 763 301 766
rect 266 716 269 763
rect 290 733 293 746
rect 258 713 269 716
rect 234 596 237 706
rect 234 593 241 596
rect 202 543 221 546
rect 202 533 205 543
rect 210 493 213 536
rect 218 523 221 543
rect 194 483 213 486
rect 194 413 197 426
rect 138 313 141 326
rect 170 323 173 396
rect 202 333 205 406
rect 178 313 181 326
rect 114 123 117 216
rect 162 123 165 216
rect 170 213 173 226
rect 170 196 173 206
rect 178 203 181 306
rect 186 196 189 216
rect 202 213 205 236
rect 210 203 213 483
rect 226 423 229 586
rect 238 546 241 593
rect 234 543 241 546
rect 218 333 221 416
rect 226 393 229 406
rect 234 356 237 543
rect 242 513 245 526
rect 258 386 261 713
rect 290 706 293 726
rect 282 703 293 706
rect 298 706 301 763
rect 306 723 309 923
rect 314 903 317 936
rect 322 923 325 943
rect 330 833 333 1193
rect 346 1193 357 1196
rect 346 1116 349 1193
rect 362 1123 365 1196
rect 346 1113 357 1116
rect 338 913 341 1006
rect 346 903 349 936
rect 354 923 357 1113
rect 370 1023 389 1026
rect 370 1013 373 1023
rect 362 993 365 1006
rect 370 933 373 1006
rect 378 1003 381 1016
rect 386 996 389 1023
rect 402 1003 405 1213
rect 418 1123 421 1216
rect 434 1203 437 1216
rect 442 1026 445 1283
rect 474 1276 477 1396
rect 482 1323 485 1406
rect 490 1313 493 1336
rect 466 1273 477 1276
rect 458 1213 461 1236
rect 458 1196 461 1206
rect 466 1203 469 1273
rect 474 1196 477 1216
rect 498 1213 501 1326
rect 506 1323 509 1423
rect 514 1333 517 1513
rect 522 1413 525 1526
rect 530 1523 533 1536
rect 538 1516 541 1553
rect 546 1533 549 1616
rect 554 1596 557 1726
rect 570 1613 573 1773
rect 594 1713 597 1726
rect 602 1723 605 1816
rect 626 1813 629 1926
rect 654 1916 657 2023
rect 666 1993 669 2016
rect 666 1933 669 1946
rect 654 1913 661 1916
rect 642 1813 645 1836
rect 642 1793 645 1806
rect 650 1723 653 1806
rect 658 1706 661 1913
rect 674 1846 677 2166
rect 682 2096 685 2343
rect 690 2303 693 2466
rect 698 2413 701 2483
rect 710 2446 713 2503
rect 730 2463 733 2536
rect 706 2443 713 2446
rect 706 2403 709 2443
rect 714 2413 717 2426
rect 722 2353 725 2406
rect 722 2333 725 2346
rect 738 2296 741 2553
rect 746 2533 749 2693
rect 766 2636 769 2763
rect 766 2633 773 2636
rect 762 2536 765 2616
rect 754 2533 765 2536
rect 746 2503 749 2526
rect 754 2313 757 2533
rect 770 2503 773 2633
rect 778 2533 781 3093
rect 786 2996 789 3086
rect 794 3013 797 3136
rect 810 3133 813 3206
rect 826 3143 829 3196
rect 834 3143 845 3146
rect 826 3133 837 3136
rect 802 3106 805 3126
rect 802 3103 809 3106
rect 786 2993 793 2996
rect 790 2846 793 2993
rect 806 2986 809 3103
rect 802 2983 809 2986
rect 802 2963 805 2983
rect 818 2963 821 3126
rect 834 3056 837 3133
rect 834 3053 841 3056
rect 826 2946 829 3046
rect 818 2943 829 2946
rect 818 2886 821 2943
rect 838 2936 841 3053
rect 834 2933 841 2936
rect 834 2896 837 2933
rect 834 2893 841 2896
rect 818 2883 829 2886
rect 786 2843 793 2846
rect 786 2776 789 2843
rect 794 2793 797 2826
rect 786 2773 793 2776
rect 790 2616 793 2773
rect 786 2613 793 2616
rect 778 2513 781 2526
rect 786 2496 789 2613
rect 794 2553 797 2596
rect 782 2493 789 2496
rect 706 2213 709 2296
rect 730 2293 741 2296
rect 714 2163 717 2286
rect 730 2226 733 2293
rect 730 2223 741 2226
rect 698 2133 701 2146
rect 722 2113 725 2126
rect 730 2096 733 2206
rect 738 2153 741 2223
rect 682 2093 693 2096
rect 690 2046 693 2093
rect 682 2043 693 2046
rect 714 2093 733 2096
rect 682 2023 685 2043
rect 682 1943 685 2016
rect 714 2013 717 2093
rect 722 2013 733 2016
rect 714 1933 717 2006
rect 738 1933 741 2146
rect 746 2033 749 2306
rect 754 2203 757 2216
rect 770 2196 773 2426
rect 782 2346 785 2493
rect 794 2423 797 2536
rect 782 2343 789 2346
rect 766 2193 773 2196
rect 766 2116 769 2193
rect 778 2123 781 2326
rect 786 2276 789 2343
rect 794 2293 797 2406
rect 786 2273 793 2276
rect 790 2116 793 2273
rect 766 2113 773 2116
rect 746 2013 749 2026
rect 754 2013 757 2086
rect 770 2023 773 2113
rect 786 2113 793 2116
rect 762 1946 765 2006
rect 762 1943 769 1946
rect 722 1853 725 1926
rect 766 1896 769 1943
rect 778 1913 781 1926
rect 762 1893 769 1896
rect 650 1703 661 1706
rect 666 1843 677 1846
rect 554 1593 565 1596
rect 562 1546 565 1593
rect 594 1563 597 1606
rect 610 1593 613 1606
rect 554 1543 565 1546
rect 530 1403 533 1516
rect 538 1513 545 1516
rect 542 1436 545 1513
rect 554 1456 557 1543
rect 554 1453 565 1456
rect 538 1433 545 1436
rect 538 1336 541 1433
rect 546 1403 549 1416
rect 530 1333 541 1336
rect 530 1256 533 1333
rect 458 1193 477 1196
rect 482 1193 485 1206
rect 514 1203 517 1256
rect 530 1253 541 1256
rect 546 1253 549 1326
rect 538 1233 541 1253
rect 554 1243 557 1336
rect 562 1303 565 1453
rect 570 1346 573 1406
rect 570 1343 581 1346
rect 570 1313 573 1336
rect 578 1323 581 1343
rect 586 1316 589 1496
rect 594 1483 597 1536
rect 618 1523 621 1616
rect 626 1613 629 1646
rect 650 1596 653 1703
rect 666 1686 669 1843
rect 674 1776 677 1816
rect 690 1813 693 1826
rect 682 1796 685 1806
rect 682 1793 709 1796
rect 674 1773 681 1776
rect 662 1683 669 1686
rect 662 1616 665 1683
rect 678 1676 681 1773
rect 674 1673 681 1676
rect 690 1676 693 1776
rect 714 1773 717 1806
rect 690 1673 701 1676
rect 662 1613 669 1616
rect 650 1593 661 1596
rect 658 1573 661 1593
rect 650 1343 653 1486
rect 666 1443 669 1613
rect 674 1593 677 1673
rect 698 1616 701 1673
rect 682 1583 685 1606
rect 690 1603 693 1616
rect 698 1613 709 1616
rect 682 1513 685 1536
rect 698 1523 701 1606
rect 706 1603 709 1613
rect 706 1523 709 1596
rect 722 1533 725 1576
rect 730 1523 733 1876
rect 746 1813 749 1826
rect 754 1806 757 1816
rect 746 1803 757 1806
rect 762 1803 765 1893
rect 746 1723 749 1803
rect 770 1676 773 1746
rect 762 1673 773 1676
rect 762 1576 765 1673
rect 762 1573 773 1576
rect 746 1523 749 1556
rect 698 1413 701 1426
rect 746 1413 749 1426
rect 754 1413 757 1536
rect 770 1483 773 1573
rect 786 1536 789 2113
rect 802 2043 805 2876
rect 826 2863 829 2883
rect 838 2846 841 2893
rect 834 2843 841 2846
rect 810 2716 813 2806
rect 818 2793 821 2806
rect 826 2743 829 2816
rect 834 2783 837 2843
rect 842 2813 845 2826
rect 834 2733 837 2746
rect 850 2716 853 3213
rect 858 3193 861 3206
rect 866 2956 869 3486
rect 906 3483 917 3486
rect 914 3356 917 3483
rect 914 3353 933 3356
rect 890 3333 909 3336
rect 890 3316 893 3333
rect 886 3313 893 3316
rect 886 3236 889 3313
rect 886 3233 893 3236
rect 890 3213 893 3233
rect 882 3163 885 3206
rect 898 3203 901 3326
rect 914 3313 917 3326
rect 874 3123 877 3136
rect 882 3123 885 3146
rect 890 3106 893 3176
rect 882 3103 893 3106
rect 882 2966 885 3103
rect 898 3023 901 3136
rect 898 2993 901 3016
rect 882 2963 889 2966
rect 810 2713 821 2716
rect 818 2646 821 2713
rect 814 2643 821 2646
rect 842 2713 853 2716
rect 862 2953 869 2956
rect 842 2646 845 2713
rect 862 2646 865 2953
rect 874 2913 877 2946
rect 874 2656 877 2906
rect 886 2826 889 2963
rect 898 2933 901 2976
rect 906 2896 909 3216
rect 914 3203 917 3216
rect 922 3193 925 3326
rect 930 3176 933 3353
rect 938 3296 941 3493
rect 966 3476 969 3593
rect 978 3566 981 3626
rect 986 3616 989 3983
rect 1002 3953 1005 4206
rect 1010 4113 1013 4126
rect 1018 4076 1021 4136
rect 1026 4096 1029 4206
rect 1042 4156 1045 4213
rect 1058 4193 1061 4226
rect 1034 4153 1045 4156
rect 1034 4113 1037 4153
rect 1026 4093 1033 4096
rect 1010 4073 1021 4076
rect 994 3933 997 3946
rect 994 3893 997 3926
rect 1002 3913 1005 3926
rect 1010 3876 1013 4073
rect 1030 4036 1033 4093
rect 1030 4033 1037 4036
rect 1002 3873 1013 3876
rect 1002 3816 1005 3873
rect 998 3813 1005 3816
rect 998 3756 1001 3813
rect 994 3753 1001 3756
rect 994 3623 997 3753
rect 1002 3706 1005 3736
rect 1010 3723 1013 3806
rect 1002 3703 1009 3706
rect 1006 3626 1009 3703
rect 1002 3623 1009 3626
rect 986 3613 997 3616
rect 978 3563 989 3566
rect 962 3473 969 3476
rect 962 3356 965 3473
rect 986 3456 989 3563
rect 978 3453 989 3456
rect 978 3376 981 3453
rect 978 3373 985 3376
rect 962 3353 973 3356
rect 946 3316 949 3336
rect 946 3313 957 3316
rect 938 3293 945 3296
rect 942 3216 945 3293
rect 926 3173 933 3176
rect 938 3213 945 3216
rect 914 3133 917 3156
rect 914 3096 917 3126
rect 926 3116 929 3173
rect 926 3113 933 3116
rect 914 3093 925 3096
rect 914 2973 917 3016
rect 922 3003 925 3093
rect 930 3043 933 3113
rect 914 2913 917 2926
rect 922 2923 925 2996
rect 906 2893 917 2896
rect 886 2823 893 2826
rect 882 2793 885 2806
rect 874 2653 881 2656
rect 842 2643 853 2646
rect 862 2643 869 2646
rect 814 2526 817 2643
rect 850 2626 853 2643
rect 826 2613 829 2626
rect 850 2623 861 2626
rect 834 2613 853 2616
rect 834 2603 837 2613
rect 858 2593 861 2623
rect 826 2533 829 2556
rect 810 2523 817 2526
rect 810 2176 813 2523
rect 834 2513 837 2536
rect 818 2283 821 2506
rect 826 2413 829 2426
rect 810 2173 817 2176
rect 814 2126 817 2173
rect 826 2143 829 2346
rect 842 2343 845 2536
rect 858 2473 861 2546
rect 834 2313 837 2326
rect 850 2313 853 2366
rect 858 2343 861 2386
rect 866 2326 869 2643
rect 878 2546 881 2653
rect 862 2323 869 2326
rect 874 2543 881 2546
rect 814 2123 821 2126
rect 850 2123 853 2216
rect 862 2146 865 2323
rect 862 2143 869 2146
rect 818 2046 821 2123
rect 810 2043 821 2046
rect 802 2003 805 2036
rect 810 1986 813 2043
rect 806 1983 813 1986
rect 806 1926 809 1983
rect 818 1936 821 2016
rect 834 2013 837 2026
rect 842 1983 845 1996
rect 818 1933 829 1936
rect 806 1923 813 1926
rect 794 1733 797 1746
rect 810 1716 813 1923
rect 826 1893 829 1926
rect 834 1913 837 1926
rect 834 1813 837 1886
rect 842 1873 845 1926
rect 850 1813 853 2046
rect 858 1893 861 2126
rect 866 1876 869 2143
rect 874 1916 877 2543
rect 882 2413 885 2526
rect 882 2333 885 2346
rect 890 2256 893 2823
rect 898 2756 901 2886
rect 914 2776 917 2893
rect 930 2803 933 3006
rect 938 2906 941 3213
rect 954 3196 957 3313
rect 946 3193 957 3196
rect 946 3083 949 3193
rect 954 3076 957 3176
rect 970 3136 973 3353
rect 982 3186 985 3373
rect 994 3193 997 3613
rect 1002 3506 1005 3623
rect 1010 3523 1013 3606
rect 1018 3526 1021 4006
rect 1026 4003 1029 4026
rect 1034 3943 1037 4033
rect 1042 4013 1045 4136
rect 1050 4123 1053 4136
rect 1074 4133 1077 4316
rect 1082 4313 1093 4316
rect 1090 4266 1093 4313
rect 1082 4263 1093 4266
rect 1082 4186 1085 4263
rect 1090 4203 1093 4226
rect 1082 4183 1089 4186
rect 1050 4013 1053 4116
rect 1074 4103 1077 4116
rect 1086 4096 1089 4183
rect 1098 4123 1101 4246
rect 1130 4243 1133 4326
rect 1146 4316 1149 4336
rect 1154 4333 1157 4346
rect 1146 4313 1157 4316
rect 1154 4236 1157 4313
rect 1178 4283 1181 4416
rect 1234 4406 1237 4516
rect 1250 4486 1253 4526
rect 1266 4503 1269 4516
rect 1290 4513 1293 4526
rect 1314 4523 1317 4536
rect 1250 4483 1261 4486
rect 1258 4436 1261 4483
rect 1186 4403 1197 4406
rect 1226 4403 1237 4406
rect 1250 4433 1261 4436
rect 1202 4326 1205 4376
rect 1226 4346 1229 4403
rect 1226 4343 1237 4346
rect 1202 4323 1213 4326
rect 1106 4183 1109 4236
rect 1146 4233 1157 4236
rect 1114 4156 1117 4206
rect 1130 4196 1133 4216
rect 1138 4203 1141 4226
rect 1146 4213 1149 4233
rect 1146 4196 1149 4206
rect 1130 4193 1149 4196
rect 1110 4153 1117 4156
rect 1082 4093 1089 4096
rect 1026 3893 1029 3936
rect 1034 3923 1037 3936
rect 1066 3916 1069 3956
rect 1074 3933 1077 4016
rect 1082 4013 1085 4093
rect 1110 4076 1113 4153
rect 1122 4083 1125 4146
rect 1138 4143 1165 4146
rect 1110 4073 1117 4076
rect 1090 4013 1093 4036
rect 1082 3993 1085 4006
rect 1098 3963 1101 4016
rect 1058 3873 1061 3916
rect 1066 3913 1073 3916
rect 1026 3823 1029 3856
rect 1026 3743 1029 3766
rect 1042 3653 1045 3846
rect 1070 3796 1073 3913
rect 1066 3793 1073 3796
rect 1066 3746 1069 3793
rect 1058 3743 1069 3746
rect 1058 3636 1061 3743
rect 1074 3716 1077 3736
rect 1070 3713 1077 3716
rect 1070 3656 1073 3713
rect 1070 3653 1077 3656
rect 1026 3613 1029 3636
rect 1050 3633 1061 3636
rect 1042 3573 1045 3606
rect 1026 3543 1029 3556
rect 1018 3523 1029 3526
rect 1002 3503 1013 3506
rect 1010 3446 1013 3503
rect 1002 3443 1013 3446
rect 1002 3376 1005 3443
rect 1026 3426 1029 3523
rect 1018 3423 1029 3426
rect 1010 3393 1013 3416
rect 1002 3373 1009 3376
rect 1006 3226 1009 3373
rect 1002 3223 1009 3226
rect 1002 3193 1005 3223
rect 1018 3213 1021 3423
rect 1050 3416 1053 3633
rect 1066 3613 1069 3626
rect 1058 3583 1061 3606
rect 1074 3553 1077 3653
rect 1066 3483 1069 3536
rect 1074 3523 1077 3546
rect 1082 3466 1085 3946
rect 1106 3856 1109 3956
rect 1114 3953 1117 4073
rect 1130 4003 1133 4016
rect 1138 3936 1141 4143
rect 1154 4126 1157 4136
rect 1162 4133 1165 4143
rect 1146 4113 1149 4126
rect 1154 4123 1173 4126
rect 1186 4123 1189 4226
rect 1194 4223 1197 4316
rect 1194 4193 1197 4206
rect 1210 4176 1213 4323
rect 1234 4223 1237 4343
rect 1250 4223 1253 4433
rect 1306 4423 1309 4516
rect 1330 4413 1333 4526
rect 1346 4523 1349 4546
rect 1354 4513 1357 4536
rect 1378 4533 1381 4583
rect 1386 4523 1389 4536
rect 1394 4523 1397 4546
rect 1402 4533 1405 4606
rect 1418 4593 1421 4606
rect 1466 4603 1469 4616
rect 1426 4503 1429 4536
rect 1434 4523 1437 4536
rect 1258 4303 1261 4336
rect 1274 4333 1277 4346
rect 1298 4333 1301 4406
rect 1306 4363 1309 4406
rect 1354 4403 1357 4426
rect 1362 4333 1365 4416
rect 1418 4403 1421 4416
rect 1322 4313 1325 4326
rect 1362 4306 1365 4326
rect 1370 4323 1373 4336
rect 1354 4303 1365 4306
rect 1354 4246 1357 4303
rect 1202 4173 1213 4176
rect 1146 3996 1149 4016
rect 1154 4003 1157 4036
rect 1162 4016 1165 4026
rect 1162 4013 1173 4016
rect 1162 3996 1165 4006
rect 1146 3993 1165 3996
rect 1130 3933 1141 3936
rect 1130 3866 1133 3933
rect 1130 3863 1141 3866
rect 1106 3853 1113 3856
rect 1090 3813 1093 3826
rect 1110 3776 1113 3853
rect 1106 3773 1113 3776
rect 1090 3723 1093 3746
rect 1090 3603 1093 3626
rect 1098 3493 1101 3656
rect 1106 3633 1109 3773
rect 1122 3733 1125 3846
rect 1130 3813 1133 3826
rect 1138 3796 1141 3863
rect 1146 3813 1149 3976
rect 1170 3973 1173 4013
rect 1134 3793 1141 3796
rect 1146 3796 1149 3806
rect 1154 3803 1157 3846
rect 1162 3796 1165 3816
rect 1146 3793 1165 3796
rect 1134 3726 1137 3793
rect 1146 3733 1149 3746
rect 1134 3723 1141 3726
rect 1138 3626 1141 3723
rect 1130 3616 1133 3626
rect 1138 3623 1149 3626
rect 1114 3596 1117 3616
rect 1122 3603 1125 3616
rect 1130 3613 1141 3616
rect 1130 3603 1141 3606
rect 1114 3593 1125 3596
rect 1122 3523 1125 3593
rect 1130 3486 1133 3556
rect 1074 3463 1085 3466
rect 1050 3413 1061 3416
rect 1042 3323 1045 3406
rect 1058 3316 1061 3413
rect 1050 3313 1061 3316
rect 1074 3316 1077 3463
rect 1090 3323 1093 3476
rect 1074 3313 1085 3316
rect 1026 3286 1029 3306
rect 1026 3283 1037 3286
rect 1034 3236 1037 3283
rect 1026 3233 1037 3236
rect 1026 3206 1029 3233
rect 1034 3213 1045 3216
rect 982 3183 989 3186
rect 962 3133 973 3136
rect 978 3133 981 3146
rect 962 3083 965 3133
rect 970 3123 981 3126
rect 986 3123 989 3183
rect 1010 3143 1013 3206
rect 1026 3203 1037 3206
rect 978 3096 981 3116
rect 986 3096 989 3116
rect 978 3093 989 3096
rect 946 3073 957 3076
rect 946 2993 949 3073
rect 946 2943 949 2956
rect 946 2913 949 2936
rect 938 2903 949 2906
rect 938 2793 941 2816
rect 914 2773 925 2776
rect 898 2753 909 2756
rect 906 2676 909 2753
rect 898 2673 909 2676
rect 898 2533 901 2673
rect 922 2656 925 2773
rect 906 2653 925 2656
rect 906 2483 909 2653
rect 922 2613 925 2636
rect 946 2613 949 2903
rect 954 2893 957 2916
rect 962 2886 965 3026
rect 970 3023 973 3066
rect 994 3046 997 3136
rect 1002 3103 1005 3126
rect 986 3043 997 3046
rect 986 2903 989 3043
rect 994 3013 997 3036
rect 1002 2886 1005 3056
rect 1010 2966 1013 3136
rect 1018 3133 1021 3196
rect 1018 3106 1021 3126
rect 1018 3103 1029 3106
rect 1018 3013 1021 3086
rect 1026 3053 1029 3103
rect 1026 2983 1029 2996
rect 1010 2963 1021 2966
rect 1018 2896 1021 2963
rect 962 2883 973 2886
rect 970 2836 973 2883
rect 962 2833 973 2836
rect 994 2883 1005 2886
rect 1010 2893 1021 2896
rect 962 2813 965 2833
rect 994 2816 997 2883
rect 1010 2873 1013 2893
rect 1034 2883 1037 3203
rect 1050 3153 1053 3313
rect 1058 3123 1061 3216
rect 1066 3213 1069 3226
rect 1066 3176 1069 3196
rect 1074 3183 1077 3206
rect 1066 3173 1077 3176
rect 1066 3106 1069 3156
rect 1062 3103 1069 3106
rect 994 2813 1005 2816
rect 1010 2813 1013 2826
rect 1034 2813 1037 2846
rect 962 2723 965 2806
rect 978 2656 981 2796
rect 978 2653 989 2656
rect 914 2586 917 2606
rect 914 2583 921 2586
rect 918 2476 921 2583
rect 914 2473 921 2476
rect 890 2253 901 2256
rect 882 1933 885 2176
rect 898 2146 901 2253
rect 914 2226 917 2473
rect 922 2323 925 2346
rect 930 2243 933 2596
rect 946 2546 949 2606
rect 954 2593 957 2606
rect 942 2543 949 2546
rect 942 2406 945 2543
rect 954 2413 957 2536
rect 962 2523 965 2536
rect 970 2423 973 2556
rect 978 2523 981 2653
rect 1002 2616 1005 2813
rect 1026 2746 1029 2806
rect 1042 2793 1045 3056
rect 1062 3046 1065 3103
rect 1074 3053 1077 3173
rect 1082 3076 1085 3313
rect 1090 3193 1093 3216
rect 1082 3073 1089 3076
rect 1050 3026 1053 3046
rect 1062 3043 1069 3046
rect 1050 3023 1057 3026
rect 1054 2856 1057 3023
rect 1050 2853 1057 2856
rect 1050 2813 1053 2853
rect 1058 2813 1061 2836
rect 1018 2743 1029 2746
rect 1018 2696 1021 2743
rect 1018 2693 1029 2696
rect 994 2613 1005 2616
rect 994 2556 997 2613
rect 994 2553 1005 2556
rect 986 2533 997 2536
rect 1002 2496 1005 2553
rect 1010 2533 1013 2606
rect 1018 2503 1021 2676
rect 1026 2586 1029 2693
rect 1034 2603 1037 2736
rect 1042 2693 1045 2726
rect 1050 2716 1053 2736
rect 1066 2723 1069 3043
rect 1074 2956 1077 3006
rect 1086 2976 1089 3073
rect 1098 2993 1101 3336
rect 1106 3323 1109 3486
rect 1122 3483 1133 3486
rect 1122 3256 1125 3483
rect 1138 3356 1141 3596
rect 1134 3353 1141 3356
rect 1134 3276 1137 3353
rect 1134 3273 1141 3276
rect 1122 3253 1133 3256
rect 1130 3236 1133 3253
rect 1106 3203 1109 3216
rect 1114 3203 1117 3236
rect 1122 3233 1133 3236
rect 1106 3126 1109 3146
rect 1106 3123 1113 3126
rect 1110 3026 1113 3123
rect 1106 3023 1113 3026
rect 1106 2976 1109 3023
rect 1086 2973 1093 2976
rect 1074 2953 1081 2956
rect 1078 2856 1081 2953
rect 1074 2853 1081 2856
rect 1050 2713 1057 2716
rect 1042 2603 1045 2686
rect 1054 2636 1057 2713
rect 1074 2683 1077 2853
rect 1090 2836 1093 2973
rect 1082 2833 1093 2836
rect 1102 2973 1109 2976
rect 1082 2676 1085 2833
rect 1102 2816 1105 2973
rect 1098 2813 1105 2816
rect 1078 2673 1085 2676
rect 1050 2633 1057 2636
rect 1026 2583 1037 2586
rect 1034 2516 1037 2583
rect 1050 2546 1053 2633
rect 1058 2593 1061 2616
rect 1066 2613 1069 2656
rect 1030 2513 1037 2516
rect 1046 2543 1053 2546
rect 1002 2493 1021 2496
rect 994 2413 997 2436
rect 1010 2413 1013 2486
rect 942 2403 949 2406
rect 890 2143 901 2146
rect 910 2223 917 2226
rect 890 2096 893 2143
rect 898 2113 901 2126
rect 890 2093 901 2096
rect 898 2026 901 2093
rect 890 2023 901 2026
rect 910 2026 913 2223
rect 910 2023 917 2026
rect 874 1913 881 1916
rect 862 1873 869 1876
rect 818 1786 821 1806
rect 818 1783 829 1786
rect 826 1726 829 1783
rect 802 1713 813 1716
rect 818 1723 829 1726
rect 802 1636 805 1713
rect 802 1633 813 1636
rect 802 1603 805 1616
rect 778 1533 789 1536
rect 794 1533 797 1556
rect 610 1333 621 1336
rect 578 1313 589 1316
rect 578 1226 581 1313
rect 602 1256 605 1306
rect 618 1273 621 1326
rect 658 1303 661 1336
rect 674 1333 677 1346
rect 722 1313 725 1326
rect 602 1253 609 1256
rect 522 1213 525 1226
rect 562 1213 565 1226
rect 578 1223 585 1226
rect 482 1133 485 1166
rect 538 1163 541 1206
rect 570 1156 573 1216
rect 554 1153 573 1156
rect 530 1123 533 1136
rect 554 1026 557 1153
rect 562 1123 565 1146
rect 570 1133 573 1153
rect 582 1146 585 1223
rect 606 1156 609 1253
rect 618 1213 621 1246
rect 626 1193 629 1206
rect 602 1153 609 1156
rect 578 1143 585 1146
rect 570 1053 573 1126
rect 578 1103 581 1143
rect 594 1133 597 1146
rect 586 1113 589 1126
rect 602 1106 605 1153
rect 610 1123 613 1136
rect 634 1113 637 1136
rect 598 1103 605 1106
rect 598 1036 601 1103
rect 598 1033 605 1036
rect 442 1023 453 1026
rect 554 1023 561 1026
rect 378 993 389 996
rect 378 906 381 993
rect 386 923 389 936
rect 394 906 397 926
rect 370 903 381 906
rect 386 903 397 906
rect 314 733 317 816
rect 338 743 341 846
rect 370 806 373 903
rect 386 813 389 903
rect 434 843 437 936
rect 442 923 445 1016
rect 450 826 453 1023
rect 458 943 477 946
rect 458 933 461 943
rect 458 913 461 926
rect 466 923 469 936
rect 474 923 477 943
rect 482 933 485 1016
rect 514 1003 517 1016
rect 514 913 517 926
rect 442 823 453 826
rect 370 803 381 806
rect 330 733 341 736
rect 346 733 349 756
rect 322 713 325 726
rect 298 703 305 706
rect 282 656 285 703
rect 282 653 293 656
rect 274 403 277 426
rect 282 413 285 526
rect 290 413 293 653
rect 302 636 305 703
rect 338 693 341 726
rect 354 703 357 726
rect 298 633 305 636
rect 298 586 301 633
rect 306 603 309 616
rect 298 583 305 586
rect 302 516 305 583
rect 298 513 305 516
rect 322 523 341 526
rect 346 523 349 606
rect 354 583 357 606
rect 362 593 365 616
rect 370 613 373 716
rect 378 693 381 803
rect 442 776 445 823
rect 458 813 461 826
rect 474 813 477 846
rect 466 783 469 806
rect 482 803 485 836
rect 530 813 533 846
rect 386 676 389 746
rect 394 723 397 736
rect 410 733 413 776
rect 442 773 453 776
rect 418 733 421 766
rect 450 743 453 773
rect 490 763 493 806
rect 538 773 541 926
rect 546 923 549 1016
rect 558 946 561 1023
rect 554 943 561 946
rect 570 943 589 946
rect 554 923 557 943
rect 570 933 573 943
rect 562 816 565 916
rect 570 893 573 926
rect 578 923 581 936
rect 586 923 589 943
rect 546 753 549 816
rect 554 813 565 816
rect 594 813 597 1016
rect 602 913 605 1033
rect 610 973 613 1106
rect 642 1096 645 1146
rect 650 1106 653 1226
rect 666 1216 669 1276
rect 746 1256 749 1346
rect 738 1253 749 1256
rect 666 1213 677 1216
rect 682 1213 685 1226
rect 658 1183 661 1206
rect 658 1123 661 1166
rect 682 1163 685 1206
rect 698 1203 701 1246
rect 722 1213 733 1216
rect 690 1106 693 1156
rect 714 1123 717 1206
rect 722 1193 725 1206
rect 650 1103 661 1106
rect 690 1103 701 1106
rect 634 1093 645 1096
rect 634 1026 637 1093
rect 658 1036 661 1103
rect 650 1033 661 1036
rect 634 1023 645 1026
rect 626 983 629 1006
rect 642 1003 645 1023
rect 650 1013 653 1033
rect 682 1003 685 1086
rect 698 1036 701 1103
rect 690 1033 701 1036
rect 642 956 645 976
rect 690 973 693 1033
rect 634 953 645 956
rect 634 906 637 953
rect 666 933 669 956
rect 738 953 741 1253
rect 746 1203 749 1216
rect 754 1203 757 1356
rect 762 1313 765 1326
rect 762 1123 765 1306
rect 778 1173 781 1533
rect 786 1513 789 1526
rect 802 1523 805 1566
rect 794 1306 797 1416
rect 802 1403 805 1426
rect 802 1313 805 1336
rect 810 1316 813 1633
rect 818 1613 821 1723
rect 834 1613 837 1706
rect 850 1676 853 1806
rect 862 1776 865 1873
rect 878 1866 881 1913
rect 890 1883 893 2023
rect 898 1923 901 2006
rect 906 1993 909 2006
rect 906 1906 909 1946
rect 902 1903 909 1906
rect 874 1863 881 1866
rect 862 1773 869 1776
rect 858 1743 861 1756
rect 866 1743 869 1773
rect 874 1726 877 1863
rect 902 1826 905 1903
rect 902 1823 909 1826
rect 846 1673 853 1676
rect 870 1723 877 1726
rect 846 1616 849 1673
rect 846 1613 853 1616
rect 818 1533 821 1546
rect 818 1506 821 1526
rect 834 1523 837 1606
rect 842 1583 845 1596
rect 850 1533 853 1613
rect 858 1526 861 1666
rect 850 1523 861 1526
rect 818 1503 829 1506
rect 826 1446 829 1503
rect 818 1443 829 1446
rect 818 1423 821 1443
rect 818 1403 821 1416
rect 842 1413 845 1426
rect 818 1333 821 1356
rect 842 1326 845 1366
rect 850 1333 853 1523
rect 858 1413 861 1446
rect 870 1416 873 1723
rect 870 1413 877 1416
rect 858 1393 869 1396
rect 858 1333 861 1346
rect 810 1313 821 1316
rect 834 1313 837 1326
rect 842 1323 853 1326
rect 794 1303 805 1306
rect 794 1203 797 1226
rect 802 1213 805 1303
rect 818 1246 821 1313
rect 810 1243 821 1246
rect 802 1163 805 1206
rect 810 1063 813 1243
rect 818 1213 821 1226
rect 834 1213 837 1246
rect 834 1163 837 1206
rect 842 1203 845 1216
rect 818 1123 821 1136
rect 746 1013 757 1016
rect 802 1013 805 1026
rect 842 1013 845 1026
rect 826 986 829 1006
rect 778 983 789 986
rect 754 933 757 946
rect 634 903 645 906
rect 402 713 405 726
rect 426 713 429 736
rect 482 733 485 746
rect 382 673 389 676
rect 382 616 385 673
rect 378 613 385 616
rect 394 613 397 696
rect 378 586 381 613
rect 386 603 397 606
rect 402 603 405 616
rect 450 613 453 726
rect 506 613 509 726
rect 530 713 533 726
rect 546 626 549 646
rect 554 633 557 813
rect 562 723 565 806
rect 570 713 573 726
rect 514 613 517 626
rect 546 623 557 626
rect 362 583 381 586
rect 298 493 301 513
rect 322 476 325 523
rect 314 473 325 476
rect 314 426 317 473
rect 314 423 325 426
rect 322 403 325 423
rect 330 413 333 426
rect 338 403 341 496
rect 230 353 237 356
rect 250 383 261 386
rect 230 306 233 353
rect 250 333 253 383
rect 298 313 301 326
rect 330 323 333 346
rect 338 313 341 326
rect 230 303 237 306
rect 170 193 189 196
rect 178 133 181 146
rect 218 123 221 216
rect 226 213 229 246
rect 234 223 237 303
rect 234 196 237 206
rect 242 203 245 216
rect 250 196 253 216
rect 266 213 269 226
rect 234 193 253 196
rect 258 123 261 206
rect 298 203 301 226
rect 306 176 309 216
rect 314 213 317 246
rect 322 203 325 216
rect 330 213 333 226
rect 354 213 357 226
rect 306 173 325 176
rect 298 133 301 146
rect 322 123 325 173
rect 362 143 365 583
rect 386 543 405 546
rect 378 523 381 536
rect 386 533 389 543
rect 394 493 397 536
rect 402 523 405 543
rect 410 533 413 596
rect 426 536 429 606
rect 514 593 517 606
rect 426 533 437 536
rect 442 533 445 546
rect 450 543 469 546
rect 386 413 389 436
rect 370 323 373 336
rect 378 296 381 406
rect 394 403 397 476
rect 418 426 421 526
rect 426 436 429 526
rect 434 456 437 533
rect 450 523 453 543
rect 458 473 461 536
rect 466 533 469 543
rect 474 503 477 536
rect 434 453 461 456
rect 426 433 437 436
rect 418 423 429 426
rect 402 396 405 416
rect 410 403 413 416
rect 418 396 421 406
rect 402 393 421 396
rect 426 386 429 423
rect 434 413 437 433
rect 442 393 445 416
rect 418 383 429 386
rect 386 343 405 346
rect 386 333 389 343
rect 386 313 389 326
rect 394 296 397 336
rect 402 323 405 343
rect 410 333 413 346
rect 378 293 397 296
rect 370 213 373 266
rect 370 196 373 206
rect 378 203 381 293
rect 386 196 389 216
rect 394 203 397 216
rect 402 213 405 226
rect 418 223 421 383
rect 458 366 461 453
rect 498 413 501 526
rect 514 523 517 536
rect 530 523 533 616
rect 546 573 549 606
rect 554 583 557 623
rect 578 606 581 776
rect 586 733 589 756
rect 594 723 597 806
rect 610 756 613 836
rect 634 813 637 826
rect 618 803 629 806
rect 634 783 637 806
rect 602 753 613 756
rect 450 363 461 366
rect 450 333 453 363
rect 474 323 477 396
rect 530 323 533 416
rect 538 413 541 546
rect 562 543 565 606
rect 570 603 589 606
rect 570 526 573 596
rect 578 533 581 566
rect 570 523 581 526
rect 586 523 589 586
rect 594 553 597 636
rect 602 593 605 753
rect 642 713 645 903
rect 674 813 677 826
rect 674 793 677 806
rect 610 613 613 656
rect 546 343 549 406
rect 402 196 405 206
rect 370 193 381 196
rect 386 193 405 196
rect 378 123 381 193
rect 410 133 413 146
rect 434 123 437 216
rect 458 203 461 226
rect 474 196 477 216
rect 482 203 485 216
rect 490 213 493 316
rect 538 306 541 336
rect 534 303 541 306
rect 506 213 509 226
rect 522 213 525 236
rect 534 226 537 303
rect 530 223 537 226
rect 530 213 533 223
rect 546 216 549 336
rect 554 333 557 356
rect 562 333 565 516
rect 578 416 581 523
rect 594 423 597 536
rect 602 503 605 526
rect 578 413 597 416
rect 610 413 613 606
rect 626 593 629 616
rect 634 603 637 616
rect 642 613 645 636
rect 658 606 661 746
rect 682 693 685 896
rect 698 813 701 866
rect 714 813 717 926
rect 778 856 781 926
rect 786 923 789 983
rect 794 933 797 986
rect 826 983 837 986
rect 778 853 789 856
rect 690 773 693 806
rect 714 793 717 806
rect 738 803 741 826
rect 746 803 749 816
rect 754 736 757 816
rect 762 783 765 806
rect 770 746 773 836
rect 778 753 781 806
rect 786 793 789 853
rect 802 833 805 976
rect 834 953 837 983
rect 850 973 853 1316
rect 858 1213 861 1236
rect 866 1163 869 1336
rect 866 1123 869 1136
rect 818 933 821 946
rect 818 903 821 926
rect 826 923 829 936
rect 794 776 797 816
rect 810 813 813 826
rect 794 773 805 776
rect 770 743 781 746
rect 746 733 773 736
rect 618 523 621 586
rect 642 583 645 606
rect 650 603 661 606
rect 626 526 629 556
rect 634 533 637 546
rect 626 523 637 526
rect 650 523 653 603
rect 682 523 685 616
rect 690 613 693 726
rect 706 613 709 716
rect 738 706 741 726
rect 730 703 741 706
rect 730 636 733 703
rect 746 696 749 733
rect 754 713 757 726
rect 746 693 757 696
rect 754 646 757 693
rect 746 643 757 646
rect 730 633 741 636
rect 690 593 693 606
rect 730 556 733 606
rect 738 603 741 633
rect 730 553 741 556
rect 634 493 637 523
rect 618 413 621 436
rect 674 416 677 496
rect 562 256 565 326
rect 570 303 573 336
rect 578 313 581 413
rect 586 383 589 406
rect 594 403 605 406
rect 538 213 549 216
rect 554 253 565 256
rect 554 213 557 253
rect 570 213 573 266
rect 594 213 597 326
rect 610 213 613 236
rect 474 193 493 196
rect 490 123 493 193
rect 498 163 501 206
rect 514 173 517 206
rect 522 193 525 206
rect 546 193 549 206
rect 530 133 533 146
rect 554 123 557 206
rect 562 183 565 206
rect 570 163 573 206
rect 610 123 613 176
rect 618 123 621 246
rect 642 193 645 206
rect 650 163 653 406
rect 658 396 661 416
rect 666 403 669 416
rect 674 413 685 416
rect 674 396 677 406
rect 658 393 677 396
rect 682 336 685 413
rect 674 333 685 336
rect 658 196 661 216
rect 666 203 669 216
rect 674 213 677 333
rect 682 313 685 326
rect 698 236 701 526
rect 730 523 733 546
rect 738 513 741 553
rect 746 533 749 643
rect 770 593 773 606
rect 706 413 709 426
rect 746 413 749 426
rect 754 413 757 536
rect 770 533 773 546
rect 778 513 781 743
rect 794 733 797 746
rect 802 696 805 773
rect 818 746 821 806
rect 826 763 829 846
rect 834 803 837 936
rect 850 933 853 946
rect 866 926 869 1096
rect 842 906 845 926
rect 858 923 869 926
rect 842 903 849 906
rect 846 836 849 903
rect 842 833 849 836
rect 842 813 845 833
rect 810 743 821 746
rect 810 733 813 743
rect 794 693 805 696
rect 810 693 813 726
rect 818 703 821 743
rect 834 733 837 756
rect 826 723 837 726
rect 842 713 845 726
rect 850 723 853 736
rect 794 606 797 693
rect 810 613 813 656
rect 794 603 805 606
rect 818 603 821 616
rect 802 423 805 603
rect 834 536 837 706
rect 842 596 845 616
rect 850 603 853 616
rect 858 613 861 923
rect 874 906 877 1413
rect 882 1303 885 1816
rect 898 1783 901 1806
rect 890 1746 893 1766
rect 890 1743 897 1746
rect 894 1566 897 1743
rect 890 1563 897 1566
rect 882 1093 885 1216
rect 882 1003 885 1026
rect 890 996 893 1563
rect 898 1486 901 1546
rect 906 1503 909 1823
rect 898 1483 905 1486
rect 902 1416 905 1483
rect 898 1413 905 1416
rect 898 1313 901 1413
rect 914 1403 917 2023
rect 922 1646 925 2216
rect 930 2176 933 2236
rect 938 2193 941 2216
rect 930 2173 937 2176
rect 934 1986 937 2173
rect 930 1983 937 1986
rect 930 1943 933 1983
rect 930 1906 933 1936
rect 938 1923 941 1966
rect 930 1903 937 1906
rect 934 1776 937 1903
rect 930 1773 937 1776
rect 930 1733 933 1773
rect 938 1673 941 1756
rect 946 1666 949 2403
rect 954 2116 957 2246
rect 962 2233 965 2396
rect 986 2346 989 2406
rect 1010 2393 1013 2406
rect 978 2343 989 2346
rect 978 2236 981 2343
rect 978 2233 989 2236
rect 962 2153 965 2206
rect 962 2133 965 2146
rect 954 2113 961 2116
rect 958 1956 961 2113
rect 970 2043 973 2206
rect 978 2143 981 2216
rect 954 1953 961 1956
rect 954 1923 957 1953
rect 962 1906 965 1936
rect 958 1903 965 1906
rect 958 1746 961 1903
rect 958 1743 965 1746
rect 954 1703 957 1726
rect 938 1663 949 1666
rect 922 1643 929 1646
rect 926 1586 929 1643
rect 922 1583 929 1586
rect 922 1413 925 1583
rect 938 1566 941 1663
rect 962 1603 965 1743
rect 970 1723 973 2036
rect 978 1943 981 2126
rect 986 2006 989 2233
rect 994 2213 997 2336
rect 1002 2293 1005 2326
rect 1018 2323 1021 2493
rect 1030 2416 1033 2513
rect 1046 2496 1049 2543
rect 1058 2513 1061 2536
rect 1066 2496 1069 2606
rect 1078 2546 1081 2673
rect 1090 2553 1093 2806
rect 1098 2766 1101 2813
rect 1106 2783 1109 2806
rect 1098 2763 1105 2766
rect 1102 2636 1105 2763
rect 1098 2633 1105 2636
rect 1098 2613 1101 2633
rect 1098 2593 1101 2606
rect 1106 2603 1109 2616
rect 1078 2543 1101 2546
rect 1026 2413 1033 2416
rect 1042 2493 1049 2496
rect 1062 2493 1069 2496
rect 1026 2306 1029 2413
rect 1042 2406 1045 2493
rect 1042 2403 1053 2406
rect 1018 2303 1029 2306
rect 1018 2236 1021 2303
rect 1018 2233 1029 2236
rect 994 2193 997 2206
rect 994 2023 997 2126
rect 986 2003 993 2006
rect 978 1813 981 1936
rect 990 1896 993 2003
rect 1002 1933 1005 2206
rect 1010 2183 1013 2196
rect 1018 2123 1021 2216
rect 1026 2106 1029 2233
rect 1022 2103 1029 2106
rect 1010 1916 1013 2076
rect 1022 2026 1025 2103
rect 1034 2073 1037 2396
rect 1050 2356 1053 2403
rect 1042 2353 1053 2356
rect 1022 2023 1029 2026
rect 986 1893 993 1896
rect 1006 1913 1013 1916
rect 978 1743 981 1806
rect 986 1753 989 1893
rect 994 1813 997 1876
rect 1006 1786 1009 1913
rect 1006 1783 1013 1786
rect 1010 1763 1013 1783
rect 978 1706 981 1736
rect 974 1703 981 1706
rect 954 1573 957 1596
rect 930 1563 941 1566
rect 906 1323 909 1346
rect 930 1333 933 1563
rect 974 1546 977 1703
rect 986 1683 989 1726
rect 994 1706 997 1736
rect 1002 1733 1005 1746
rect 1010 1733 1013 1746
rect 1018 1723 1021 2006
rect 1026 1996 1029 2023
rect 1034 2013 1037 2026
rect 1026 1993 1033 1996
rect 1030 1836 1033 1993
rect 1026 1833 1033 1836
rect 1026 1706 1029 1833
rect 994 1703 1005 1706
rect 946 1533 949 1546
rect 970 1543 977 1546
rect 938 1486 941 1506
rect 970 1486 973 1543
rect 938 1483 945 1486
rect 942 1376 945 1483
rect 966 1483 973 1486
rect 954 1393 957 1436
rect 942 1373 949 1376
rect 898 1133 901 1216
rect 914 1213 917 1296
rect 906 1166 909 1206
rect 922 1183 925 1196
rect 906 1163 917 1166
rect 914 1146 917 1163
rect 906 1083 909 1146
rect 914 1143 921 1146
rect 918 1076 921 1143
rect 930 1126 933 1306
rect 946 1216 949 1373
rect 966 1346 969 1483
rect 966 1343 973 1346
rect 962 1313 965 1326
rect 970 1296 973 1343
rect 978 1333 981 1536
rect 986 1356 989 1676
rect 1002 1636 1005 1703
rect 998 1633 1005 1636
rect 1018 1703 1029 1706
rect 1018 1636 1021 1703
rect 1018 1633 1029 1636
rect 998 1576 1001 1633
rect 1010 1613 1021 1616
rect 994 1573 1001 1576
rect 994 1533 997 1573
rect 1026 1536 1029 1633
rect 1034 1603 1037 1816
rect 1010 1533 1029 1536
rect 994 1513 997 1526
rect 1010 1426 1013 1533
rect 1018 1523 1029 1526
rect 1034 1513 1037 1526
rect 1010 1423 1017 1426
rect 994 1403 997 1416
rect 1002 1373 1005 1416
rect 986 1353 997 1356
rect 962 1293 973 1296
rect 962 1226 965 1293
rect 962 1223 973 1226
rect 938 1213 949 1216
rect 938 1133 941 1213
rect 970 1203 973 1223
rect 962 1193 973 1196
rect 946 1126 949 1146
rect 930 1123 941 1126
rect 946 1123 957 1126
rect 914 1073 921 1076
rect 898 1003 901 1016
rect 906 1013 909 1026
rect 890 993 901 996
rect 870 903 877 906
rect 870 846 873 903
rect 870 843 877 846
rect 866 813 869 826
rect 874 693 877 843
rect 882 813 885 936
rect 898 856 901 993
rect 914 923 917 1073
rect 922 1013 925 1056
rect 922 993 933 996
rect 938 986 941 1123
rect 954 1026 957 1123
rect 946 1023 957 1026
rect 946 1003 949 1023
rect 930 983 941 986
rect 930 966 933 983
rect 926 963 933 966
rect 926 906 929 963
rect 926 903 933 906
rect 894 853 901 856
rect 894 776 897 853
rect 914 813 917 826
rect 894 773 901 776
rect 866 613 869 626
rect 882 613 893 616
rect 858 596 861 606
rect 842 593 861 596
rect 810 516 813 536
rect 834 533 853 536
rect 858 533 861 556
rect 810 513 821 516
rect 794 413 805 416
rect 818 406 821 513
rect 722 393 725 406
rect 810 403 821 406
rect 842 403 845 526
rect 850 523 853 533
rect 858 433 861 526
rect 866 523 869 536
rect 722 313 725 326
rect 690 233 701 236
rect 674 196 677 206
rect 658 193 677 196
rect 642 133 645 146
rect 682 123 685 216
rect 690 143 693 233
rect 698 213 701 226
rect 706 203 709 216
rect 714 203 725 206
rect 730 203 733 276
rect 738 263 741 316
rect 738 236 741 256
rect 738 233 749 236
rect 738 213 741 233
rect 754 213 757 226
rect 722 123 725 203
rect 746 123 749 206
rect 754 193 757 206
rect 778 203 781 326
rect 810 323 813 403
rect 810 203 813 216
rect 818 213 821 236
rect 826 203 829 256
rect 834 213 837 226
rect 834 183 837 206
rect 850 203 853 326
rect 858 323 861 416
rect 882 413 885 426
rect 890 306 893 586
rect 898 553 901 773
rect 930 766 933 903
rect 946 886 949 976
rect 946 883 965 886
rect 926 763 933 766
rect 906 713 909 726
rect 914 723 917 756
rect 926 686 929 763
rect 946 713 949 726
rect 926 683 933 686
rect 914 613 917 626
rect 930 596 933 683
rect 930 593 949 596
rect 914 543 941 546
rect 914 533 917 543
rect 906 313 909 326
rect 914 316 917 526
rect 922 513 925 526
rect 930 396 933 416
rect 938 403 941 536
rect 946 533 949 593
rect 962 583 965 883
rect 978 803 981 1316
rect 994 1236 997 1353
rect 1014 1346 1017 1423
rect 1026 1383 1029 1416
rect 1034 1403 1037 1416
rect 1014 1343 1021 1346
rect 986 1233 997 1236
rect 986 1176 989 1233
rect 994 1203 997 1216
rect 1002 1203 1005 1216
rect 1010 1213 1013 1336
rect 1018 1303 1021 1343
rect 1034 1293 1037 1326
rect 1042 1313 1045 2353
rect 1062 2336 1065 2493
rect 1074 2403 1077 2536
rect 1082 2523 1093 2526
rect 1098 2523 1101 2543
rect 1082 2413 1085 2516
rect 1106 2446 1109 2536
rect 1114 2513 1117 3006
rect 1122 2983 1125 3233
rect 1130 3213 1133 3226
rect 1138 3213 1141 3273
rect 1146 3233 1149 3623
rect 1154 3613 1157 3646
rect 1170 3586 1173 3956
rect 1178 3773 1181 3816
rect 1186 3756 1189 4016
rect 1194 3803 1197 3856
rect 1182 3753 1189 3756
rect 1182 3626 1185 3753
rect 1182 3623 1189 3626
rect 1194 3623 1197 3766
rect 1202 3746 1205 4173
rect 1250 4123 1253 4216
rect 1274 4213 1277 4226
rect 1290 4223 1293 4246
rect 1354 4243 1365 4246
rect 1282 4083 1285 4136
rect 1298 4103 1301 4136
rect 1282 4046 1285 4076
rect 1274 4043 1285 4046
rect 1218 4013 1221 4026
rect 1226 3956 1229 4036
rect 1258 4013 1261 4026
rect 1274 3996 1277 4043
rect 1274 3993 1285 3996
rect 1218 3953 1229 3956
rect 1218 3933 1221 3953
rect 1210 3763 1213 3826
rect 1218 3793 1221 3926
rect 1242 3923 1245 3936
rect 1202 3743 1209 3746
rect 1166 3583 1173 3586
rect 1166 3516 1169 3583
rect 1178 3523 1181 3606
rect 1186 3566 1189 3623
rect 1194 3583 1197 3606
rect 1206 3576 1209 3743
rect 1218 3613 1221 3726
rect 1242 3723 1245 3816
rect 1250 3763 1253 3806
rect 1258 3786 1261 3806
rect 1258 3783 1269 3786
rect 1282 3783 1285 3993
rect 1250 3733 1253 3746
rect 1266 3726 1269 3783
rect 1258 3723 1269 3726
rect 1258 3706 1261 3723
rect 1254 3703 1261 3706
rect 1254 3636 1257 3703
rect 1242 3623 1245 3636
rect 1254 3633 1261 3636
rect 1202 3573 1209 3576
rect 1186 3563 1193 3566
rect 1190 3516 1193 3563
rect 1166 3513 1173 3516
rect 1170 3456 1173 3513
rect 1166 3453 1173 3456
rect 1186 3513 1193 3516
rect 1186 3456 1189 3513
rect 1186 3453 1193 3456
rect 1154 3413 1157 3426
rect 1166 3376 1169 3453
rect 1190 3376 1193 3453
rect 1166 3373 1173 3376
rect 1154 3306 1157 3326
rect 1154 3303 1161 3306
rect 1158 3236 1161 3303
rect 1170 3253 1173 3373
rect 1186 3373 1193 3376
rect 1186 3323 1189 3373
rect 1202 3306 1205 3573
rect 1226 3533 1229 3606
rect 1250 3603 1253 3616
rect 1242 3533 1245 3546
rect 1250 3533 1253 3566
rect 1226 3493 1229 3526
rect 1258 3513 1261 3633
rect 1266 3596 1269 3686
rect 1290 3626 1293 3726
rect 1298 3723 1301 3896
rect 1306 3766 1309 4086
rect 1314 4073 1317 4226
rect 1322 4203 1325 4226
rect 1330 4213 1349 4216
rect 1354 4213 1357 4226
rect 1330 4123 1333 4206
rect 1346 4186 1349 4213
rect 1354 4193 1357 4206
rect 1362 4203 1365 4243
rect 1346 4183 1357 4186
rect 1354 4106 1357 4183
rect 1378 4126 1381 4346
rect 1442 4343 1445 4596
rect 1458 4413 1461 4526
rect 1474 4506 1477 4536
rect 1498 4523 1501 4556
rect 1506 4533 1509 4606
rect 1522 4553 1525 4616
rect 1578 4576 1581 4606
rect 1562 4573 1581 4576
rect 1514 4516 1517 4526
rect 1506 4513 1517 4516
rect 1474 4503 1485 4506
rect 1482 4426 1485 4503
rect 1474 4423 1485 4426
rect 1402 4213 1405 4226
rect 1346 4103 1357 4106
rect 1370 4123 1381 4126
rect 1346 3996 1349 4103
rect 1346 3993 1357 3996
rect 1314 3893 1317 3976
rect 1354 3973 1357 3993
rect 1370 3966 1373 4123
rect 1386 4103 1389 4136
rect 1394 4133 1397 4206
rect 1410 4203 1413 4316
rect 1426 4223 1445 4226
rect 1426 4213 1429 4223
rect 1418 4203 1429 4206
rect 1402 4123 1405 4196
rect 1434 4193 1437 4216
rect 1410 4113 1413 4136
rect 1434 4056 1437 4136
rect 1442 4123 1445 4223
rect 1450 4123 1453 4206
rect 1434 4053 1441 4056
rect 1418 3993 1421 4016
rect 1438 3976 1441 4053
rect 1362 3963 1373 3966
rect 1434 3973 1441 3976
rect 1346 3903 1349 3936
rect 1362 3933 1365 3963
rect 1434 3936 1437 3973
rect 1430 3933 1437 3936
rect 1450 3933 1453 4016
rect 1458 3946 1461 4336
rect 1474 4333 1477 4423
rect 1490 4333 1493 4406
rect 1466 4323 1485 4326
rect 1490 4213 1493 4306
rect 1498 4203 1501 4316
rect 1506 4306 1509 4513
rect 1514 4413 1517 4506
rect 1522 4406 1525 4476
rect 1562 4446 1565 4573
rect 1586 4533 1589 4546
rect 1594 4523 1597 4536
rect 1610 4533 1613 4616
rect 1650 4533 1653 4606
rect 1658 4533 1661 4616
rect 1666 4603 1669 4616
rect 1602 4513 1605 4526
rect 1618 4493 1621 4526
rect 1626 4513 1629 4526
rect 1682 4523 1685 4736
rect 1730 4553 1733 4646
rect 1794 4613 1797 4646
rect 1938 4636 1941 4726
rect 1934 4633 1941 4636
rect 1858 4613 1861 4626
rect 1562 4443 1581 4446
rect 1538 4413 1541 4426
rect 1514 4403 1525 4406
rect 1530 4393 1533 4406
rect 1546 4393 1549 4406
rect 1554 4403 1557 4416
rect 1562 4383 1565 4406
rect 1578 4343 1581 4443
rect 1602 4393 1605 4416
rect 1538 4333 1549 4336
rect 1626 4333 1629 4346
rect 1506 4303 1517 4306
rect 1514 4246 1517 4303
rect 1506 4243 1517 4246
rect 1546 4246 1549 4326
rect 1578 4313 1581 4326
rect 1642 4323 1645 4426
rect 1658 4333 1661 4416
rect 1546 4243 1557 4246
rect 1498 4113 1501 4126
rect 1458 3943 1477 3946
rect 1410 3913 1413 3926
rect 1314 3813 1317 3876
rect 1322 3793 1325 3826
rect 1330 3783 1333 3806
rect 1306 3763 1317 3766
rect 1314 3656 1317 3763
rect 1338 3723 1341 3796
rect 1354 3753 1357 3816
rect 1362 3803 1365 3896
rect 1430 3876 1433 3933
rect 1426 3873 1433 3876
rect 1370 3793 1373 3806
rect 1378 3723 1381 3816
rect 1410 3783 1413 3816
rect 1426 3796 1429 3873
rect 1442 3803 1445 3926
rect 1458 3903 1461 3926
rect 1474 3896 1477 3943
rect 1490 3933 1493 4016
rect 1498 3993 1501 4006
rect 1506 3926 1509 4243
rect 1514 4213 1517 4226
rect 1538 4196 1541 4206
rect 1554 4203 1557 4243
rect 1562 4196 1565 4216
rect 1570 4203 1573 4266
rect 1538 4193 1565 4196
rect 1514 3936 1517 4006
rect 1522 4003 1525 4016
rect 1514 3933 1525 3936
rect 1466 3893 1477 3896
rect 1498 3893 1501 3926
rect 1506 3923 1517 3926
rect 1426 3793 1437 3796
rect 1394 3723 1397 3746
rect 1418 3713 1421 3736
rect 1306 3653 1317 3656
rect 1290 3623 1301 3626
rect 1274 3613 1293 3616
rect 1298 3613 1301 3623
rect 1266 3593 1277 3596
rect 1210 3346 1213 3416
rect 1210 3343 1221 3346
rect 1194 3303 1205 3306
rect 1154 3233 1161 3236
rect 1194 3236 1197 3303
rect 1210 3246 1213 3326
rect 1218 3323 1221 3343
rect 1234 3303 1237 3406
rect 1210 3243 1221 3246
rect 1194 3233 1205 3236
rect 1154 3213 1157 3233
rect 1130 3186 1133 3206
rect 1130 3183 1137 3186
rect 1122 2716 1125 2936
rect 1134 2896 1137 3183
rect 1146 3163 1149 3206
rect 1154 3186 1157 3196
rect 1170 3193 1173 3206
rect 1178 3203 1181 3216
rect 1154 3183 1165 3186
rect 1146 3003 1149 3126
rect 1154 3083 1157 3146
rect 1154 3013 1157 3026
rect 1130 2893 1137 2896
rect 1130 2806 1133 2893
rect 1138 2813 1141 2876
rect 1130 2803 1141 2806
rect 1130 2733 1133 2746
rect 1122 2713 1129 2716
rect 1126 2646 1129 2713
rect 1126 2643 1133 2646
rect 1090 2443 1109 2446
rect 1074 2346 1077 2396
rect 1074 2343 1081 2346
rect 1050 2316 1053 2336
rect 1062 2333 1069 2336
rect 1050 2313 1057 2316
rect 1054 2226 1057 2313
rect 1050 2223 1057 2226
rect 1050 1813 1053 2223
rect 1058 2193 1061 2206
rect 1058 2003 1061 2136
rect 1058 1813 1061 1956
rect 1050 1786 1053 1806
rect 1050 1783 1057 1786
rect 1054 1446 1057 1783
rect 1050 1443 1057 1446
rect 1050 1213 1053 1443
rect 1066 1413 1069 2333
rect 1078 2156 1081 2343
rect 1074 2153 1081 2156
rect 1074 1833 1077 2153
rect 1082 2123 1085 2136
rect 1082 1583 1085 2076
rect 1090 1863 1093 2443
rect 1106 2413 1117 2416
rect 1098 2086 1101 2336
rect 1106 2306 1109 2406
rect 1114 2383 1117 2413
rect 1122 2376 1125 2616
rect 1130 2523 1133 2643
rect 1138 2506 1141 2803
rect 1146 2606 1149 2996
rect 1162 2993 1165 3183
rect 1170 3123 1173 3186
rect 1178 3133 1181 3166
rect 1186 3143 1189 3216
rect 1202 3166 1205 3233
rect 1198 3163 1205 3166
rect 1186 3113 1189 3136
rect 1198 3096 1201 3163
rect 1218 3156 1221 3243
rect 1210 3153 1221 3156
rect 1154 2903 1157 2976
rect 1154 2743 1157 2816
rect 1154 2723 1157 2736
rect 1162 2706 1165 2986
rect 1170 2813 1173 3086
rect 1178 3003 1181 3026
rect 1178 2806 1181 2936
rect 1170 2803 1181 2806
rect 1170 2723 1173 2803
rect 1186 2766 1189 3096
rect 1198 3093 1205 3096
rect 1210 3093 1213 3153
rect 1218 3123 1221 3136
rect 1202 3076 1205 3093
rect 1202 3073 1213 3076
rect 1210 2996 1213 3073
rect 1194 2966 1197 2996
rect 1202 2993 1213 2996
rect 1202 2973 1205 2993
rect 1194 2963 1205 2966
rect 1194 2913 1197 2926
rect 1202 2923 1205 2963
rect 1218 2913 1221 2956
rect 1234 2946 1237 3256
rect 1250 3193 1253 3426
rect 1258 3413 1261 3496
rect 1274 3406 1277 3593
rect 1290 3553 1293 3613
rect 1298 3533 1301 3606
rect 1306 3596 1309 3653
rect 1314 3613 1317 3636
rect 1394 3626 1397 3706
rect 1434 3703 1437 3793
rect 1466 3736 1469 3893
rect 1482 3813 1501 3816
rect 1506 3803 1509 3916
rect 1458 3733 1469 3736
rect 1482 3733 1485 3746
rect 1458 3676 1461 3733
rect 1466 3723 1477 3726
rect 1458 3673 1469 3676
rect 1394 3623 1401 3626
rect 1306 3593 1313 3596
rect 1310 3526 1313 3593
rect 1330 3533 1333 3606
rect 1354 3603 1357 3616
rect 1266 3403 1277 3406
rect 1266 3256 1269 3403
rect 1290 3363 1293 3526
rect 1306 3523 1313 3526
rect 1306 3436 1309 3523
rect 1322 3493 1325 3526
rect 1302 3433 1309 3436
rect 1282 3323 1285 3336
rect 1302 3326 1305 3433
rect 1314 3333 1317 3426
rect 1322 3393 1325 3406
rect 1290 3283 1293 3326
rect 1302 3323 1309 3326
rect 1306 3266 1309 3323
rect 1262 3253 1269 3256
rect 1298 3263 1309 3266
rect 1250 3123 1253 3146
rect 1250 3036 1253 3116
rect 1262 3096 1265 3253
rect 1274 3103 1277 3246
rect 1298 3186 1301 3263
rect 1298 3183 1309 3186
rect 1290 3133 1293 3166
rect 1262 3093 1269 3096
rect 1242 3033 1253 3036
rect 1242 3023 1245 3033
rect 1234 2943 1241 2946
rect 1226 2913 1229 2936
rect 1194 2833 1197 2866
rect 1182 2763 1189 2766
rect 1162 2703 1173 2706
rect 1154 2623 1157 2676
rect 1170 2636 1173 2703
rect 1182 2686 1185 2763
rect 1182 2683 1189 2686
rect 1162 2633 1173 2636
rect 1146 2603 1153 2606
rect 1134 2503 1141 2506
rect 1134 2426 1137 2503
rect 1150 2496 1153 2603
rect 1146 2493 1153 2496
rect 1134 2423 1141 2426
rect 1130 2393 1133 2406
rect 1114 2373 1125 2376
rect 1114 2323 1117 2373
rect 1138 2353 1141 2423
rect 1130 2316 1133 2326
rect 1122 2313 1133 2316
rect 1106 2303 1113 2306
rect 1110 2106 1113 2303
rect 1122 2213 1125 2313
rect 1138 2296 1141 2336
rect 1134 2293 1141 2296
rect 1134 2226 1137 2293
rect 1130 2223 1137 2226
rect 1122 2123 1125 2146
rect 1130 2106 1133 2223
rect 1138 2193 1141 2216
rect 1110 2103 1117 2106
rect 1098 2083 1105 2086
rect 1102 1866 1105 2083
rect 1098 1863 1105 1866
rect 1098 1843 1101 1863
rect 1114 1836 1117 2103
rect 1126 2103 1133 2106
rect 1126 2016 1129 2103
rect 1138 2023 1141 2126
rect 1146 2096 1149 2493
rect 1162 2416 1165 2633
rect 1170 2613 1181 2616
rect 1186 2546 1189 2683
rect 1178 2543 1189 2546
rect 1202 2546 1205 2906
rect 1238 2886 1241 2943
rect 1250 2916 1253 3033
rect 1250 2913 1261 2916
rect 1234 2883 1241 2886
rect 1210 2786 1213 2866
rect 1234 2863 1237 2883
rect 1250 2866 1253 2886
rect 1250 2863 1257 2866
rect 1226 2803 1229 2856
rect 1254 2796 1257 2863
rect 1250 2793 1257 2796
rect 1210 2783 1221 2786
rect 1210 2723 1213 2736
rect 1218 2653 1221 2783
rect 1226 2663 1229 2736
rect 1250 2733 1253 2793
rect 1218 2593 1221 2626
rect 1202 2543 1221 2546
rect 1178 2436 1181 2543
rect 1194 2516 1197 2536
rect 1190 2513 1197 2516
rect 1202 2513 1205 2526
rect 1190 2456 1193 2513
rect 1210 2466 1213 2536
rect 1218 2533 1221 2543
rect 1234 2533 1237 2606
rect 1250 2523 1253 2656
rect 1258 2623 1261 2646
rect 1202 2463 1213 2466
rect 1190 2453 1197 2456
rect 1178 2433 1189 2436
rect 1162 2413 1173 2416
rect 1186 2413 1189 2433
rect 1154 2363 1157 2406
rect 1154 2323 1157 2356
rect 1170 2346 1173 2413
rect 1194 2393 1197 2453
rect 1162 2343 1173 2346
rect 1162 2226 1165 2343
rect 1162 2223 1169 2226
rect 1178 2223 1181 2326
rect 1154 2113 1157 2216
rect 1166 2176 1169 2223
rect 1178 2193 1181 2206
rect 1202 2176 1205 2463
rect 1210 2423 1245 2426
rect 1234 2403 1237 2416
rect 1210 2376 1213 2396
rect 1210 2373 1229 2376
rect 1226 2266 1229 2373
rect 1166 2173 1173 2176
rect 1170 2106 1173 2173
rect 1162 2103 1173 2106
rect 1186 2173 1205 2176
rect 1218 2263 1229 2266
rect 1146 2093 1153 2096
rect 1150 2016 1153 2093
rect 1126 2013 1133 2016
rect 1130 1893 1133 2013
rect 1146 2013 1153 2016
rect 1130 1846 1133 1866
rect 1106 1833 1117 1836
rect 1126 1843 1133 1846
rect 1098 1723 1101 1746
rect 1090 1603 1093 1616
rect 1098 1613 1101 1656
rect 1098 1553 1101 1606
rect 1074 1513 1077 1536
rect 1098 1526 1101 1546
rect 1082 1503 1085 1526
rect 1094 1523 1101 1526
rect 1094 1436 1097 1523
rect 1094 1433 1101 1436
rect 1066 1393 1069 1406
rect 1066 1366 1069 1386
rect 1066 1363 1073 1366
rect 1058 1313 1061 1336
rect 1026 1193 1029 1206
rect 1058 1196 1061 1306
rect 1070 1236 1073 1363
rect 1082 1273 1085 1396
rect 1090 1323 1093 1416
rect 1098 1306 1101 1433
rect 1094 1303 1101 1306
rect 1042 1193 1061 1196
rect 1066 1233 1073 1236
rect 986 1173 1005 1176
rect 1002 1026 1005 1173
rect 1042 1166 1045 1193
rect 986 1023 1005 1026
rect 1026 1163 1045 1166
rect 986 1003 989 1023
rect 1026 1016 1029 1163
rect 1050 1136 1053 1176
rect 1042 1133 1053 1136
rect 1042 1036 1045 1133
rect 1058 1103 1061 1126
rect 1042 1033 1053 1036
rect 1026 1013 1037 1016
rect 1010 983 1013 996
rect 1034 946 1037 1013
rect 1034 943 1045 946
rect 994 913 997 926
rect 1018 923 1029 926
rect 1034 913 1037 926
rect 1042 906 1045 943
rect 1026 903 1045 906
rect 978 783 981 796
rect 1002 793 1005 806
rect 994 733 997 746
rect 1010 733 1013 746
rect 978 603 981 696
rect 978 573 981 596
rect 1002 593 1005 606
rect 1018 583 1021 616
rect 986 543 989 566
rect 1002 543 1013 546
rect 994 523 997 536
rect 1026 533 1029 903
rect 1042 793 1045 816
rect 1050 803 1053 1033
rect 1050 766 1053 786
rect 1042 763 1053 766
rect 1042 616 1045 763
rect 1042 613 1053 616
rect 1034 593 1045 596
rect 1034 523 1037 546
rect 1050 533 1053 613
rect 1058 603 1061 1066
rect 1066 906 1069 1233
rect 1074 1136 1077 1216
rect 1094 1146 1097 1303
rect 1094 1143 1101 1146
rect 1074 1133 1085 1136
rect 1074 1053 1077 1126
rect 1082 1123 1085 1133
rect 1098 1126 1101 1143
rect 1106 1133 1109 1833
rect 1114 1723 1117 1816
rect 1126 1776 1129 1843
rect 1126 1773 1133 1776
rect 1122 1716 1125 1736
rect 1114 1713 1125 1716
rect 1114 1613 1117 1713
rect 1130 1706 1133 1773
rect 1146 1766 1149 2013
rect 1162 1953 1165 2103
rect 1186 1976 1189 2173
rect 1218 2166 1221 2263
rect 1242 2226 1245 2246
rect 1210 2163 1221 2166
rect 1234 2223 1245 2226
rect 1210 2116 1213 2163
rect 1202 2113 1213 2116
rect 1202 1996 1205 2113
rect 1202 1993 1213 1996
rect 1186 1973 1205 1976
rect 1170 1933 1173 1946
rect 1154 1913 1157 1926
rect 1194 1913 1197 1926
rect 1202 1896 1205 1973
rect 1122 1703 1133 1706
rect 1142 1763 1149 1766
rect 1122 1606 1125 1703
rect 1142 1696 1145 1763
rect 1130 1676 1133 1696
rect 1142 1693 1149 1696
rect 1130 1673 1137 1676
rect 1118 1603 1125 1606
rect 1118 1466 1121 1603
rect 1134 1576 1137 1673
rect 1114 1463 1121 1466
rect 1130 1573 1137 1576
rect 1114 1316 1117 1463
rect 1122 1333 1125 1346
rect 1130 1333 1133 1573
rect 1146 1543 1149 1693
rect 1154 1536 1157 1846
rect 1170 1826 1173 1896
rect 1198 1893 1205 1896
rect 1170 1823 1177 1826
rect 1162 1603 1165 1816
rect 1174 1746 1177 1823
rect 1170 1743 1177 1746
rect 1146 1533 1157 1536
rect 1138 1503 1141 1526
rect 1138 1393 1141 1416
rect 1138 1343 1141 1386
rect 1114 1313 1125 1316
rect 1138 1313 1141 1326
rect 1098 1123 1109 1126
rect 1082 1096 1085 1116
rect 1082 1093 1093 1096
rect 1074 923 1077 1026
rect 1090 916 1093 1093
rect 1106 1056 1109 1123
rect 1102 1053 1109 1056
rect 1102 996 1105 1053
rect 1122 1046 1125 1313
rect 1146 1306 1149 1533
rect 1154 1513 1157 1526
rect 1162 1523 1165 1536
rect 1154 1333 1157 1416
rect 1170 1413 1173 1743
rect 1186 1736 1189 1836
rect 1198 1756 1201 1893
rect 1198 1753 1205 1756
rect 1186 1733 1193 1736
rect 1178 1693 1181 1726
rect 1190 1686 1193 1733
rect 1186 1683 1193 1686
rect 1178 1523 1181 1616
rect 1186 1513 1189 1683
rect 1170 1366 1173 1406
rect 1170 1363 1177 1366
rect 1162 1333 1165 1356
rect 1114 1043 1125 1046
rect 1138 1303 1149 1306
rect 1114 1003 1117 1043
rect 1122 1013 1125 1026
rect 1102 993 1109 996
rect 1082 913 1093 916
rect 1066 903 1073 906
rect 1070 816 1073 903
rect 1066 813 1073 816
rect 1066 733 1069 813
rect 1074 773 1077 796
rect 1082 783 1085 913
rect 1106 896 1109 993
rect 1138 973 1141 1303
rect 1162 1196 1165 1326
rect 1174 1286 1177 1363
rect 1174 1283 1181 1286
rect 1154 1193 1165 1196
rect 1154 1026 1157 1193
rect 1170 1176 1173 1276
rect 1166 1173 1173 1176
rect 1166 1046 1169 1173
rect 1166 1043 1173 1046
rect 1154 1023 1165 1026
rect 1154 986 1157 1006
rect 1146 983 1157 986
rect 1122 943 1141 946
rect 1122 933 1125 943
rect 1098 893 1109 896
rect 1130 893 1133 936
rect 1138 923 1141 943
rect 1146 923 1149 983
rect 1098 836 1101 893
rect 1098 833 1109 836
rect 1090 813 1101 816
rect 1106 803 1109 833
rect 1114 813 1117 886
rect 1074 723 1077 756
rect 1090 696 1093 746
rect 1114 726 1117 806
rect 1130 743 1133 876
rect 1114 723 1125 726
rect 1082 693 1093 696
rect 1066 613 1077 616
rect 1082 606 1085 693
rect 1066 603 1085 606
rect 1090 603 1093 616
rect 946 396 949 416
rect 954 403 957 416
rect 962 413 965 506
rect 1050 473 1053 526
rect 1066 523 1069 603
rect 978 413 981 426
rect 986 413 989 436
rect 1018 413 1021 426
rect 1090 406 1093 556
rect 1098 523 1101 616
rect 1106 506 1109 696
rect 1122 646 1125 723
rect 1114 643 1125 646
rect 1114 603 1117 643
rect 1130 603 1133 626
rect 1138 613 1141 726
rect 1154 693 1157 976
rect 1162 903 1165 1023
rect 1162 676 1165 856
rect 1158 673 1165 676
rect 1146 613 1149 656
rect 1158 596 1161 673
rect 1102 503 1109 506
rect 1102 426 1105 503
rect 1102 423 1109 426
rect 962 396 965 406
rect 930 393 941 396
rect 946 393 965 396
rect 938 386 941 393
rect 938 383 949 386
rect 922 343 941 346
rect 922 323 925 343
rect 914 313 925 316
rect 890 303 909 306
rect 858 213 861 236
rect 874 193 877 206
rect 810 123 813 166
rect 882 163 885 216
rect 834 133 837 156
rect 850 133 853 146
rect 874 123 877 136
rect 890 123 893 206
rect 898 193 901 206
rect 906 153 909 303
rect 914 133 917 216
rect 922 133 925 313
rect 930 253 933 336
rect 938 333 941 343
rect 938 213 941 326
rect 946 323 949 383
rect 1066 356 1069 406
rect 1090 403 1097 406
rect 1082 383 1085 396
rect 1094 356 1097 403
rect 1058 353 1069 356
rect 1058 333 1061 353
rect 1074 343 1077 356
rect 1090 353 1097 356
rect 946 293 949 316
rect 970 313 973 326
rect 978 303 981 326
rect 1010 313 1013 326
rect 898 123 909 126
rect 930 123 933 206
rect 954 196 957 216
rect 962 203 965 226
rect 970 213 973 286
rect 970 196 973 206
rect 954 193 973 196
rect 986 123 989 216
rect 1018 193 1021 206
rect 1074 203 1077 336
rect 1090 333 1093 353
rect 1106 333 1109 423
rect 1114 403 1117 576
rect 1122 403 1125 416
rect 1138 393 1141 526
rect 1146 523 1149 596
rect 1158 593 1165 596
rect 1162 573 1165 593
rect 1154 513 1157 536
rect 1162 413 1165 526
rect 1170 486 1173 1043
rect 1178 966 1181 1283
rect 1186 986 1189 1366
rect 1194 1113 1197 1636
rect 1202 1176 1205 1753
rect 1210 1706 1213 1993
rect 1218 1886 1221 2106
rect 1234 2046 1237 2223
rect 1250 2123 1253 2426
rect 1234 2043 1245 2046
rect 1234 2013 1237 2026
rect 1234 1993 1237 2006
rect 1242 1976 1245 2043
rect 1250 2006 1253 2116
rect 1266 2073 1269 3093
rect 1274 2893 1277 2936
rect 1290 2883 1293 3126
rect 1298 3063 1301 3136
rect 1298 2933 1301 2986
rect 1306 2846 1309 3183
rect 1314 3093 1317 3116
rect 1322 3113 1325 3316
rect 1338 3286 1341 3536
rect 1386 3523 1389 3616
rect 1398 3526 1401 3623
rect 1410 3543 1413 3626
rect 1426 3586 1429 3606
rect 1422 3583 1429 3586
rect 1450 3586 1453 3666
rect 1458 3603 1461 3616
rect 1450 3583 1457 3586
rect 1394 3523 1401 3526
rect 1394 3506 1397 3523
rect 1386 3503 1397 3506
rect 1386 3396 1389 3503
rect 1410 3486 1413 3526
rect 1422 3516 1425 3583
rect 1422 3513 1429 3516
rect 1402 3483 1413 3486
rect 1402 3426 1405 3483
rect 1402 3423 1413 3426
rect 1410 3403 1413 3423
rect 1418 3413 1421 3496
rect 1426 3403 1429 3513
rect 1386 3393 1397 3396
rect 1362 3303 1365 3336
rect 1338 3283 1349 3286
rect 1346 3216 1349 3283
rect 1338 3213 1349 3216
rect 1338 3193 1341 3213
rect 1362 3176 1365 3196
rect 1354 3173 1365 3176
rect 1338 3113 1341 3126
rect 1354 3116 1357 3173
rect 1370 3123 1373 3286
rect 1394 3223 1397 3393
rect 1434 3386 1437 3556
rect 1430 3383 1437 3386
rect 1410 3313 1413 3326
rect 1402 3276 1405 3306
rect 1402 3273 1413 3276
rect 1410 3216 1413 3273
rect 1430 3246 1433 3383
rect 1430 3243 1437 3246
rect 1402 3213 1413 3216
rect 1386 3133 1389 3156
rect 1354 3113 1365 3116
rect 1314 3003 1317 3046
rect 1330 3003 1333 3056
rect 1314 2916 1317 2966
rect 1322 2933 1325 2956
rect 1362 2943 1365 3113
rect 1378 3013 1381 3026
rect 1378 2923 1389 2926
rect 1314 2913 1325 2916
rect 1346 2913 1357 2916
rect 1302 2843 1309 2846
rect 1274 2793 1277 2816
rect 1274 2593 1277 2726
rect 1290 2723 1293 2806
rect 1302 2736 1305 2843
rect 1322 2836 1325 2913
rect 1314 2833 1325 2836
rect 1302 2733 1309 2736
rect 1290 2713 1301 2716
rect 1290 2656 1293 2713
rect 1282 2653 1293 2656
rect 1282 2623 1285 2653
rect 1282 2613 1301 2616
rect 1306 2603 1309 2733
rect 1314 2716 1317 2833
rect 1322 2733 1325 2816
rect 1338 2803 1341 2816
rect 1314 2713 1321 2716
rect 1354 2713 1357 2913
rect 1378 2816 1381 2836
rect 1370 2813 1381 2816
rect 1370 2756 1373 2813
rect 1370 2753 1377 2756
rect 1318 2596 1321 2713
rect 1282 2423 1285 2596
rect 1314 2593 1321 2596
rect 1314 2546 1317 2593
rect 1314 2543 1321 2546
rect 1298 2423 1301 2526
rect 1306 2416 1309 2536
rect 1318 2416 1321 2543
rect 1274 2393 1277 2416
rect 1290 2413 1309 2416
rect 1314 2413 1321 2416
rect 1282 2233 1285 2366
rect 1290 2056 1293 2413
rect 1298 2393 1301 2406
rect 1298 2203 1301 2326
rect 1306 2133 1309 2406
rect 1314 2306 1317 2413
rect 1322 2323 1325 2396
rect 1330 2386 1333 2686
rect 1362 2673 1365 2736
rect 1374 2626 1377 2753
rect 1374 2623 1381 2626
rect 1346 2593 1349 2606
rect 1338 2483 1341 2526
rect 1354 2516 1357 2556
rect 1370 2533 1373 2606
rect 1378 2596 1381 2623
rect 1386 2613 1389 2923
rect 1394 2833 1397 3066
rect 1402 3053 1405 3213
rect 1426 3076 1429 3226
rect 1418 3073 1429 3076
rect 1418 2976 1421 3073
rect 1418 2973 1429 2976
rect 1402 2936 1405 2956
rect 1426 2953 1429 2973
rect 1402 2933 1409 2936
rect 1406 2826 1409 2933
rect 1402 2823 1409 2826
rect 1378 2593 1385 2596
rect 1382 2526 1385 2593
rect 1378 2523 1385 2526
rect 1346 2443 1349 2516
rect 1354 2513 1365 2516
rect 1362 2446 1365 2513
rect 1354 2443 1365 2446
rect 1354 2426 1357 2443
rect 1350 2423 1357 2426
rect 1338 2403 1341 2416
rect 1330 2383 1337 2386
rect 1334 2316 1337 2383
rect 1350 2366 1353 2423
rect 1362 2373 1365 2426
rect 1370 2403 1373 2416
rect 1350 2363 1357 2366
rect 1354 2346 1357 2363
rect 1354 2343 1365 2346
rect 1330 2313 1337 2316
rect 1314 2303 1321 2306
rect 1290 2053 1297 2056
rect 1250 2003 1261 2006
rect 1274 2003 1277 2026
rect 1238 1973 1245 1976
rect 1238 1916 1241 1973
rect 1250 1923 1253 1996
rect 1258 1953 1261 2003
rect 1282 1923 1285 2046
rect 1294 1926 1297 2053
rect 1306 2003 1309 2116
rect 1318 1996 1321 2303
rect 1314 1993 1321 1996
rect 1314 1933 1317 1993
rect 1290 1923 1297 1926
rect 1306 1923 1317 1926
rect 1238 1913 1245 1916
rect 1218 1883 1229 1886
rect 1226 1733 1229 1883
rect 1242 1833 1245 1913
rect 1290 1903 1293 1923
rect 1306 1903 1309 1923
rect 1322 1886 1325 1916
rect 1314 1883 1325 1886
rect 1234 1813 1245 1816
rect 1234 1796 1237 1813
rect 1250 1803 1253 1826
rect 1274 1816 1277 1836
rect 1314 1826 1317 1883
rect 1314 1823 1325 1826
rect 1234 1793 1241 1796
rect 1218 1723 1229 1726
rect 1238 1716 1241 1793
rect 1258 1736 1261 1816
rect 1266 1803 1269 1816
rect 1274 1813 1285 1816
rect 1282 1746 1285 1813
rect 1274 1743 1285 1746
rect 1258 1733 1265 1736
rect 1234 1713 1241 1716
rect 1210 1703 1221 1706
rect 1218 1626 1221 1703
rect 1210 1623 1221 1626
rect 1210 1573 1213 1623
rect 1234 1613 1237 1713
rect 1250 1663 1253 1726
rect 1262 1636 1265 1733
rect 1274 1706 1277 1743
rect 1306 1733 1317 1736
rect 1322 1733 1325 1823
rect 1298 1723 1309 1726
rect 1274 1703 1285 1706
rect 1258 1633 1265 1636
rect 1258 1613 1261 1633
rect 1282 1626 1285 1703
rect 1274 1623 1285 1626
rect 1226 1533 1229 1606
rect 1234 1603 1245 1606
rect 1210 1303 1213 1526
rect 1218 1413 1221 1426
rect 1218 1253 1221 1326
rect 1210 1193 1213 1206
rect 1202 1173 1209 1176
rect 1206 1106 1209 1173
rect 1218 1133 1221 1216
rect 1226 1156 1229 1336
rect 1234 1323 1237 1566
rect 1242 1306 1245 1576
rect 1274 1563 1277 1623
rect 1250 1516 1253 1536
rect 1274 1533 1277 1556
rect 1250 1513 1257 1516
rect 1254 1446 1257 1513
rect 1250 1443 1257 1446
rect 1250 1413 1253 1443
rect 1258 1413 1261 1426
rect 1266 1403 1269 1526
rect 1274 1426 1277 1516
rect 1282 1443 1285 1526
rect 1298 1523 1301 1606
rect 1306 1506 1309 1626
rect 1298 1503 1309 1506
rect 1274 1423 1285 1426
rect 1258 1333 1261 1356
rect 1266 1333 1269 1346
rect 1250 1313 1253 1326
rect 1242 1303 1253 1306
rect 1266 1303 1269 1326
rect 1250 1246 1253 1303
rect 1282 1296 1285 1423
rect 1298 1306 1301 1503
rect 1298 1303 1309 1306
rect 1274 1293 1285 1296
rect 1274 1256 1277 1293
rect 1306 1283 1309 1303
rect 1314 1266 1317 1716
rect 1330 1616 1333 2313
rect 1346 2213 1349 2336
rect 1362 2266 1365 2343
rect 1358 2263 1365 2266
rect 1358 2206 1361 2263
rect 1378 2256 1381 2523
rect 1394 2386 1397 2616
rect 1402 2606 1405 2823
rect 1402 2603 1409 2606
rect 1406 2466 1409 2603
rect 1418 2586 1421 2946
rect 1434 2703 1437 3243
rect 1442 3223 1445 3546
rect 1454 3506 1457 3583
rect 1466 3533 1469 3673
rect 1498 3603 1501 3796
rect 1514 3713 1517 3923
rect 1522 3896 1525 3933
rect 1522 3893 1529 3896
rect 1526 3826 1529 3893
rect 1538 3873 1541 4136
rect 1554 4093 1557 4193
rect 1602 4186 1605 4276
rect 1666 4246 1669 4386
rect 1674 4313 1677 4336
rect 1682 4333 1685 4486
rect 1690 4453 1693 4536
rect 1722 4533 1733 4536
rect 1698 4376 1701 4416
rect 1746 4413 1749 4426
rect 1762 4413 1765 4546
rect 1810 4543 1813 4606
rect 1890 4573 1893 4616
rect 1898 4613 1901 4626
rect 1898 4566 1901 4606
rect 1890 4563 1901 4566
rect 1810 4513 1813 4526
rect 1850 4426 1853 4536
rect 1866 4523 1869 4546
rect 1874 4523 1877 4556
rect 1890 4523 1893 4563
rect 1906 4533 1909 4576
rect 1778 4393 1781 4416
rect 1786 4413 1789 4426
rect 1826 4423 1853 4426
rect 1802 4403 1805 4416
rect 1698 4373 1717 4376
rect 1658 4243 1669 4246
rect 1586 4183 1605 4186
rect 1562 4003 1565 4136
rect 1586 4046 1589 4183
rect 1610 4133 1613 4216
rect 1618 4133 1621 4196
rect 1642 4193 1645 4216
rect 1658 4156 1661 4243
rect 1658 4153 1669 4156
rect 1586 4043 1605 4046
rect 1570 3986 1573 4016
rect 1586 4013 1589 4026
rect 1566 3983 1573 3986
rect 1554 3836 1557 3926
rect 1566 3916 1569 3983
rect 1578 3933 1581 4006
rect 1594 4003 1597 4016
rect 1566 3913 1573 3916
rect 1570 3893 1573 3913
rect 1602 3856 1605 4043
rect 1610 4013 1613 4126
rect 1626 4023 1629 4126
rect 1634 4103 1637 4136
rect 1642 4003 1645 4136
rect 1658 4126 1661 4136
rect 1650 4123 1661 4126
rect 1666 4123 1669 4153
rect 1650 4106 1653 4123
rect 1650 4103 1661 4106
rect 1658 3996 1661 4103
rect 1674 4036 1677 4156
rect 1690 4133 1693 4256
rect 1706 4133 1709 4296
rect 1714 4276 1717 4373
rect 1826 4346 1829 4423
rect 1842 4396 1845 4406
rect 1850 4403 1853 4423
rect 1858 4396 1861 4416
rect 1842 4393 1861 4396
rect 1866 4393 1869 4406
rect 1826 4343 1837 4346
rect 1762 4323 1765 4336
rect 1794 4303 1797 4326
rect 1802 4323 1805 4336
rect 1714 4273 1721 4276
rect 1718 4216 1721 4273
rect 1810 4263 1813 4326
rect 1834 4316 1837 4343
rect 1842 4343 1861 4346
rect 1842 4333 1845 4343
rect 1850 4316 1853 4336
rect 1858 4323 1861 4343
rect 1834 4313 1853 4316
rect 1850 4236 1853 4313
rect 1866 4303 1869 4336
rect 1834 4233 1853 4236
rect 1714 4213 1721 4216
rect 1714 4176 1717 4213
rect 1738 4193 1741 4206
rect 1786 4193 1789 4216
rect 1818 4183 1821 4216
rect 1826 4213 1829 4226
rect 1714 4173 1721 4176
rect 1718 4126 1721 4173
rect 1770 4133 1773 4176
rect 1826 4136 1829 4206
rect 1834 4203 1837 4233
rect 1842 4213 1845 4226
rect 1850 4183 1853 4206
rect 1650 3993 1661 3996
rect 1670 4033 1677 4036
rect 1714 4123 1721 4126
rect 1610 3923 1613 3936
rect 1650 3923 1653 3993
rect 1670 3986 1673 4033
rect 1690 3993 1693 4006
rect 1670 3983 1677 3986
rect 1522 3823 1529 3826
rect 1538 3833 1557 3836
rect 1522 3636 1525 3823
rect 1530 3743 1533 3806
rect 1538 3793 1541 3833
rect 1554 3803 1557 3833
rect 1594 3853 1605 3856
rect 1626 3856 1629 3876
rect 1626 3853 1637 3856
rect 1530 3723 1533 3736
rect 1538 3733 1541 3756
rect 1546 3723 1549 3766
rect 1554 3733 1557 3796
rect 1578 3793 1581 3816
rect 1594 3776 1597 3853
rect 1634 3776 1637 3853
rect 1594 3773 1601 3776
rect 1570 3726 1573 3746
rect 1514 3633 1525 3636
rect 1514 3576 1517 3633
rect 1530 3603 1533 3616
rect 1498 3573 1517 3576
rect 1450 3503 1457 3506
rect 1450 3396 1453 3503
rect 1458 3413 1461 3486
rect 1490 3403 1493 3416
rect 1450 3393 1457 3396
rect 1454 3236 1457 3393
rect 1450 3233 1457 3236
rect 1442 3203 1445 3216
rect 1442 3123 1445 3136
rect 1450 3076 1453 3233
rect 1458 3203 1461 3216
rect 1466 3203 1469 3316
rect 1482 3216 1485 3326
rect 1474 3213 1485 3216
rect 1490 3203 1493 3216
rect 1498 3166 1501 3573
rect 1514 3523 1517 3536
rect 1522 3533 1525 3586
rect 1554 3583 1557 3616
rect 1530 3483 1533 3526
rect 1546 3436 1549 3536
rect 1562 3523 1565 3726
rect 1570 3723 1581 3726
rect 1578 3666 1581 3723
rect 1598 3706 1601 3773
rect 1626 3773 1637 3776
rect 1626 3736 1629 3773
rect 1666 3763 1669 3816
rect 1610 3713 1613 3736
rect 1618 3733 1629 3736
rect 1598 3703 1605 3706
rect 1570 3663 1581 3666
rect 1570 3456 1573 3663
rect 1602 3626 1605 3703
rect 1650 3666 1653 3726
rect 1646 3663 1653 3666
rect 1598 3623 1605 3626
rect 1578 3533 1581 3596
rect 1586 3523 1589 3536
rect 1598 3526 1601 3623
rect 1610 3533 1613 3616
rect 1626 3533 1629 3616
rect 1634 3613 1637 3636
rect 1646 3576 1649 3663
rect 1646 3573 1653 3576
rect 1674 3573 1677 3983
rect 1714 3976 1717 4123
rect 1730 4006 1733 4106
rect 1754 4046 1757 4126
rect 1762 4073 1765 4126
rect 1754 4043 1761 4046
rect 1738 4013 1741 4026
rect 1710 3973 1717 3976
rect 1710 3926 1713 3973
rect 1722 3933 1725 4006
rect 1730 4003 1741 4006
rect 1738 3946 1741 4003
rect 1758 3976 1761 4043
rect 1770 4013 1773 4126
rect 1778 4056 1781 4126
rect 1786 4123 1789 4136
rect 1778 4053 1789 4056
rect 1778 4013 1781 4026
rect 1786 4003 1789 4053
rect 1754 3973 1761 3976
rect 1738 3943 1745 3946
rect 1698 3913 1701 3926
rect 1710 3923 1717 3926
rect 1730 3923 1733 3936
rect 1690 3793 1693 3806
rect 1690 3733 1693 3746
rect 1682 3613 1685 3626
rect 1714 3603 1717 3923
rect 1730 3813 1733 3876
rect 1742 3866 1745 3943
rect 1738 3863 1745 3866
rect 1730 3723 1733 3786
rect 1738 3686 1741 3863
rect 1754 3856 1757 3973
rect 1762 3873 1765 3926
rect 1802 3923 1805 4126
rect 1810 4073 1813 4136
rect 1818 4133 1829 4136
rect 1754 3853 1765 3856
rect 1762 3776 1765 3853
rect 1794 3813 1797 3876
rect 1818 3846 1821 4133
rect 1858 4123 1861 4266
rect 1882 4263 1885 4426
rect 1906 4423 1909 4526
rect 1914 4513 1917 4526
rect 1866 4193 1869 4216
rect 1898 4203 1901 4226
rect 1906 4203 1909 4216
rect 1826 4013 1829 4106
rect 1866 4096 1869 4126
rect 1882 4123 1885 4136
rect 1858 4093 1869 4096
rect 1834 4003 1837 4086
rect 1858 4006 1861 4093
rect 1858 4003 1869 4006
rect 1826 3943 1845 3946
rect 1826 3933 1829 3943
rect 1826 3866 1829 3926
rect 1834 3873 1837 3936
rect 1842 3923 1845 3943
rect 1850 3923 1853 3936
rect 1858 3923 1861 3986
rect 1866 3913 1869 4003
rect 1874 3996 1877 4076
rect 1914 4066 1917 4416
rect 1922 4403 1925 4626
rect 1934 4586 1937 4633
rect 1954 4593 1957 4606
rect 2002 4603 2005 4616
rect 1934 4583 1941 4586
rect 1938 4566 1941 4583
rect 1938 4563 1949 4566
rect 1930 4523 1933 4536
rect 1946 4446 1949 4563
rect 1970 4543 1989 4546
rect 1970 4533 1973 4543
rect 1970 4483 1973 4526
rect 1978 4523 1981 4536
rect 1986 4523 1989 4543
rect 1994 4533 1997 4586
rect 2034 4533 2037 4616
rect 2042 4603 2045 4616
rect 2002 4493 2005 4526
rect 2066 4523 2069 4606
rect 2074 4523 2077 4536
rect 2082 4473 2085 4526
rect 2106 4503 2109 4666
rect 2642 4656 2645 4726
rect 2642 4653 2649 4656
rect 2138 4593 2141 4606
rect 2186 4603 2189 4616
rect 2122 4533 2125 4576
rect 2146 4533 2149 4546
rect 2170 4536 2173 4596
rect 2166 4533 2173 4536
rect 2218 4533 2221 4616
rect 2226 4603 2229 4616
rect 2234 4586 2237 4606
rect 2226 4583 2237 4586
rect 2138 4513 2141 4526
rect 1938 4443 1949 4446
rect 1930 4413 1933 4426
rect 1938 4406 1941 4443
rect 1930 4403 1941 4406
rect 1930 4333 1933 4403
rect 1946 4396 1949 4426
rect 1938 4393 1949 4396
rect 1938 4296 1941 4393
rect 1954 4333 1957 4416
rect 1962 4403 1965 4416
rect 1986 4323 1989 4356
rect 1994 4323 1997 4336
rect 1994 4303 1997 4316
rect 1938 4293 1957 4296
rect 1930 4236 1933 4266
rect 1954 4236 1957 4293
rect 1922 4233 1933 4236
rect 1946 4233 1957 4236
rect 1922 4203 1925 4233
rect 1938 4153 1941 4216
rect 1938 4133 1941 4146
rect 1946 4106 1949 4233
rect 1954 4183 1957 4206
rect 1962 4166 1965 4216
rect 1970 4183 1973 4206
rect 1978 4203 1981 4226
rect 1986 4213 1989 4276
rect 2002 4216 2005 4376
rect 2010 4353 2013 4416
rect 2050 4393 2053 4406
rect 2018 4346 2021 4366
rect 2066 4346 2069 4416
rect 2010 4343 2021 4346
rect 2062 4343 2069 4346
rect 2010 4333 2013 4343
rect 2010 4323 2021 4326
rect 2026 4286 2029 4336
rect 2034 4293 2037 4336
rect 2026 4283 2037 4286
rect 1994 4213 2005 4216
rect 1962 4163 1973 4166
rect 2010 4163 2013 4206
rect 2026 4196 2029 4206
rect 2034 4203 2037 4283
rect 2042 4213 2045 4326
rect 2050 4216 2053 4326
rect 2062 4296 2065 4343
rect 2090 4336 2093 4406
rect 2114 4396 2117 4416
rect 2122 4403 2125 4436
rect 2130 4396 2133 4406
rect 2114 4393 2133 4396
rect 2074 4333 2093 4336
rect 2074 4306 2077 4333
rect 2098 4323 2101 4336
rect 2074 4303 2093 4306
rect 2138 4303 2141 4456
rect 2154 4443 2157 4526
rect 2166 4416 2169 4533
rect 2178 4453 2181 4526
rect 2226 4523 2229 4583
rect 2194 4456 2197 4476
rect 2194 4453 2201 4456
rect 2166 4413 2173 4416
rect 2178 4413 2181 4426
rect 2186 4413 2189 4436
rect 2062 4293 2069 4296
rect 2050 4213 2061 4216
rect 2050 4196 2053 4206
rect 2026 4193 2053 4196
rect 1898 4063 1917 4066
rect 1938 4103 1949 4106
rect 1882 4013 1885 4046
rect 1874 3993 1885 3996
rect 1882 3906 1885 3993
rect 1898 3956 1901 4063
rect 1826 3863 1837 3866
rect 1810 3843 1821 3846
rect 1754 3773 1765 3776
rect 1802 3773 1805 3816
rect 1754 3706 1757 3773
rect 1810 3756 1813 3843
rect 1818 3793 1821 3816
rect 1770 3723 1773 3736
rect 1778 3713 1781 3756
rect 1802 3753 1813 3756
rect 1786 3733 1789 3746
rect 1754 3703 1765 3706
rect 1738 3683 1749 3686
rect 1730 3613 1733 3626
rect 1650 3536 1653 3573
rect 1650 3533 1661 3536
rect 1674 3533 1685 3536
rect 1598 3523 1605 3526
rect 1650 3523 1653 3533
rect 1542 3433 1549 3436
rect 1562 3453 1573 3456
rect 1514 3303 1517 3406
rect 1490 3163 1501 3166
rect 1490 3116 1493 3163
rect 1514 3123 1517 3156
rect 1490 3113 1501 3116
rect 1450 3073 1461 3076
rect 1442 2983 1445 3016
rect 1458 2956 1461 3073
rect 1498 3046 1501 3113
rect 1450 2953 1461 2956
rect 1482 3043 1501 3046
rect 1482 2956 1485 3043
rect 1522 3036 1525 3206
rect 1530 3203 1533 3366
rect 1542 3236 1545 3433
rect 1562 3426 1565 3453
rect 1554 3423 1565 3426
rect 1542 3233 1549 3236
rect 1506 3033 1525 3036
rect 1482 2953 1493 2956
rect 1450 2746 1453 2953
rect 1458 2903 1461 2926
rect 1466 2913 1469 2936
rect 1490 2836 1493 2953
rect 1506 2886 1509 3033
rect 1514 2983 1517 3016
rect 1522 3003 1525 3026
rect 1538 3013 1541 3216
rect 1546 3106 1549 3233
rect 1554 3203 1557 3423
rect 1562 3366 1565 3416
rect 1562 3363 1573 3366
rect 1570 3226 1573 3363
rect 1562 3223 1573 3226
rect 1562 3206 1565 3223
rect 1586 3213 1589 3326
rect 1602 3306 1605 3523
rect 1674 3453 1677 3533
rect 1706 3516 1709 3576
rect 1698 3513 1709 3516
rect 1698 3436 1701 3513
rect 1722 3456 1725 3526
rect 1730 3493 1733 3576
rect 1738 3533 1741 3676
rect 1746 3666 1749 3683
rect 1746 3663 1753 3666
rect 1750 3566 1753 3663
rect 1746 3563 1753 3566
rect 1746 3526 1749 3563
rect 1762 3546 1765 3703
rect 1802 3656 1805 3753
rect 1802 3653 1813 3656
rect 1738 3523 1749 3526
rect 1754 3543 1765 3546
rect 1722 3453 1729 3456
rect 1698 3433 1705 3436
rect 1626 3323 1629 3416
rect 1658 3393 1661 3406
rect 1666 3333 1669 3376
rect 1674 3333 1677 3346
rect 1682 3306 1685 3326
rect 1602 3303 1613 3306
rect 1610 3216 1613 3303
rect 1674 3303 1685 3306
rect 1674 3236 1677 3303
rect 1674 3233 1685 3236
rect 1610 3213 1621 3216
rect 1562 3203 1581 3206
rect 1570 3133 1581 3136
rect 1554 3123 1573 3126
rect 1586 3106 1589 3206
rect 1594 3193 1597 3206
rect 1594 3123 1597 3156
rect 1546 3103 1557 3106
rect 1554 3036 1557 3103
rect 1546 3033 1557 3036
rect 1578 3103 1589 3106
rect 1538 2933 1541 2966
rect 1530 2903 1533 2926
rect 1546 2886 1549 3033
rect 1578 3016 1581 3103
rect 1506 2883 1517 2886
rect 1490 2833 1501 2836
rect 1458 2803 1461 2826
rect 1466 2813 1477 2816
rect 1446 2743 1453 2746
rect 1446 2676 1449 2743
rect 1458 2726 1461 2736
rect 1466 2733 1469 2806
rect 1482 2793 1485 2806
rect 1458 2723 1477 2726
rect 1458 2683 1461 2723
rect 1434 2603 1437 2676
rect 1446 2673 1453 2676
rect 1450 2653 1453 2673
rect 1418 2583 1437 2586
rect 1418 2533 1429 2536
rect 1418 2476 1421 2533
rect 1418 2473 1425 2476
rect 1406 2463 1413 2466
rect 1410 2443 1413 2463
rect 1422 2426 1425 2473
rect 1434 2463 1437 2583
rect 1458 2566 1461 2606
rect 1450 2563 1461 2566
rect 1450 2486 1453 2563
rect 1466 2493 1469 2706
rect 1474 2596 1477 2656
rect 1482 2613 1485 2736
rect 1490 2723 1493 2816
rect 1498 2803 1501 2833
rect 1514 2826 1517 2883
rect 1506 2823 1517 2826
rect 1538 2883 1549 2886
rect 1506 2783 1509 2823
rect 1538 2816 1541 2883
rect 1538 2813 1549 2816
rect 1530 2733 1533 2796
rect 1546 2716 1549 2813
rect 1554 2803 1557 3016
rect 1578 3013 1589 3016
rect 1562 2976 1565 2996
rect 1562 2973 1569 2976
rect 1566 2896 1569 2973
rect 1586 2956 1589 3013
rect 1594 3003 1597 3116
rect 1618 3076 1621 3213
rect 1602 3073 1621 3076
rect 1602 2976 1605 3073
rect 1618 2993 1621 3056
rect 1642 3046 1645 3136
rect 1674 3133 1677 3206
rect 1682 3163 1685 3233
rect 1690 3203 1693 3416
rect 1702 3376 1705 3433
rect 1726 3376 1729 3453
rect 1702 3373 1709 3376
rect 1706 3226 1709 3373
rect 1722 3373 1729 3376
rect 1722 3246 1725 3373
rect 1738 3356 1741 3523
rect 1754 3426 1757 3543
rect 1778 3533 1781 3636
rect 1786 3613 1789 3626
rect 1786 3596 1789 3606
rect 1794 3603 1797 3636
rect 1802 3596 1805 3616
rect 1786 3593 1805 3596
rect 1810 3583 1813 3653
rect 1754 3423 1761 3426
rect 1746 3373 1749 3416
rect 1758 3356 1761 3423
rect 1734 3353 1741 3356
rect 1754 3353 1761 3356
rect 1734 3266 1737 3353
rect 1754 3333 1757 3353
rect 1770 3343 1773 3526
rect 1786 3516 1789 3566
rect 1818 3536 1821 3746
rect 1826 3733 1829 3806
rect 1834 3623 1837 3863
rect 1842 3783 1845 3816
rect 1858 3636 1861 3906
rect 1854 3633 1861 3636
rect 1874 3903 1885 3906
rect 1894 3953 1901 3956
rect 1894 3906 1897 3953
rect 1894 3903 1901 3906
rect 1826 3593 1829 3616
rect 1842 3576 1845 3596
rect 1854 3586 1857 3633
rect 1874 3623 1877 3903
rect 1882 3803 1893 3806
rect 1882 3793 1885 3803
rect 1898 3736 1901 3903
rect 1914 3883 1917 4056
rect 1938 3903 1941 4103
rect 1970 4096 1973 4163
rect 1962 4093 1973 4096
rect 1962 4036 1965 4093
rect 1962 4033 1973 4036
rect 1946 3923 1949 4016
rect 1914 3803 1917 3876
rect 1922 3813 1933 3816
rect 1938 3813 1941 3836
rect 1890 3733 1901 3736
rect 1922 3733 1925 3813
rect 1930 3803 1941 3806
rect 1946 3786 1949 3826
rect 1938 3783 1949 3786
rect 1890 3653 1893 3733
rect 1874 3603 1877 3616
rect 1854 3583 1861 3586
rect 1794 3533 1805 3536
rect 1814 3533 1821 3536
rect 1838 3573 1845 3576
rect 1782 3513 1789 3516
rect 1782 3356 1785 3513
rect 1802 3486 1805 3526
rect 1794 3483 1805 3486
rect 1782 3353 1789 3356
rect 1734 3263 1741 3266
rect 1722 3243 1733 3246
rect 1706 3223 1713 3226
rect 1642 3043 1653 3046
rect 1650 2996 1653 3043
rect 1666 3013 1669 3056
rect 1682 3043 1685 3126
rect 1690 3053 1693 3136
rect 1698 3123 1701 3216
rect 1710 3116 1713 3223
rect 1706 3113 1713 3116
rect 1706 3026 1709 3113
rect 1722 3096 1725 3236
rect 1698 3023 1709 3026
rect 1718 3093 1725 3096
rect 1642 2993 1653 2996
rect 1602 2973 1629 2976
rect 1578 2933 1581 2956
rect 1586 2953 1597 2956
rect 1578 2913 1581 2926
rect 1594 2906 1597 2953
rect 1618 2923 1621 2966
rect 1586 2903 1597 2906
rect 1566 2893 1573 2896
rect 1570 2826 1573 2893
rect 1562 2823 1573 2826
rect 1538 2713 1549 2716
rect 1538 2636 1541 2713
rect 1538 2633 1549 2636
rect 1474 2593 1481 2596
rect 1478 2486 1481 2593
rect 1490 2533 1493 2546
rect 1450 2483 1461 2486
rect 1418 2423 1425 2426
rect 1418 2403 1421 2423
rect 1442 2413 1445 2426
rect 1458 2403 1461 2483
rect 1474 2483 1481 2486
rect 1490 2523 1501 2526
rect 1386 2383 1397 2386
rect 1386 2363 1389 2383
rect 1394 2356 1397 2376
rect 1394 2353 1405 2356
rect 1402 2266 1405 2353
rect 1394 2263 1405 2266
rect 1378 2253 1385 2256
rect 1354 2203 1361 2206
rect 1354 2146 1357 2203
rect 1382 2176 1385 2253
rect 1378 2173 1385 2176
rect 1378 2146 1381 2173
rect 1354 2143 1365 2146
rect 1346 2116 1349 2136
rect 1338 2013 1341 2116
rect 1346 2113 1353 2116
rect 1350 2046 1353 2113
rect 1346 2043 1353 2046
rect 1346 2023 1349 2043
rect 1362 2016 1365 2143
rect 1354 2013 1365 2016
rect 1374 2143 1381 2146
rect 1394 2146 1397 2263
rect 1402 2193 1405 2216
rect 1426 2203 1429 2236
rect 1394 2143 1413 2146
rect 1442 2143 1445 2186
rect 1338 1916 1341 1936
rect 1338 1913 1345 1916
rect 1342 1736 1345 1913
rect 1338 1733 1345 1736
rect 1338 1713 1341 1733
rect 1354 1633 1357 2013
rect 1374 2006 1377 2143
rect 1386 2106 1389 2136
rect 1386 2103 1397 2106
rect 1394 2056 1397 2103
rect 1386 2053 1397 2056
rect 1386 2013 1389 2053
rect 1410 2036 1413 2143
rect 1450 2133 1453 2146
rect 1458 2123 1461 2166
rect 1466 2153 1469 2256
rect 1402 2033 1413 2036
rect 1474 2033 1477 2483
rect 1490 2413 1493 2523
rect 1506 2516 1509 2536
rect 1506 2513 1513 2516
rect 1498 2396 1501 2496
rect 1510 2446 1513 2513
rect 1522 2493 1525 2616
rect 1546 2613 1549 2633
rect 1554 2613 1557 2686
rect 1562 2673 1565 2823
rect 1578 2743 1581 2806
rect 1562 2593 1565 2616
rect 1530 2533 1533 2546
rect 1570 2543 1573 2646
rect 1530 2483 1533 2516
rect 1546 2513 1549 2526
rect 1506 2443 1513 2446
rect 1506 2423 1509 2443
rect 1506 2413 1517 2416
rect 1490 2393 1501 2396
rect 1490 2246 1493 2393
rect 1490 2243 1501 2246
rect 1482 2213 1485 2226
rect 1482 2133 1485 2206
rect 1490 2193 1493 2206
rect 1374 2003 1381 2006
rect 1370 1923 1373 1936
rect 1378 1906 1381 2003
rect 1402 1976 1405 2033
rect 1394 1973 1405 1976
rect 1370 1903 1381 1906
rect 1370 1826 1373 1903
rect 1362 1823 1373 1826
rect 1362 1726 1365 1823
rect 1370 1813 1381 1816
rect 1370 1733 1373 1813
rect 1386 1773 1389 1926
rect 1394 1876 1397 1973
rect 1394 1873 1401 1876
rect 1398 1756 1401 1873
rect 1418 1863 1421 1946
rect 1426 1833 1429 2016
rect 1458 2003 1461 2026
rect 1490 2023 1493 2126
rect 1466 1973 1469 2006
rect 1474 1996 1477 2016
rect 1474 1993 1481 1996
rect 1458 1933 1461 1946
rect 1434 1813 1437 1926
rect 1478 1906 1481 1993
rect 1474 1903 1481 1906
rect 1490 1903 1493 1926
rect 1394 1753 1401 1756
rect 1394 1733 1397 1753
rect 1362 1723 1381 1726
rect 1378 1696 1381 1723
rect 1394 1713 1397 1726
rect 1410 1723 1413 1806
rect 1378 1693 1397 1696
rect 1346 1616 1349 1626
rect 1330 1613 1337 1616
rect 1346 1613 1357 1616
rect 1322 1523 1325 1606
rect 1334 1546 1337 1613
rect 1362 1603 1365 1616
rect 1370 1613 1373 1636
rect 1394 1606 1397 1693
rect 1418 1653 1421 1736
rect 1434 1633 1437 1726
rect 1442 1696 1445 1716
rect 1442 1693 1449 1696
rect 1378 1603 1397 1606
rect 1330 1543 1337 1546
rect 1330 1506 1333 1543
rect 1346 1536 1349 1586
rect 1346 1533 1353 1536
rect 1326 1503 1333 1506
rect 1326 1386 1329 1503
rect 1338 1453 1341 1526
rect 1350 1466 1353 1533
rect 1346 1463 1353 1466
rect 1346 1393 1349 1463
rect 1378 1416 1381 1603
rect 1394 1433 1397 1526
rect 1418 1426 1421 1576
rect 1434 1533 1437 1616
rect 1446 1546 1449 1693
rect 1466 1656 1469 1816
rect 1474 1813 1477 1903
rect 1498 1896 1501 2243
rect 1506 2133 1509 2406
rect 1522 2286 1525 2466
rect 1538 2436 1541 2506
rect 1562 2456 1565 2536
rect 1534 2433 1541 2436
rect 1558 2453 1565 2456
rect 1534 2316 1537 2433
rect 1546 2323 1549 2426
rect 1534 2313 1541 2316
rect 1522 2283 1529 2286
rect 1514 2163 1517 2276
rect 1526 2226 1529 2283
rect 1522 2223 1529 2226
rect 1506 2113 1509 2126
rect 1506 2006 1509 2106
rect 1514 2013 1517 2156
rect 1506 2003 1517 2006
rect 1498 1893 1509 1896
rect 1514 1876 1517 2003
rect 1498 1873 1517 1876
rect 1498 1786 1501 1873
rect 1522 1793 1525 2223
rect 1538 2216 1541 2313
rect 1558 2306 1561 2453
rect 1554 2303 1561 2306
rect 1554 2236 1557 2303
rect 1554 2233 1565 2236
rect 1538 2213 1545 2216
rect 1530 1933 1533 2206
rect 1542 2116 1545 2213
rect 1554 2133 1557 2216
rect 1562 2116 1565 2233
rect 1570 2166 1573 2446
rect 1578 2253 1581 2526
rect 1586 2396 1589 2903
rect 1594 2813 1597 2826
rect 1594 2803 1605 2806
rect 1594 2723 1597 2803
rect 1610 2766 1613 2816
rect 1606 2763 1613 2766
rect 1606 2706 1609 2763
rect 1626 2733 1629 2973
rect 1642 2913 1645 2993
rect 1666 2933 1669 2996
rect 1698 2976 1701 3023
rect 1718 3006 1721 3093
rect 1718 3003 1725 3006
rect 1722 2983 1725 3003
rect 1698 2973 1709 2976
rect 1706 2936 1709 2973
rect 1698 2933 1709 2936
rect 1698 2856 1701 2933
rect 1698 2853 1709 2856
rect 1706 2836 1709 2853
rect 1642 2803 1645 2836
rect 1602 2703 1609 2706
rect 1602 2556 1605 2703
rect 1602 2553 1613 2556
rect 1594 2513 1597 2526
rect 1594 2413 1597 2426
rect 1586 2393 1593 2396
rect 1590 2236 1593 2393
rect 1602 2366 1605 2406
rect 1610 2393 1613 2553
rect 1618 2506 1621 2666
rect 1626 2523 1629 2606
rect 1650 2603 1653 2746
rect 1666 2723 1669 2826
rect 1674 2803 1677 2816
rect 1682 2813 1685 2836
rect 1698 2833 1709 2836
rect 1698 2776 1701 2833
rect 1698 2773 1709 2776
rect 1682 2713 1685 2736
rect 1706 2733 1709 2773
rect 1714 2696 1717 2716
rect 1706 2693 1717 2696
rect 1706 2636 1709 2693
rect 1706 2633 1717 2636
rect 1658 2613 1677 2616
rect 1666 2516 1669 2606
rect 1682 2523 1685 2606
rect 1690 2533 1693 2616
rect 1714 2603 1717 2633
rect 1722 2553 1725 2926
rect 1730 2576 1733 3243
rect 1738 2996 1741 3263
rect 1746 3216 1749 3326
rect 1754 3233 1757 3326
rect 1746 3213 1757 3216
rect 1746 3193 1749 3206
rect 1746 3133 1749 3186
rect 1746 3013 1749 3046
rect 1738 2993 1745 2996
rect 1742 2846 1745 2993
rect 1754 2923 1757 3213
rect 1762 3183 1765 3276
rect 1770 3163 1773 3266
rect 1778 3246 1781 3336
rect 1786 3263 1789 3353
rect 1794 3333 1797 3483
rect 1802 3413 1805 3456
rect 1814 3426 1817 3533
rect 1814 3423 1821 3426
rect 1802 3323 1805 3336
rect 1778 3243 1789 3246
rect 1770 3073 1773 3136
rect 1786 3066 1789 3243
rect 1802 3196 1805 3306
rect 1798 3193 1805 3196
rect 1798 3096 1801 3193
rect 1810 3103 1813 3406
rect 1798 3093 1805 3096
rect 1778 3063 1789 3066
rect 1778 3023 1781 3063
rect 1778 3006 1781 3016
rect 1778 3003 1789 3006
rect 1762 2933 1773 2936
rect 1738 2843 1745 2846
rect 1738 2713 1741 2843
rect 1746 2813 1749 2826
rect 1770 2783 1773 2806
rect 1754 2733 1757 2766
rect 1770 2733 1781 2736
rect 1786 2726 1789 2986
rect 1802 2836 1805 3093
rect 1818 3086 1821 3423
rect 1826 3413 1829 3526
rect 1838 3506 1841 3573
rect 1858 3563 1861 3583
rect 1898 3566 1901 3626
rect 1906 3613 1909 3726
rect 1938 3676 1941 3783
rect 1938 3673 1949 3676
rect 1922 3626 1925 3646
rect 1918 3623 1925 3626
rect 1874 3563 1901 3566
rect 1918 3566 1921 3623
rect 1938 3566 1941 3656
rect 1946 3593 1949 3673
rect 1954 3643 1957 4026
rect 1970 3976 1973 4033
rect 1994 3993 1997 4006
rect 2010 3983 2013 4006
rect 2026 4003 2029 4126
rect 1962 3973 1973 3976
rect 1962 3823 1965 3973
rect 1962 3743 1965 3816
rect 1970 3793 1973 3886
rect 1994 3836 1997 3926
rect 2042 3906 2045 4016
rect 2058 4013 2061 4213
rect 2066 4006 2069 4293
rect 2090 4186 2093 4303
rect 2146 4213 2149 4326
rect 2170 4256 2173 4413
rect 2198 4406 2201 4453
rect 2218 4413 2221 4426
rect 2194 4403 2201 4406
rect 2194 4346 2197 4403
rect 2194 4343 2205 4346
rect 2202 4296 2205 4343
rect 2218 4303 2221 4326
rect 2194 4293 2205 4296
rect 2170 4253 2181 4256
rect 2178 4193 2181 4253
rect 2034 3903 2045 3906
rect 2050 4003 2069 4006
rect 2074 4183 2093 4186
rect 2034 3856 2037 3903
rect 2034 3853 2045 3856
rect 1986 3833 1997 3836
rect 1986 3803 1989 3833
rect 2002 3793 2005 3806
rect 1962 3733 1981 3736
rect 1954 3613 1957 3626
rect 1962 3616 1965 3676
rect 1962 3613 1973 3616
rect 1978 3613 1981 3733
rect 1986 3723 1989 3766
rect 2018 3746 2021 3796
rect 2026 3763 2029 3816
rect 2018 3743 2029 3746
rect 1994 3703 1997 3736
rect 2026 3726 2029 3743
rect 2034 3733 2037 3786
rect 2010 3713 2013 3726
rect 2018 3723 2029 3726
rect 1962 3583 1965 3606
rect 1918 3563 1925 3566
rect 1938 3563 1949 3566
rect 1838 3503 1845 3506
rect 1842 3483 1845 3503
rect 1834 3413 1837 3446
rect 1866 3413 1869 3526
rect 1874 3456 1877 3563
rect 1906 3533 1909 3556
rect 1922 3546 1925 3563
rect 1922 3543 1933 3546
rect 1882 3476 1885 3496
rect 1882 3473 1893 3476
rect 1874 3453 1881 3456
rect 1878 3406 1881 3453
rect 1826 3393 1829 3406
rect 1842 3356 1845 3406
rect 1834 3353 1845 3356
rect 1826 3313 1829 3326
rect 1834 3323 1837 3353
rect 1842 3336 1845 3353
rect 1874 3403 1881 3406
rect 1842 3333 1853 3336
rect 1842 3306 1845 3326
rect 1838 3303 1845 3306
rect 1794 2833 1805 2836
rect 1814 3083 1821 3086
rect 1794 2796 1797 2833
rect 1802 2813 1805 2826
rect 1814 2806 1817 3083
rect 1826 3036 1829 3296
rect 1838 3236 1841 3303
rect 1838 3233 1845 3236
rect 1842 3213 1845 3233
rect 1834 3133 1837 3206
rect 1850 3203 1853 3333
rect 1866 3313 1869 3326
rect 1874 3293 1877 3403
rect 1890 3376 1893 3473
rect 1914 3413 1917 3486
rect 1930 3466 1933 3543
rect 1922 3463 1933 3466
rect 1882 3373 1893 3376
rect 1882 3276 1885 3373
rect 1874 3273 1885 3276
rect 1826 3033 1837 3036
rect 1826 2813 1829 3026
rect 1814 2803 1821 2806
rect 1794 2793 1801 2796
rect 1762 2723 1789 2726
rect 1786 2706 1789 2723
rect 1778 2703 1789 2706
rect 1746 2576 1749 2656
rect 1778 2636 1781 2703
rect 1798 2696 1801 2793
rect 1818 2746 1821 2803
rect 1834 2786 1837 3033
rect 1842 3013 1845 3126
rect 1858 3123 1861 3216
rect 1874 3166 1877 3273
rect 1890 3176 1893 3356
rect 1922 3353 1925 3463
rect 1946 3446 1949 3563
rect 1970 3493 1973 3613
rect 1986 3603 1989 3626
rect 1994 3613 1997 3676
rect 1986 3496 1989 3596
rect 1982 3493 1989 3496
rect 1938 3443 1949 3446
rect 1982 3446 1985 3493
rect 1982 3443 1989 3446
rect 1914 3216 1917 3346
rect 1930 3303 1933 3416
rect 1938 3306 1941 3443
rect 1986 3426 1989 3443
rect 1994 3433 1997 3486
rect 1954 3423 1981 3426
rect 1986 3423 1993 3426
rect 1946 3396 1949 3406
rect 1954 3403 1957 3423
rect 1962 3396 1965 3416
rect 1970 3403 1973 3416
rect 1978 3403 1981 3423
rect 1946 3393 1965 3396
rect 1990 3346 1993 3423
rect 1954 3333 1957 3346
rect 1990 3343 1997 3346
rect 1938 3303 1949 3306
rect 1914 3213 1925 3216
rect 1890 3173 1897 3176
rect 1874 3163 1885 3166
rect 1866 3123 1869 3146
rect 1882 3106 1885 3163
rect 1842 2903 1845 2936
rect 1850 2836 1853 2926
rect 1842 2833 1853 2836
rect 1858 2833 1861 3106
rect 1874 3103 1885 3106
rect 1874 2946 1877 3103
rect 1894 3096 1897 3173
rect 1890 3093 1897 3096
rect 1890 2956 1893 3093
rect 1898 3013 1901 3026
rect 1890 2953 1897 2956
rect 1874 2943 1885 2946
rect 1874 2893 1877 2926
rect 1842 2803 1845 2833
rect 1834 2783 1853 2786
rect 1858 2783 1861 2806
rect 1850 2766 1853 2783
rect 1882 2766 1885 2943
rect 1894 2836 1897 2953
rect 1906 2923 1909 3206
rect 1922 3146 1925 3213
rect 1946 3203 1949 3303
rect 1986 3213 1989 3326
rect 1994 3276 1997 3343
rect 2002 3293 2005 3656
rect 2018 3553 2021 3723
rect 2042 3626 2045 3853
rect 2050 3653 2053 4003
rect 2058 3923 2061 3996
rect 2074 3936 2077 4183
rect 2082 4033 2085 4126
rect 2082 3996 2085 4016
rect 2090 4003 2093 4016
rect 2098 4013 2101 4076
rect 2106 4053 2109 4166
rect 2122 4063 2125 4126
rect 2138 4116 2141 4136
rect 2178 4123 2181 4176
rect 2186 4133 2189 4146
rect 2138 4113 2149 4116
rect 2130 4046 2133 4096
rect 2122 4043 2133 4046
rect 2106 4013 2109 4036
rect 2098 3996 2101 4006
rect 2082 3993 2101 3996
rect 2122 3996 2125 4043
rect 2146 4036 2149 4113
rect 2186 4106 2189 4126
rect 2138 4033 2149 4036
rect 2178 4103 2189 4106
rect 2178 4036 2181 4103
rect 2178 4033 2189 4036
rect 2138 4003 2141 4033
rect 2122 3993 2133 3996
rect 2066 3933 2077 3936
rect 2066 3736 2069 3933
rect 2082 3923 2085 3986
rect 2074 3816 2077 3836
rect 2074 3813 2081 3816
rect 2078 3746 2081 3813
rect 2058 3733 2069 3736
rect 2074 3743 2081 3746
rect 2058 3646 2061 3733
rect 2074 3723 2077 3743
rect 2090 3733 2093 3816
rect 2082 3703 2085 3726
rect 2098 3703 2101 3766
rect 2106 3756 2109 3936
rect 2130 3846 2133 3993
rect 2146 3983 2149 4016
rect 2186 4013 2189 4033
rect 2146 3956 2149 3976
rect 2146 3953 2157 3956
rect 2154 3866 2157 3953
rect 2146 3863 2157 3866
rect 2130 3843 2137 3846
rect 2134 3786 2137 3843
rect 2134 3783 2141 3786
rect 2106 3753 2117 3756
rect 2114 3736 2117 3753
rect 2058 3643 2065 3646
rect 2042 3623 2053 3626
rect 2026 3523 2029 3536
rect 2042 3523 2045 3616
rect 2010 3413 2013 3436
rect 2018 3276 2021 3456
rect 1994 3273 2005 3276
rect 2002 3206 2005 3273
rect 1918 3143 1925 3146
rect 1918 3096 1921 3143
rect 1930 3103 1933 3136
rect 1938 3133 1941 3156
rect 1938 3106 1941 3126
rect 1954 3123 1957 3206
rect 1970 3123 1973 3206
rect 1994 3203 2005 3206
rect 2014 3273 2021 3276
rect 1994 3116 1997 3203
rect 2014 3186 2017 3273
rect 2026 3253 2029 3466
rect 2034 3413 2037 3496
rect 2050 3433 2053 3623
rect 2062 3566 2065 3643
rect 2082 3566 2085 3696
rect 2106 3633 2109 3736
rect 2114 3733 2121 3736
rect 2130 3733 2133 3776
rect 2118 3666 2121 3733
rect 2114 3663 2121 3666
rect 2062 3563 2069 3566
rect 2058 3393 2061 3446
rect 2066 3403 2069 3563
rect 2078 3563 2085 3566
rect 2050 3333 2053 3346
rect 2078 3336 2081 3563
rect 2090 3533 2093 3626
rect 2098 3536 2101 3616
rect 2114 3603 2117 3663
rect 2138 3566 2141 3783
rect 2122 3563 2141 3566
rect 2098 3533 2109 3536
rect 2090 3413 2093 3526
rect 2106 3456 2109 3533
rect 2098 3453 2109 3456
rect 2122 3456 2125 3563
rect 2146 3466 2149 3863
rect 2154 3813 2157 3836
rect 2154 3733 2165 3736
rect 2170 3733 2173 3746
rect 2154 3723 2165 3726
rect 2178 3656 2181 3826
rect 2186 3763 2189 3816
rect 2178 3653 2185 3656
rect 2154 3613 2157 3626
rect 2146 3463 2153 3466
rect 2122 3453 2141 3456
rect 2074 3333 2081 3336
rect 2034 3296 2037 3326
rect 2034 3293 2045 3296
rect 2042 3226 2045 3293
rect 2066 3256 2069 3296
rect 2074 3263 2077 3333
rect 2066 3253 2077 3256
rect 2026 3203 2029 3226
rect 2034 3223 2045 3226
rect 2010 3183 2017 3186
rect 2010 3126 2013 3183
rect 2034 3166 2037 3223
rect 2066 3213 2069 3236
rect 2026 3163 2037 3166
rect 2026 3133 2029 3163
rect 2042 3153 2045 3206
rect 2010 3123 2021 3126
rect 1986 3113 1997 3116
rect 1938 3103 1965 3106
rect 1918 3093 1925 3096
rect 1850 2763 1861 2766
rect 1818 2743 1825 2746
rect 1794 2693 1801 2696
rect 1778 2633 1789 2636
rect 1778 2593 1781 2616
rect 1730 2573 1737 2576
rect 1746 2573 1757 2576
rect 1666 2513 1693 2516
rect 1618 2503 1637 2506
rect 1634 2376 1637 2503
rect 1690 2456 1693 2513
rect 1686 2453 1693 2456
rect 1666 2403 1669 2416
rect 1674 2403 1677 2416
rect 1626 2373 1637 2376
rect 1686 2376 1689 2453
rect 1714 2443 1717 2536
rect 1734 2506 1737 2573
rect 1730 2503 1737 2506
rect 1686 2373 1693 2376
rect 1602 2363 1613 2366
rect 1610 2323 1613 2363
rect 1626 2316 1629 2373
rect 1618 2313 1629 2316
rect 1618 2243 1621 2313
rect 1586 2233 1593 2236
rect 1570 2163 1577 2166
rect 1542 2113 1549 2116
rect 1546 2026 1549 2113
rect 1538 2023 1549 2026
rect 1558 2113 1565 2116
rect 1530 1863 1533 1926
rect 1498 1783 1509 1786
rect 1506 1716 1509 1783
rect 1530 1723 1533 1816
rect 1538 1796 1541 2023
rect 1558 2016 1561 2113
rect 1574 2106 1577 2163
rect 1570 2103 1577 2106
rect 1570 2026 1573 2103
rect 1570 2023 1577 2026
rect 1558 2013 1565 2016
rect 1546 1916 1549 2006
rect 1562 1993 1565 2013
rect 1546 1913 1557 1916
rect 1546 1813 1549 1906
rect 1538 1793 1545 1796
rect 1542 1716 1545 1793
rect 1506 1713 1517 1716
rect 1466 1653 1477 1656
rect 1474 1576 1477 1653
rect 1490 1613 1493 1626
rect 1442 1543 1449 1546
rect 1466 1573 1477 1576
rect 1514 1573 1517 1713
rect 1538 1713 1545 1716
rect 1538 1636 1541 1713
rect 1538 1633 1545 1636
rect 1530 1613 1533 1626
rect 1466 1543 1469 1573
rect 1442 1523 1445 1543
rect 1414 1423 1421 1426
rect 1326 1383 1333 1386
rect 1330 1363 1333 1383
rect 1322 1333 1333 1336
rect 1306 1263 1317 1266
rect 1274 1253 1285 1256
rect 1250 1243 1261 1246
rect 1234 1213 1237 1226
rect 1234 1193 1237 1206
rect 1226 1153 1245 1156
rect 1234 1126 1237 1146
rect 1230 1123 1237 1126
rect 1202 1103 1209 1106
rect 1194 993 1197 1016
rect 1186 983 1197 986
rect 1178 963 1185 966
rect 1182 896 1185 963
rect 1178 893 1185 896
rect 1178 873 1181 893
rect 1178 813 1181 836
rect 1194 803 1197 983
rect 1178 646 1181 736
rect 1186 723 1189 736
rect 1194 733 1197 746
rect 1194 703 1197 726
rect 1178 643 1197 646
rect 1178 576 1181 616
rect 1186 603 1189 636
rect 1178 573 1189 576
rect 1178 503 1181 526
rect 1186 523 1189 573
rect 1194 533 1197 643
rect 1202 596 1205 1103
rect 1210 976 1213 1016
rect 1218 1003 1221 1106
rect 1230 1036 1233 1123
rect 1230 1033 1237 1036
rect 1210 973 1221 976
rect 1210 806 1213 936
rect 1218 913 1221 973
rect 1226 933 1229 996
rect 1218 816 1221 906
rect 1226 873 1229 926
rect 1234 923 1237 1033
rect 1218 813 1229 816
rect 1234 813 1237 826
rect 1210 803 1221 806
rect 1210 733 1221 736
rect 1210 633 1213 726
rect 1226 706 1229 813
rect 1242 743 1245 1153
rect 1258 1026 1261 1243
rect 1282 1186 1285 1253
rect 1306 1196 1309 1263
rect 1322 1213 1325 1326
rect 1338 1286 1341 1326
rect 1346 1303 1349 1336
rect 1354 1313 1357 1336
rect 1370 1323 1373 1416
rect 1378 1413 1389 1416
rect 1386 1316 1389 1413
rect 1414 1366 1417 1423
rect 1378 1313 1389 1316
rect 1402 1363 1417 1366
rect 1338 1283 1349 1286
rect 1346 1236 1349 1283
rect 1338 1233 1349 1236
rect 1322 1203 1333 1206
rect 1306 1193 1317 1196
rect 1274 1183 1285 1186
rect 1274 1166 1277 1183
rect 1270 1163 1277 1166
rect 1270 1096 1273 1163
rect 1290 1133 1293 1166
rect 1314 1146 1317 1193
rect 1314 1143 1325 1146
rect 1338 1143 1341 1233
rect 1378 1216 1381 1313
rect 1378 1213 1385 1216
rect 1354 1146 1357 1166
rect 1354 1143 1361 1146
rect 1322 1096 1325 1143
rect 1338 1123 1341 1136
rect 1270 1093 1277 1096
rect 1274 1076 1277 1093
rect 1314 1093 1325 1096
rect 1274 1073 1285 1076
rect 1258 1023 1265 1026
rect 1250 923 1253 1016
rect 1262 966 1265 1023
rect 1282 976 1285 1073
rect 1314 1026 1317 1093
rect 1358 1086 1361 1143
rect 1370 1103 1373 1206
rect 1382 1156 1385 1213
rect 1402 1163 1405 1363
rect 1426 1353 1429 1416
rect 1434 1403 1437 1456
rect 1426 1213 1429 1326
rect 1466 1313 1469 1526
rect 1482 1523 1485 1536
rect 1490 1513 1493 1536
rect 1482 1413 1485 1426
rect 1490 1403 1493 1446
rect 1498 1406 1501 1546
rect 1530 1533 1533 1606
rect 1542 1566 1545 1633
rect 1538 1563 1545 1566
rect 1506 1413 1509 1436
rect 1498 1403 1509 1406
rect 1474 1343 1493 1346
rect 1474 1333 1477 1343
rect 1378 1153 1385 1156
rect 1258 963 1265 966
rect 1274 973 1285 976
rect 1306 1023 1317 1026
rect 1354 1083 1361 1086
rect 1306 976 1309 1023
rect 1306 973 1317 976
rect 1250 813 1253 876
rect 1258 853 1261 963
rect 1266 933 1269 946
rect 1274 926 1277 973
rect 1266 923 1277 926
rect 1258 813 1261 836
rect 1266 806 1269 923
rect 1258 803 1269 806
rect 1226 703 1237 706
rect 1234 646 1237 703
rect 1226 643 1237 646
rect 1210 613 1213 626
rect 1226 616 1229 643
rect 1258 626 1261 803
rect 1250 623 1261 626
rect 1226 613 1237 616
rect 1202 593 1209 596
rect 1218 593 1221 606
rect 1206 526 1209 593
rect 1202 523 1209 526
rect 1170 483 1181 486
rect 1178 416 1181 483
rect 1202 456 1205 523
rect 1218 513 1221 526
rect 1202 453 1213 456
rect 1170 413 1181 416
rect 1082 203 1085 216
rect 1090 213 1093 246
rect 1098 203 1101 236
rect 1010 133 1013 156
rect 1050 133 1053 146
rect 1074 133 1077 156
rect 1106 143 1109 216
rect 1114 213 1117 346
rect 1130 333 1133 386
rect 1122 303 1125 326
rect 1138 273 1141 346
rect 1146 323 1149 336
rect 1162 323 1165 346
rect 1170 333 1173 413
rect 1130 213 1133 226
rect 1058 113 1061 126
rect 1098 113 1101 126
rect 1138 123 1141 216
rect 1146 186 1149 206
rect 1154 203 1157 256
rect 1162 196 1165 216
rect 1170 203 1173 216
rect 1178 213 1181 226
rect 1178 196 1181 206
rect 1154 186 1157 196
rect 1162 193 1181 196
rect 1146 183 1157 186
rect 1154 123 1157 183
rect 1186 133 1189 396
rect 1210 376 1213 453
rect 1226 413 1229 536
rect 1234 523 1237 613
rect 1234 413 1237 446
rect 1250 406 1253 623
rect 1274 616 1277 916
rect 1282 803 1285 826
rect 1282 733 1285 796
rect 1290 773 1293 816
rect 1298 783 1301 806
rect 1266 613 1285 616
rect 1266 526 1269 613
rect 1282 603 1293 606
rect 1274 533 1285 536
rect 1266 523 1277 526
rect 1274 506 1277 523
rect 1274 503 1281 506
rect 1250 403 1261 406
rect 1258 383 1261 403
rect 1202 373 1213 376
rect 1202 333 1205 373
rect 1250 333 1253 356
rect 1266 333 1269 476
rect 1278 406 1281 503
rect 1274 403 1281 406
rect 1290 403 1293 576
rect 1298 513 1301 726
rect 1314 696 1317 973
rect 1330 923 1333 1016
rect 1354 903 1357 1083
rect 1378 946 1381 1153
rect 1386 1123 1389 1136
rect 1418 1013 1421 1166
rect 1434 1143 1453 1146
rect 1434 1133 1437 1143
rect 1442 1103 1445 1136
rect 1450 1123 1453 1143
rect 1466 1136 1469 1226
rect 1482 1213 1485 1336
rect 1490 1323 1493 1343
rect 1498 1333 1501 1386
rect 1490 1203 1493 1256
rect 1466 1133 1477 1136
rect 1418 996 1421 1006
rect 1426 1003 1429 1016
rect 1434 996 1437 1016
rect 1466 1013 1469 1126
rect 1474 1093 1477 1133
rect 1418 993 1437 996
rect 1442 983 1445 1006
rect 1378 943 1385 946
rect 1370 856 1373 936
rect 1346 853 1373 856
rect 1338 796 1341 816
rect 1346 803 1349 853
rect 1354 813 1357 846
rect 1354 796 1357 806
rect 1338 793 1357 796
rect 1322 733 1325 746
rect 1338 733 1341 766
rect 1362 723 1365 816
rect 1370 763 1373 853
rect 1382 756 1385 943
rect 1394 873 1397 926
rect 1402 883 1405 936
rect 1418 866 1421 936
rect 1426 933 1429 946
rect 1466 913 1469 926
rect 1474 916 1477 1036
rect 1482 933 1485 1126
rect 1506 1103 1509 1403
rect 1522 1333 1525 1356
rect 1538 1316 1541 1563
rect 1554 1523 1557 1913
rect 1562 1713 1565 1986
rect 1574 1886 1577 2023
rect 1586 1903 1589 2233
rect 1594 2203 1597 2216
rect 1634 2203 1637 2226
rect 1658 2223 1661 2336
rect 1674 2313 1677 2366
rect 1666 2136 1669 2266
rect 1690 2153 1693 2373
rect 1714 2326 1717 2396
rect 1722 2333 1725 2416
rect 1706 2143 1709 2326
rect 1714 2323 1725 2326
rect 1722 2213 1725 2323
rect 1730 2306 1733 2503
rect 1754 2403 1757 2573
rect 1778 2486 1781 2556
rect 1774 2483 1781 2486
rect 1774 2376 1777 2483
rect 1770 2373 1777 2376
rect 1738 2323 1741 2336
rect 1730 2303 1741 2306
rect 1610 2063 1613 2136
rect 1642 2133 1669 2136
rect 1714 2133 1717 2206
rect 1642 2123 1645 2133
rect 1650 2083 1653 2126
rect 1682 2083 1685 2126
rect 1626 2013 1629 2066
rect 1738 2063 1741 2303
rect 1754 2123 1757 2336
rect 1770 2326 1773 2373
rect 1786 2333 1789 2633
rect 1794 2376 1797 2693
rect 1810 2643 1813 2736
rect 1822 2646 1825 2743
rect 1834 2733 1845 2736
rect 1818 2643 1825 2646
rect 1802 2513 1805 2526
rect 1818 2486 1821 2643
rect 1826 2613 1829 2626
rect 1834 2573 1837 2726
rect 1858 2706 1861 2763
rect 1850 2703 1861 2706
rect 1874 2763 1885 2766
rect 1890 2833 1897 2836
rect 1850 2683 1853 2703
rect 1874 2636 1877 2763
rect 1890 2746 1893 2833
rect 1886 2743 1893 2746
rect 1886 2676 1889 2743
rect 1898 2733 1901 2816
rect 1898 2683 1901 2726
rect 1906 2703 1909 2906
rect 1914 2723 1917 2736
rect 1886 2673 1893 2676
rect 1874 2633 1885 2636
rect 1842 2593 1845 2616
rect 1850 2573 1853 2616
rect 1874 2583 1877 2616
rect 1882 2566 1885 2633
rect 1874 2563 1885 2566
rect 1810 2483 1821 2486
rect 1826 2533 1845 2536
rect 1802 2393 1805 2466
rect 1794 2373 1801 2376
rect 1798 2326 1801 2373
rect 1810 2343 1813 2483
rect 1826 2413 1829 2533
rect 1834 2486 1837 2526
rect 1842 2513 1845 2526
rect 1850 2503 1853 2556
rect 1834 2483 1845 2486
rect 1842 2426 1845 2483
rect 1874 2446 1877 2563
rect 1890 2546 1893 2673
rect 1922 2653 1925 3093
rect 1946 3013 1949 3026
rect 1954 2996 1957 3096
rect 1962 3086 1965 3103
rect 1962 3083 1969 3086
rect 1966 3006 1969 3083
rect 1986 3066 1989 3113
rect 1986 3063 1997 3066
rect 1950 2993 1957 2996
rect 1962 3003 1969 3006
rect 1930 2726 1933 2896
rect 1938 2733 1941 2936
rect 1950 2926 1953 2993
rect 1962 2963 1965 3003
rect 1950 2923 1957 2926
rect 1946 2803 1949 2906
rect 1954 2813 1957 2923
rect 1962 2833 1965 2936
rect 1970 2923 1973 2986
rect 1986 2973 1989 3026
rect 1994 2906 1997 3063
rect 2002 2933 2005 3106
rect 1994 2903 2005 2906
rect 1970 2796 1973 2816
rect 1978 2803 1981 2826
rect 1986 2813 1989 2896
rect 2002 2836 2005 2903
rect 1994 2833 2005 2836
rect 1986 2796 1989 2806
rect 1994 2803 1997 2833
rect 2018 2826 2021 3123
rect 2018 2823 2025 2826
rect 1970 2793 1989 2796
rect 1930 2723 1941 2726
rect 1938 2706 1941 2723
rect 1938 2703 1949 2706
rect 1898 2596 1901 2606
rect 1906 2603 1909 2626
rect 1914 2596 1917 2616
rect 1930 2613 1933 2666
rect 1946 2636 1949 2703
rect 1938 2633 1949 2636
rect 1938 2613 1941 2633
rect 1978 2626 1981 2706
rect 1986 2636 1989 2786
rect 2010 2723 2013 2816
rect 2022 2716 2025 2823
rect 2018 2713 2025 2716
rect 1986 2633 2005 2636
rect 1978 2623 1989 2626
rect 1898 2593 1917 2596
rect 1886 2543 1893 2546
rect 1886 2466 1889 2543
rect 1886 2463 1893 2466
rect 1874 2443 1885 2446
rect 1842 2423 1853 2426
rect 1818 2373 1821 2406
rect 1850 2403 1853 2423
rect 1834 2346 1837 2396
rect 1830 2343 1837 2346
rect 1770 2323 1781 2326
rect 1778 2306 1781 2323
rect 1794 2323 1801 2326
rect 1778 2303 1785 2306
rect 1770 2256 1773 2286
rect 1766 2253 1773 2256
rect 1766 2186 1769 2253
rect 1782 2246 1785 2303
rect 1778 2243 1785 2246
rect 1766 2183 1773 2186
rect 1762 2106 1765 2166
rect 1754 2103 1765 2106
rect 1754 2046 1757 2103
rect 1754 2043 1765 2046
rect 1610 1923 1613 2006
rect 1642 1923 1645 1936
rect 1574 1883 1581 1886
rect 1578 1706 1581 1883
rect 1570 1703 1581 1706
rect 1570 1573 1573 1703
rect 1562 1403 1565 1426
rect 1578 1363 1581 1526
rect 1594 1446 1597 1866
rect 1618 1813 1621 1826
rect 1602 1723 1605 1736
rect 1618 1733 1621 1746
rect 1610 1693 1613 1726
rect 1626 1646 1629 1806
rect 1642 1783 1645 1816
rect 1650 1736 1653 1806
rect 1666 1803 1669 2016
rect 1698 1793 1701 1936
rect 1714 1923 1717 2016
rect 1746 1993 1749 2006
rect 1762 1966 1765 2043
rect 1746 1963 1765 1966
rect 1706 1783 1709 1806
rect 1714 1743 1717 1816
rect 1722 1803 1725 1856
rect 1746 1836 1749 1963
rect 1770 1846 1773 2183
rect 1778 2163 1781 2243
rect 1794 2146 1797 2323
rect 1818 2313 1821 2336
rect 1830 2296 1833 2343
rect 1818 2293 1833 2296
rect 1818 2176 1821 2293
rect 1818 2173 1837 2176
rect 1794 2143 1801 2146
rect 1786 2123 1789 2136
rect 1798 2086 1801 2143
rect 1834 2133 1837 2173
rect 1842 2166 1845 2336
rect 1850 2283 1853 2396
rect 1858 2333 1861 2426
rect 1882 2393 1885 2443
rect 1866 2313 1869 2326
rect 1882 2296 1885 2316
rect 1874 2293 1885 2296
rect 1874 2196 1877 2293
rect 1874 2193 1885 2196
rect 1882 2173 1885 2193
rect 1842 2163 1853 2166
rect 1798 2083 1805 2086
rect 1778 2003 1781 2056
rect 1802 1996 1805 2083
rect 1794 1993 1805 1996
rect 1794 1946 1797 1993
rect 1786 1943 1797 1946
rect 1786 1866 1789 1943
rect 1802 1876 1805 1936
rect 1802 1873 1809 1876
rect 1786 1863 1797 1866
rect 1770 1843 1777 1846
rect 1746 1833 1765 1836
rect 1730 1803 1733 1816
rect 1650 1733 1661 1736
rect 1634 1706 1637 1726
rect 1634 1703 1645 1706
rect 1618 1643 1629 1646
rect 1602 1513 1605 1526
rect 1594 1443 1605 1446
rect 1602 1376 1605 1443
rect 1586 1373 1605 1376
rect 1530 1313 1541 1316
rect 1530 1246 1533 1313
rect 1546 1283 1549 1326
rect 1554 1323 1557 1336
rect 1578 1316 1581 1336
rect 1530 1243 1541 1246
rect 1522 1213 1525 1226
rect 1514 1203 1525 1206
rect 1522 1113 1525 1203
rect 1530 1193 1533 1206
rect 1538 1196 1541 1243
rect 1546 1203 1549 1226
rect 1538 1193 1545 1196
rect 1490 923 1493 1006
rect 1498 923 1501 936
rect 1506 933 1509 1016
rect 1530 1013 1533 1126
rect 1542 1096 1545 1193
rect 1554 1163 1557 1316
rect 1570 1313 1581 1316
rect 1570 1246 1573 1313
rect 1586 1256 1589 1373
rect 1594 1333 1605 1336
rect 1610 1333 1613 1376
rect 1602 1313 1605 1326
rect 1618 1283 1621 1643
rect 1642 1636 1645 1703
rect 1634 1633 1645 1636
rect 1626 1503 1629 1526
rect 1634 1523 1637 1633
rect 1642 1513 1645 1526
rect 1658 1506 1661 1733
rect 1690 1653 1693 1726
rect 1698 1723 1701 1736
rect 1642 1503 1661 1506
rect 1642 1456 1645 1503
rect 1642 1453 1649 1456
rect 1626 1413 1629 1426
rect 1646 1376 1649 1453
rect 1642 1373 1649 1376
rect 1634 1313 1637 1326
rect 1642 1316 1645 1373
rect 1650 1323 1653 1336
rect 1658 1333 1661 1436
rect 1666 1413 1669 1426
rect 1698 1333 1701 1406
rect 1706 1353 1709 1616
rect 1714 1503 1717 1736
rect 1722 1723 1725 1796
rect 1730 1733 1733 1786
rect 1754 1733 1757 1806
rect 1762 1746 1765 1833
rect 1774 1766 1777 1843
rect 1774 1763 1781 1766
rect 1762 1743 1769 1746
rect 1738 1666 1741 1726
rect 1738 1663 1749 1666
rect 1730 1533 1733 1616
rect 1738 1583 1741 1606
rect 1746 1566 1749 1663
rect 1754 1613 1757 1726
rect 1766 1656 1769 1743
rect 1762 1653 1769 1656
rect 1762 1633 1765 1653
rect 1738 1563 1749 1566
rect 1738 1466 1741 1563
rect 1746 1533 1749 1556
rect 1754 1523 1757 1546
rect 1762 1533 1765 1616
rect 1778 1576 1781 1763
rect 1794 1736 1797 1863
rect 1806 1806 1809 1873
rect 1818 1813 1821 1926
rect 1826 1923 1829 2066
rect 1806 1803 1821 1806
rect 1770 1573 1781 1576
rect 1790 1733 1797 1736
rect 1790 1576 1793 1733
rect 1790 1573 1797 1576
rect 1730 1463 1741 1466
rect 1730 1413 1733 1463
rect 1730 1396 1733 1406
rect 1738 1403 1741 1436
rect 1746 1396 1749 1416
rect 1754 1403 1757 1506
rect 1770 1456 1773 1573
rect 1778 1533 1781 1546
rect 1770 1453 1777 1456
rect 1730 1393 1749 1396
rect 1642 1313 1661 1316
rect 1586 1253 1593 1256
rect 1570 1243 1581 1246
rect 1570 1213 1573 1226
rect 1578 1193 1581 1243
rect 1590 1176 1593 1253
rect 1610 1213 1613 1226
rect 1590 1173 1605 1176
rect 1570 1133 1573 1166
rect 1586 1106 1589 1146
rect 1586 1103 1597 1106
rect 1542 1093 1549 1096
rect 1546 956 1549 1093
rect 1570 993 1573 1006
rect 1538 953 1549 956
rect 1474 913 1493 916
rect 1394 863 1421 866
rect 1394 813 1397 863
rect 1418 853 1421 863
rect 1442 806 1445 846
rect 1450 813 1453 826
rect 1442 803 1453 806
rect 1378 753 1385 756
rect 1314 693 1325 696
rect 1322 636 1325 693
rect 1314 633 1325 636
rect 1306 613 1309 626
rect 1306 533 1309 566
rect 1314 526 1317 633
rect 1322 533 1325 606
rect 1330 573 1333 606
rect 1306 523 1317 526
rect 1330 523 1333 536
rect 1306 413 1309 523
rect 1202 313 1205 326
rect 1194 243 1197 266
rect 1194 166 1197 216
rect 1210 213 1213 246
rect 1202 193 1205 206
rect 1218 203 1221 326
rect 1234 213 1237 326
rect 1274 323 1277 403
rect 1306 386 1309 406
rect 1298 383 1309 386
rect 1234 183 1237 206
rect 1194 163 1213 166
rect 1242 163 1245 216
rect 1250 213 1253 276
rect 1258 203 1261 316
rect 1298 276 1301 383
rect 1298 273 1309 276
rect 1306 253 1309 273
rect 1314 233 1317 366
rect 1322 343 1325 416
rect 1330 333 1333 426
rect 1338 363 1341 616
rect 1346 593 1349 616
rect 1346 543 1365 546
rect 1346 523 1349 543
rect 1354 523 1357 536
rect 1362 533 1365 543
rect 1378 503 1381 753
rect 1418 723 1421 766
rect 1426 703 1429 736
rect 1450 676 1453 803
rect 1474 793 1477 906
rect 1490 786 1493 913
rect 1498 803 1501 856
rect 1482 783 1493 786
rect 1474 733 1477 746
rect 1466 723 1477 726
rect 1450 673 1477 676
rect 1394 523 1397 556
rect 1426 523 1429 616
rect 1458 593 1461 606
rect 1474 553 1477 673
rect 1370 393 1373 406
rect 1394 376 1397 416
rect 1386 373 1397 376
rect 1338 266 1341 336
rect 1346 333 1357 336
rect 1346 273 1349 326
rect 1338 263 1357 266
rect 1266 213 1269 226
rect 1322 193 1325 206
rect 1210 123 1213 163
rect 1266 123 1269 166
rect 1298 133 1301 156
rect 1330 123 1333 216
rect 1338 213 1341 236
rect 1346 196 1349 206
rect 1354 203 1357 263
rect 1362 223 1365 326
rect 1370 323 1373 336
rect 1378 333 1381 346
rect 1386 323 1389 373
rect 1394 323 1397 356
rect 1434 353 1437 536
rect 1442 506 1445 536
rect 1482 523 1485 783
rect 1498 756 1501 796
rect 1506 783 1509 816
rect 1522 813 1525 926
rect 1538 906 1541 953
rect 1562 933 1565 946
rect 1586 923 1589 1016
rect 1594 1013 1597 1103
rect 1602 926 1605 1173
rect 1626 1146 1629 1166
rect 1658 1163 1661 1313
rect 1682 1306 1685 1326
rect 1674 1303 1685 1306
rect 1674 1246 1677 1303
rect 1674 1243 1685 1246
rect 1674 1176 1677 1216
rect 1670 1173 1677 1176
rect 1626 1143 1637 1146
rect 1634 1066 1637 1143
rect 1650 1123 1653 1136
rect 1670 1096 1673 1173
rect 1682 1103 1685 1243
rect 1690 1203 1693 1326
rect 1706 1283 1709 1326
rect 1738 1323 1741 1376
rect 1746 1333 1749 1346
rect 1690 1123 1693 1136
rect 1722 1133 1725 1206
rect 1730 1186 1733 1216
rect 1738 1203 1741 1296
rect 1754 1293 1757 1396
rect 1762 1373 1765 1446
rect 1774 1366 1777 1453
rect 1786 1393 1789 1556
rect 1770 1363 1777 1366
rect 1762 1313 1765 1326
rect 1746 1213 1749 1286
rect 1770 1276 1773 1363
rect 1778 1333 1781 1346
rect 1786 1313 1789 1336
rect 1762 1273 1773 1276
rect 1730 1183 1737 1186
rect 1670 1093 1677 1096
rect 1618 1063 1637 1066
rect 1610 973 1613 1006
rect 1618 966 1621 1063
rect 1626 1003 1629 1056
rect 1674 1046 1677 1093
rect 1666 1043 1677 1046
rect 1634 1013 1645 1016
rect 1618 963 1629 966
rect 1602 923 1613 926
rect 1538 903 1549 906
rect 1530 813 1533 826
rect 1514 773 1517 806
rect 1522 783 1525 806
rect 1498 753 1509 756
rect 1490 723 1493 736
rect 1506 636 1509 753
rect 1530 713 1533 726
rect 1538 723 1541 736
rect 1490 613 1493 636
rect 1498 633 1509 636
rect 1490 506 1493 556
rect 1442 503 1453 506
rect 1450 446 1453 503
rect 1442 443 1453 446
rect 1482 503 1493 506
rect 1362 196 1365 216
rect 1370 203 1373 256
rect 1378 213 1381 296
rect 1346 193 1365 196
rect 1378 193 1381 206
rect 1386 123 1389 216
rect 1402 213 1405 226
rect 1402 123 1405 206
rect 1410 173 1413 216
rect 1418 196 1421 216
rect 1426 203 1429 216
rect 1434 213 1437 236
rect 1442 223 1445 443
rect 1450 413 1453 426
rect 1458 406 1461 416
rect 1450 403 1461 406
rect 1450 323 1453 403
rect 1482 376 1485 503
rect 1482 373 1493 376
rect 1474 333 1477 346
rect 1434 196 1437 206
rect 1418 193 1437 196
rect 1450 123 1453 216
rect 1458 213 1461 236
rect 1466 203 1469 266
rect 1490 233 1493 373
rect 1498 343 1501 633
rect 1506 503 1509 606
rect 1514 546 1517 616
rect 1530 613 1533 626
rect 1522 563 1525 606
rect 1514 543 1533 546
rect 1514 403 1517 526
rect 1522 473 1525 536
rect 1530 533 1533 543
rect 1538 523 1541 556
rect 1546 523 1549 903
rect 1578 733 1581 806
rect 1570 713 1573 726
rect 1586 716 1589 816
rect 1602 813 1605 836
rect 1594 753 1597 806
rect 1610 763 1613 923
rect 1626 876 1629 963
rect 1622 873 1629 876
rect 1622 826 1625 873
rect 1634 833 1637 1013
rect 1642 923 1645 1006
rect 1650 1003 1653 1036
rect 1650 923 1653 936
rect 1618 823 1625 826
rect 1586 713 1597 716
rect 1594 656 1597 713
rect 1594 653 1601 656
rect 1598 576 1601 653
rect 1594 573 1601 576
rect 1594 513 1597 573
rect 1610 523 1613 616
rect 1618 593 1621 823
rect 1634 753 1637 806
rect 1642 803 1645 916
rect 1666 896 1669 1043
rect 1674 1013 1677 1036
rect 1658 893 1669 896
rect 1682 893 1685 936
rect 1690 923 1693 996
rect 1698 933 1701 946
rect 1722 926 1725 1126
rect 1734 1116 1737 1183
rect 1762 1166 1765 1273
rect 1762 1163 1773 1166
rect 1746 1143 1765 1146
rect 1746 1133 1749 1143
rect 1734 1113 1741 1116
rect 1738 1046 1741 1113
rect 1754 1103 1757 1136
rect 1762 1123 1765 1143
rect 1730 1043 1741 1046
rect 1730 1013 1733 1043
rect 1730 1003 1741 1006
rect 1746 1003 1749 1026
rect 1754 1013 1765 1016
rect 1722 923 1733 926
rect 1746 906 1749 986
rect 1770 983 1773 1163
rect 1778 1133 1781 1296
rect 1778 1113 1781 1126
rect 1786 1013 1789 1216
rect 1794 1006 1797 1573
rect 1802 1166 1805 1726
rect 1818 1723 1821 1803
rect 1842 1793 1845 1926
rect 1850 1896 1853 2163
rect 1866 2133 1877 2136
rect 1866 2093 1869 2133
rect 1890 2123 1893 2463
rect 1898 2416 1901 2586
rect 1922 2536 1925 2606
rect 1906 2423 1909 2536
rect 1914 2533 1925 2536
rect 1938 2416 1941 2606
rect 1954 2503 1957 2536
rect 1898 2413 1909 2416
rect 1898 2306 1901 2406
rect 1906 2323 1909 2413
rect 1922 2413 1941 2416
rect 1922 2396 1925 2413
rect 1946 2403 1949 2426
rect 1918 2393 1925 2396
rect 1918 2306 1921 2393
rect 1898 2303 1905 2306
rect 1918 2303 1925 2306
rect 1902 2226 1905 2303
rect 1898 2223 1905 2226
rect 1898 2203 1901 2223
rect 1866 1923 1869 1936
rect 1882 1933 1885 1946
rect 1906 1923 1909 2016
rect 1914 1976 1917 2286
rect 1922 2216 1925 2303
rect 1930 2223 1933 2396
rect 1954 2326 1957 2416
rect 1962 2393 1965 2406
rect 1970 2386 1973 2616
rect 1986 2603 1989 2623
rect 1994 2603 1997 2626
rect 2002 2596 2005 2633
rect 1994 2593 2005 2596
rect 1978 2513 1981 2526
rect 1970 2383 1981 2386
rect 1994 2383 1997 2593
rect 2018 2533 2021 2713
rect 2034 2603 2037 3146
rect 2050 3083 2053 3166
rect 2058 3133 2069 3136
rect 2066 3116 2069 3126
rect 2058 3113 2069 3116
rect 2050 2916 2053 3006
rect 2058 3003 2061 3113
rect 2074 3093 2077 3253
rect 2082 3233 2085 3326
rect 2090 3273 2093 3406
rect 2098 3403 2101 3453
rect 2106 3413 2109 3436
rect 2138 3403 2141 3453
rect 2150 3376 2153 3463
rect 2146 3373 2153 3376
rect 2090 3213 2093 3226
rect 2098 3146 2101 3326
rect 2106 3203 2109 3216
rect 2098 3143 2105 3146
rect 2066 2993 2069 3006
rect 2074 2983 2077 3086
rect 2082 3013 2085 3136
rect 2090 3003 2093 3136
rect 2102 3026 2105 3143
rect 2098 3023 2105 3026
rect 2098 3003 2101 3023
rect 2082 2983 2093 2986
rect 2050 2913 2069 2916
rect 2050 2746 2053 2896
rect 2050 2743 2057 2746
rect 2054 2686 2057 2743
rect 2066 2723 2069 2913
rect 2082 2893 2085 2983
rect 2098 2873 2101 2996
rect 2114 2983 2117 3366
rect 2146 3356 2149 3373
rect 2162 3363 2165 3646
rect 2182 3576 2185 3653
rect 2178 3573 2185 3576
rect 2170 3523 2173 3536
rect 2178 3356 2181 3573
rect 2186 3533 2189 3556
rect 2130 3353 2149 3356
rect 2174 3353 2181 3356
rect 2130 3333 2133 3353
rect 2146 3333 2149 3346
rect 2122 3323 2133 3326
rect 2122 3203 2125 3256
rect 2122 3123 2125 3136
rect 2130 3106 2133 3266
rect 2126 3103 2133 3106
rect 2126 2946 2129 3103
rect 2138 2983 2141 3216
rect 2146 2993 2149 3326
rect 2174 3296 2177 3353
rect 2186 3313 2189 3326
rect 2170 3293 2177 3296
rect 2154 3203 2165 3206
rect 2154 3173 2157 3203
rect 2170 3153 2173 3293
rect 2186 3136 2189 3216
rect 2194 3213 2197 4293
rect 2234 4236 2237 4516
rect 2242 4503 2245 4556
rect 2274 4473 2277 4526
rect 2290 4496 2293 4536
rect 2298 4523 2301 4606
rect 2314 4603 2317 4616
rect 2322 4533 2325 4616
rect 2378 4603 2381 4616
rect 2330 4533 2333 4566
rect 2370 4533 2381 4536
rect 2386 4533 2389 4556
rect 2394 4533 2397 4586
rect 2290 4493 2301 4496
rect 2282 4413 2285 4486
rect 2298 4436 2301 4493
rect 2290 4433 2301 4436
rect 2266 4393 2269 4406
rect 2282 4383 2285 4406
rect 2290 4403 2293 4433
rect 2314 4416 2317 4526
rect 2322 4513 2325 4526
rect 2378 4493 2381 4526
rect 2394 4513 2397 4526
rect 2298 4396 2301 4416
rect 2306 4403 2309 4416
rect 2314 4413 2325 4416
rect 2378 4413 2381 4426
rect 2418 4413 2421 4426
rect 2314 4396 2317 4406
rect 2298 4393 2317 4396
rect 2322 4356 2325 4413
rect 2394 4393 2397 4406
rect 2426 4393 2429 4606
rect 2530 4576 2533 4606
rect 2562 4603 2565 4616
rect 2578 4576 2581 4606
rect 2602 4603 2605 4616
rect 2646 4586 2649 4653
rect 2834 4616 2837 4686
rect 3034 4626 3037 4646
rect 2642 4583 2649 4586
rect 2530 4573 2541 4576
rect 2578 4573 2597 4576
rect 2458 4516 2461 4536
rect 2450 4513 2461 4516
rect 2450 4466 2453 4513
rect 2466 4493 2469 4526
rect 2474 4486 2477 4536
rect 2482 4503 2485 4526
rect 2474 4483 2485 4486
rect 2450 4463 2461 4466
rect 2458 4393 2461 4463
rect 2482 4436 2485 4483
rect 2474 4433 2485 4436
rect 2474 4416 2477 4433
rect 2466 4413 2477 4416
rect 2506 4413 2509 4426
rect 2514 4403 2517 4416
rect 2306 4353 2325 4356
rect 2242 4323 2253 4326
rect 2258 4303 2261 4326
rect 2306 4323 2309 4353
rect 2314 4343 2333 4346
rect 2314 4333 2317 4343
rect 2322 4323 2325 4336
rect 2330 4323 2333 4343
rect 2338 4333 2341 4386
rect 2378 4316 2381 4336
rect 2370 4313 2381 4316
rect 2230 4233 2237 4236
rect 2202 4173 2205 4206
rect 2202 4123 2205 4136
rect 2210 4013 2213 4126
rect 2218 4123 2221 4196
rect 2230 4126 2233 4233
rect 2242 4213 2245 4226
rect 2258 4213 2261 4246
rect 2370 4236 2373 4313
rect 2386 4296 2389 4326
rect 2394 4303 2397 4326
rect 2386 4293 2397 4296
rect 2370 4233 2381 4236
rect 2282 4213 2285 4226
rect 2242 4133 2245 4206
rect 2258 4163 2261 4206
rect 2230 4123 2237 4126
rect 2218 3933 2221 4016
rect 2234 3916 2237 4123
rect 2250 4113 2253 4126
rect 2258 3936 2261 4126
rect 2290 4113 2293 4126
rect 2306 4096 2309 4166
rect 2338 4143 2341 4216
rect 2362 4176 2365 4216
rect 2378 4213 2381 4233
rect 2394 4213 2397 4293
rect 2370 4193 2373 4206
rect 2362 4173 2377 4176
rect 2338 4123 2341 4136
rect 2362 4133 2365 4146
rect 2298 4093 2309 4096
rect 2282 4003 2285 4016
rect 2298 3996 2301 4093
rect 2314 4003 2317 4106
rect 2330 4013 2333 4066
rect 2338 4006 2341 4076
rect 2374 4066 2377 4173
rect 2386 4073 2389 4206
rect 2402 4193 2405 4326
rect 2410 4276 2413 4326
rect 2434 4303 2437 4326
rect 2410 4273 2421 4276
rect 2418 4226 2421 4273
rect 2410 4223 2421 4226
rect 2410 4203 2413 4223
rect 2402 4123 2405 4146
rect 2410 4133 2413 4166
rect 2450 4143 2453 4276
rect 2482 4216 2485 4336
rect 2458 4173 2461 4206
rect 2374 4063 2381 4066
rect 2362 4013 2365 4056
rect 2338 4003 2349 4006
rect 2298 3993 2309 3996
rect 2258 3933 2269 3936
rect 2226 3913 2237 3916
rect 2202 3813 2205 3836
rect 2210 3723 2213 3876
rect 2226 3826 2229 3913
rect 2226 3823 2237 3826
rect 2226 3776 2229 3806
rect 2234 3783 2237 3823
rect 2242 3796 2245 3926
rect 2266 3866 2269 3933
rect 2250 3863 2269 3866
rect 2250 3803 2253 3863
rect 2258 3813 2261 3826
rect 2290 3816 2293 3936
rect 2306 3833 2309 3993
rect 2322 3923 2325 3986
rect 2346 3933 2349 4003
rect 2378 3976 2381 4063
rect 2394 4003 2397 4016
rect 2402 4003 2405 4016
rect 2418 4006 2421 4036
rect 2426 4013 2429 4136
rect 2442 4123 2445 4136
rect 2466 4133 2469 4216
rect 2482 4213 2493 4216
rect 2474 4193 2477 4206
rect 2450 4123 2461 4126
rect 2490 4096 2493 4213
rect 2514 4176 2517 4386
rect 2522 4353 2525 4536
rect 2538 4523 2541 4573
rect 2554 4446 2557 4526
rect 2570 4473 2573 4526
rect 2546 4443 2557 4446
rect 2546 4416 2549 4443
rect 2562 4416 2565 4436
rect 2530 4396 2533 4416
rect 2538 4403 2541 4416
rect 2546 4413 2557 4416
rect 2562 4413 2569 4416
rect 2578 4413 2581 4426
rect 2546 4396 2549 4406
rect 2530 4393 2549 4396
rect 2554 4363 2557 4413
rect 2530 4323 2533 4336
rect 2538 4333 2549 4336
rect 2554 4333 2557 4356
rect 2538 4213 2541 4326
rect 2546 4323 2549 4333
rect 2566 4326 2569 4413
rect 2594 4383 2597 4573
rect 2642 4456 2645 4583
rect 2658 4533 2661 4616
rect 2682 4576 2685 4606
rect 2706 4603 2709 4616
rect 2722 4593 2725 4606
rect 2746 4603 2749 4616
rect 2682 4573 2693 4576
rect 2634 4453 2645 4456
rect 2618 4413 2621 4426
rect 2634 4396 2637 4453
rect 2666 4413 2677 4416
rect 2634 4393 2645 4396
rect 2562 4323 2569 4326
rect 2578 4323 2589 4326
rect 2562 4256 2565 4323
rect 2554 4253 2565 4256
rect 2530 4176 2533 4196
rect 2514 4173 2533 4176
rect 2554 4176 2557 4253
rect 2594 4213 2597 4336
rect 2602 4333 2605 4366
rect 2610 4323 2613 4376
rect 2642 4373 2645 4393
rect 2674 4383 2677 4413
rect 2602 4213 2605 4246
rect 2554 4173 2565 4176
rect 2530 4133 2533 4173
rect 2562 4136 2565 4173
rect 2594 4143 2613 4146
rect 2562 4133 2573 4136
rect 2594 4133 2597 4143
rect 2506 4113 2509 4126
rect 2546 4113 2549 4126
rect 2482 4093 2493 4096
rect 2482 4073 2485 4093
rect 2554 4083 2557 4126
rect 2418 4003 2429 4006
rect 2434 4003 2437 4056
rect 2530 4046 2533 4076
rect 2522 4043 2533 4046
rect 2466 4003 2469 4016
rect 2474 4013 2485 4016
rect 2506 4003 2509 4016
rect 2522 3996 2525 4043
rect 2554 4003 2557 4036
rect 2370 3973 2381 3976
rect 2354 3923 2365 3926
rect 2370 3846 2373 3973
rect 2378 3886 2381 3946
rect 2386 3906 2389 3996
rect 2522 3993 2533 3996
rect 2394 3923 2397 3936
rect 2386 3903 2397 3906
rect 2442 3903 2445 3926
rect 2450 3923 2453 3946
rect 2378 3883 2385 3886
rect 2354 3843 2373 3846
rect 2266 3803 2269 3816
rect 2242 3793 2261 3796
rect 2226 3773 2237 3776
rect 2202 3583 2205 3616
rect 2210 3613 2213 3696
rect 2226 3676 2229 3746
rect 2234 3723 2237 3773
rect 2242 3733 2245 3766
rect 2242 3723 2253 3726
rect 2218 3673 2229 3676
rect 2210 3593 2213 3606
rect 2218 3576 2221 3673
rect 2226 3593 2229 3616
rect 2242 3613 2245 3723
rect 2258 3636 2261 3793
rect 2282 3643 2285 3816
rect 2290 3813 2301 3816
rect 2298 3766 2301 3813
rect 2290 3763 2301 3766
rect 2290 3743 2293 3763
rect 2314 3733 2317 3766
rect 2258 3633 2265 3636
rect 2250 3613 2253 3626
rect 2214 3573 2221 3576
rect 2214 3526 2217 3573
rect 2226 3533 2229 3566
rect 2234 3533 2237 3606
rect 2262 3586 2265 3633
rect 2258 3583 2265 3586
rect 2258 3563 2261 3583
rect 2202 3513 2205 3526
rect 2214 3523 2221 3526
rect 2218 3433 2221 3523
rect 2258 3466 2261 3486
rect 2254 3463 2261 3466
rect 2210 3333 2237 3336
rect 2210 3213 2213 3333
rect 2226 3226 2229 3326
rect 2234 3313 2237 3326
rect 2218 3223 2229 3226
rect 2194 3183 2197 3206
rect 2218 3143 2221 3223
rect 2226 3203 2229 3216
rect 2242 3166 2245 3426
rect 2234 3163 2245 3166
rect 2154 3123 2157 3136
rect 2154 3013 2157 3026
rect 2126 2943 2133 2946
rect 2130 2926 2133 2943
rect 2138 2933 2141 2946
rect 2146 2933 2149 2966
rect 2082 2773 2085 2836
rect 2122 2813 2125 2926
rect 2130 2923 2137 2926
rect 2098 2783 2101 2806
rect 2050 2683 2057 2686
rect 2042 2603 2045 2616
rect 2050 2596 2053 2683
rect 2074 2663 2077 2726
rect 2082 2703 2085 2736
rect 2098 2636 2101 2766
rect 2134 2746 2137 2923
rect 2134 2743 2141 2746
rect 2122 2723 2133 2726
rect 2122 2706 2125 2723
rect 2138 2716 2141 2743
rect 2114 2703 2125 2706
rect 2130 2713 2141 2716
rect 2114 2646 2117 2703
rect 2114 2643 2125 2646
rect 2034 2593 2053 2596
rect 2090 2633 2101 2636
rect 2034 2526 2037 2593
rect 2090 2556 2093 2633
rect 2106 2566 2109 2626
rect 2114 2593 2117 2606
rect 2122 2603 2125 2643
rect 2130 2586 2133 2713
rect 2126 2583 2133 2586
rect 2106 2563 2117 2566
rect 2090 2553 2101 2556
rect 2018 2513 2021 2526
rect 2026 2523 2037 2526
rect 2026 2413 2029 2523
rect 2074 2516 2077 2536
rect 2070 2513 2077 2516
rect 1946 2323 1957 2326
rect 1922 2213 1933 2216
rect 1938 2203 1941 2236
rect 1946 2213 1949 2323
rect 1978 2286 1981 2383
rect 1970 2283 1981 2286
rect 1954 2186 1957 2206
rect 1946 2183 1957 2186
rect 1946 2056 1949 2183
rect 1962 2133 1965 2226
rect 1970 2196 1973 2283
rect 1994 2213 1997 2326
rect 1970 2193 1981 2196
rect 1978 2146 1981 2193
rect 1970 2143 1981 2146
rect 1946 2053 1957 2056
rect 1930 1996 1933 2006
rect 1938 2003 1941 2036
rect 1946 1996 1949 2016
rect 1954 2003 1957 2053
rect 1970 2013 1973 2143
rect 1930 1993 1949 1996
rect 1914 1973 1925 1976
rect 1922 1916 1925 1973
rect 1914 1913 1925 1916
rect 1850 1893 1861 1896
rect 1858 1836 1861 1893
rect 1882 1846 1885 1866
rect 1882 1843 1893 1846
rect 1858 1833 1877 1836
rect 1858 1803 1861 1816
rect 1842 1776 1845 1786
rect 1834 1773 1845 1776
rect 1834 1653 1837 1773
rect 1866 1756 1869 1796
rect 1858 1753 1869 1756
rect 1858 1666 1861 1753
rect 1874 1673 1877 1833
rect 1890 1786 1893 1843
rect 1882 1783 1893 1786
rect 1914 1783 1917 1913
rect 1954 1906 1957 1926
rect 1962 1923 1965 2006
rect 2018 1976 2021 2386
rect 2034 2333 2037 2366
rect 2042 2273 2045 2476
rect 2050 2376 2053 2456
rect 2058 2413 2061 2506
rect 2070 2376 2073 2513
rect 2082 2403 2085 2526
rect 2090 2403 2093 2416
rect 2050 2373 2057 2376
rect 2070 2373 2077 2376
rect 2054 2226 2057 2373
rect 2074 2356 2077 2373
rect 2074 2353 2085 2356
rect 2054 2223 2061 2226
rect 2050 2123 2053 2206
rect 2058 2106 2061 2223
rect 2050 2103 2061 2106
rect 2050 2056 2053 2103
rect 2050 2053 2061 2056
rect 2058 2033 2061 2053
rect 1970 1923 1973 1976
rect 2018 1973 2029 1976
rect 2018 1943 2021 1973
rect 2034 1906 2037 1926
rect 2050 1923 2053 2016
rect 1950 1903 1957 1906
rect 2026 1903 2037 1906
rect 1950 1836 1953 1903
rect 1950 1833 1957 1836
rect 1858 1663 1869 1666
rect 1834 1516 1837 1526
rect 1842 1523 1845 1616
rect 1850 1516 1853 1526
rect 1866 1516 1869 1663
rect 1874 1533 1877 1546
rect 1834 1513 1853 1516
rect 1858 1513 1869 1516
rect 1858 1496 1861 1513
rect 1850 1493 1861 1496
rect 1850 1406 1853 1493
rect 1866 1413 1869 1506
rect 1882 1456 1885 1783
rect 1890 1723 1901 1726
rect 1906 1723 1909 1766
rect 1914 1733 1917 1776
rect 1890 1543 1893 1606
rect 1890 1523 1893 1536
rect 1898 1533 1901 1723
rect 1922 1706 1925 1816
rect 1930 1783 1933 1806
rect 1938 1803 1941 1826
rect 1954 1733 1957 1833
rect 1962 1813 1965 1886
rect 2026 1836 2029 1903
rect 2050 1896 2053 1916
rect 2046 1893 2053 1896
rect 2026 1833 2037 1836
rect 2002 1803 2005 1816
rect 2034 1813 2037 1833
rect 1954 1713 1957 1726
rect 1914 1703 1925 1706
rect 1914 1636 1917 1703
rect 1914 1633 1925 1636
rect 1922 1613 1925 1633
rect 1930 1603 1933 1706
rect 1938 1613 1941 1696
rect 1898 1523 1909 1526
rect 1914 1516 1917 1546
rect 1922 1523 1925 1566
rect 1906 1513 1917 1516
rect 1906 1496 1909 1513
rect 1902 1493 1909 1496
rect 1882 1453 1893 1456
rect 1818 1393 1821 1406
rect 1850 1403 1869 1406
rect 1818 1313 1821 1326
rect 1826 1323 1829 1346
rect 1858 1313 1861 1326
rect 1802 1163 1813 1166
rect 1810 1146 1813 1163
rect 1810 1143 1817 1146
rect 1814 1076 1817 1143
rect 1810 1073 1817 1076
rect 1810 1056 1813 1073
rect 1802 1053 1813 1056
rect 1802 1013 1805 1053
rect 1826 1006 1829 1136
rect 1834 1106 1837 1136
rect 1842 1123 1845 1216
rect 1850 1123 1853 1136
rect 1834 1103 1841 1106
rect 1838 1036 1841 1103
rect 1834 1033 1841 1036
rect 1834 1013 1837 1033
rect 1850 1013 1853 1096
rect 1866 1026 1869 1403
rect 1890 1376 1893 1453
rect 1902 1436 1905 1493
rect 1902 1433 1909 1436
rect 1906 1413 1909 1433
rect 1914 1413 1917 1506
rect 1930 1503 1933 1536
rect 1946 1533 1949 1606
rect 1946 1403 1949 1526
rect 1954 1513 1957 1616
rect 1954 1396 1957 1496
rect 1962 1413 1965 1526
rect 1970 1493 1973 1726
rect 1978 1723 1981 1756
rect 2002 1716 2005 1736
rect 1994 1713 2005 1716
rect 1994 1666 1997 1713
rect 2010 1696 2013 1746
rect 2034 1733 2037 1806
rect 2046 1796 2049 1893
rect 2058 1803 2061 1936
rect 2066 1913 2069 2346
rect 2082 2236 2085 2353
rect 2098 2306 2101 2553
rect 2114 2466 2117 2563
rect 2126 2526 2129 2583
rect 2138 2533 2141 2656
rect 2126 2523 2133 2526
rect 2106 2463 2117 2466
rect 2106 2386 2109 2463
rect 2114 2403 2117 2446
rect 2106 2383 2113 2386
rect 2074 2233 2085 2236
rect 2094 2303 2101 2306
rect 2094 2236 2097 2303
rect 2110 2296 2113 2383
rect 2106 2293 2113 2296
rect 2094 2233 2101 2236
rect 2074 2093 2077 2233
rect 2090 2203 2093 2216
rect 2082 1976 2085 2146
rect 2074 1973 2085 1976
rect 2074 1896 2077 1973
rect 2070 1893 2077 1896
rect 2070 1826 2073 1893
rect 2070 1823 2077 1826
rect 2046 1793 2053 1796
rect 2066 1793 2069 1806
rect 2074 1803 2077 1823
rect 2026 1713 2029 1726
rect 2042 1723 2045 1776
rect 2010 1693 2021 1696
rect 1994 1663 2005 1666
rect 1994 1603 1997 1646
rect 2002 1546 2005 1663
rect 2018 1626 2021 1693
rect 2010 1623 2021 1626
rect 2010 1603 2013 1623
rect 2034 1596 2037 1616
rect 2026 1593 2037 1596
rect 2002 1543 2013 1546
rect 1986 1503 1989 1526
rect 1994 1473 1997 1536
rect 2010 1466 2013 1543
rect 2002 1463 2013 1466
rect 2002 1443 2005 1463
rect 2026 1456 2029 1593
rect 2042 1576 2045 1676
rect 2038 1573 2045 1576
rect 2038 1476 2041 1573
rect 2038 1473 2045 1476
rect 2026 1453 2037 1456
rect 1970 1413 1973 1426
rect 1882 1373 1893 1376
rect 1882 1356 1885 1373
rect 1878 1353 1885 1356
rect 1878 1296 1881 1353
rect 1906 1333 1909 1396
rect 1946 1393 1957 1396
rect 1930 1323 1933 1336
rect 1946 1306 1949 1393
rect 1938 1303 1949 1306
rect 1878 1293 1885 1296
rect 1882 1146 1885 1293
rect 1938 1226 1941 1303
rect 1938 1223 1949 1226
rect 1890 1196 1893 1216
rect 1890 1193 1901 1196
rect 1946 1193 1949 1223
rect 1954 1196 1957 1216
rect 1962 1203 1965 1316
rect 1970 1213 1973 1406
rect 1994 1403 1997 1436
rect 2010 1413 2013 1426
rect 1978 1346 1981 1366
rect 1978 1343 1985 1346
rect 1982 1206 1985 1343
rect 1970 1196 1973 1206
rect 1954 1193 1973 1196
rect 1978 1203 1985 1206
rect 1878 1143 1885 1146
rect 1878 1046 1881 1143
rect 1898 1136 1901 1193
rect 1978 1186 1981 1203
rect 1970 1183 1981 1186
rect 1890 1133 1901 1136
rect 1890 1046 1893 1133
rect 1946 1123 1949 1136
rect 1970 1076 1973 1183
rect 1986 1133 1989 1146
rect 1994 1116 1997 1396
rect 2002 1366 2005 1386
rect 2002 1363 2009 1366
rect 2018 1363 2021 1436
rect 2026 1403 2029 1416
rect 2034 1383 2037 1453
rect 2006 1236 2009 1363
rect 1962 1073 1973 1076
rect 1990 1113 1997 1116
rect 2002 1233 2009 1236
rect 1878 1043 1885 1046
rect 1890 1043 1901 1046
rect 1866 1023 1873 1026
rect 1762 943 1781 946
rect 1762 933 1765 943
rect 1754 913 1757 926
rect 1762 906 1765 926
rect 1746 903 1765 906
rect 1770 893 1773 936
rect 1778 923 1781 943
rect 1786 933 1789 1006
rect 1794 1003 1813 1006
rect 1826 1003 1845 1006
rect 1858 1003 1861 1016
rect 1786 923 1797 926
rect 1802 923 1805 946
rect 1658 776 1661 893
rect 1666 813 1669 826
rect 1698 816 1701 876
rect 1786 843 1789 923
rect 1810 853 1813 1003
rect 1834 913 1837 926
rect 1842 893 1845 1003
rect 1858 976 1861 996
rect 1870 976 1873 1023
rect 1882 993 1885 1043
rect 1854 973 1861 976
rect 1866 973 1873 976
rect 1854 896 1857 973
rect 1866 953 1869 973
rect 1898 956 1901 1043
rect 1938 1013 1941 1026
rect 1962 976 1965 1073
rect 1978 1013 1981 1026
rect 1954 973 1965 976
rect 1882 913 1885 956
rect 1898 953 1909 956
rect 1906 906 1909 953
rect 1930 923 1933 936
rect 1954 933 1957 973
rect 1898 903 1909 906
rect 1854 893 1861 896
rect 1674 783 1677 806
rect 1690 803 1693 816
rect 1698 813 1709 816
rect 1658 773 1685 776
rect 1658 733 1661 766
rect 1682 756 1685 773
rect 1682 753 1689 756
rect 1686 696 1689 753
rect 1682 693 1689 696
rect 1642 593 1645 606
rect 1658 603 1661 616
rect 1666 603 1677 606
rect 1682 603 1685 693
rect 1698 616 1701 813
rect 1714 776 1717 816
rect 1706 773 1717 776
rect 1722 776 1725 836
rect 1778 813 1781 836
rect 1730 793 1733 806
rect 1722 773 1729 776
rect 1706 723 1709 773
rect 1726 686 1729 773
rect 1738 723 1741 756
rect 1762 706 1765 726
rect 1754 703 1765 706
rect 1726 683 1741 686
rect 1694 613 1701 616
rect 1642 436 1645 536
rect 1650 523 1653 536
rect 1658 533 1661 546
rect 1666 513 1669 603
rect 1694 556 1697 613
rect 1694 553 1701 556
rect 1642 433 1653 436
rect 1546 393 1549 416
rect 1602 413 1605 426
rect 1642 413 1645 426
rect 1626 383 1629 406
rect 1498 333 1509 336
rect 1514 333 1533 336
rect 1498 293 1501 333
rect 1498 193 1501 216
rect 1506 213 1509 326
rect 1514 323 1517 333
rect 1522 286 1525 326
rect 1530 323 1533 333
rect 1586 306 1589 326
rect 1514 283 1525 286
rect 1578 303 1589 306
rect 1514 213 1517 283
rect 1578 236 1581 303
rect 1610 256 1613 346
rect 1626 293 1629 336
rect 1642 333 1645 406
rect 1650 393 1653 433
rect 1658 386 1661 426
rect 1666 403 1669 476
rect 1682 473 1685 536
rect 1690 426 1693 536
rect 1674 423 1693 426
rect 1698 423 1701 553
rect 1706 523 1709 606
rect 1714 593 1717 606
rect 1730 603 1733 616
rect 1738 596 1741 683
rect 1754 646 1757 703
rect 1754 643 1765 646
rect 1746 603 1749 626
rect 1738 593 1749 596
rect 1714 513 1717 526
rect 1722 506 1725 536
rect 1738 533 1741 586
rect 1746 523 1749 593
rect 1754 586 1757 616
rect 1762 603 1765 643
rect 1770 613 1773 806
rect 1786 803 1789 826
rect 1802 816 1805 846
rect 1802 813 1813 816
rect 1818 813 1821 826
rect 1802 793 1805 806
rect 1810 776 1813 813
rect 1802 773 1813 776
rect 1786 613 1789 706
rect 1802 636 1805 773
rect 1826 766 1829 886
rect 1858 856 1861 893
rect 1834 813 1837 856
rect 1854 853 1861 856
rect 1834 773 1837 806
rect 1842 803 1845 816
rect 1854 796 1857 853
rect 1874 813 1877 836
rect 1854 793 1861 796
rect 1898 793 1901 903
rect 1858 776 1861 793
rect 1858 773 1869 776
rect 1818 763 1829 766
rect 1802 633 1813 636
rect 1810 613 1813 633
rect 1754 583 1773 586
rect 1650 383 1661 386
rect 1674 386 1677 423
rect 1682 396 1685 406
rect 1690 403 1693 416
rect 1698 396 1701 416
rect 1682 393 1701 396
rect 1706 393 1709 406
rect 1674 383 1685 386
rect 1634 313 1637 326
rect 1602 253 1613 256
rect 1578 233 1589 236
rect 1482 133 1485 146
rect 1506 123 1509 206
rect 1514 193 1517 206
rect 1570 123 1573 216
rect 1578 203 1581 216
rect 1586 213 1589 233
rect 1602 133 1605 253
rect 1650 213 1653 383
rect 1666 223 1669 336
rect 1674 323 1677 336
rect 1682 213 1685 383
rect 1690 303 1693 336
rect 1698 273 1701 326
rect 1634 123 1637 206
rect 1650 203 1661 206
rect 1674 183 1677 206
rect 1682 193 1685 206
rect 1714 203 1717 506
rect 1722 503 1733 506
rect 1730 456 1733 503
rect 1722 453 1733 456
rect 1722 433 1725 453
rect 1722 323 1725 336
rect 1746 333 1749 346
rect 1746 313 1749 326
rect 1754 296 1757 416
rect 1762 413 1765 536
rect 1770 513 1773 583
rect 1778 516 1781 606
rect 1818 603 1821 763
rect 1826 723 1829 736
rect 1858 713 1861 726
rect 1786 543 1805 546
rect 1786 523 1789 543
rect 1794 516 1797 536
rect 1802 533 1805 543
rect 1778 513 1797 516
rect 1794 413 1797 513
rect 1802 493 1805 526
rect 1818 413 1821 526
rect 1826 513 1829 616
rect 1834 533 1837 626
rect 1842 543 1861 546
rect 1842 523 1845 543
rect 1850 503 1853 536
rect 1858 533 1861 543
rect 1858 513 1861 526
rect 1858 413 1861 496
rect 1866 453 1869 773
rect 1874 733 1877 766
rect 1882 733 1893 736
rect 1922 726 1925 916
rect 1938 913 1941 926
rect 1938 813 1941 826
rect 1938 763 1941 806
rect 1946 803 1949 836
rect 1954 813 1957 926
rect 1978 913 1981 926
rect 1990 896 1993 1113
rect 2002 903 2005 1233
rect 2010 1106 2013 1216
rect 2034 1213 2037 1326
rect 2042 1223 2045 1473
rect 2050 1373 2053 1793
rect 2058 1626 2061 1706
rect 2058 1623 2065 1626
rect 2062 1556 2065 1623
rect 2074 1603 2077 1626
rect 2058 1553 2065 1556
rect 2058 1516 2061 1553
rect 2082 1546 2085 1906
rect 2090 1743 2093 2176
rect 2098 2146 2101 2233
rect 2106 2166 2109 2293
rect 2122 2213 2125 2326
rect 2130 2306 2133 2523
rect 2146 2456 2149 2876
rect 2154 2856 2157 3006
rect 2162 2963 2165 3056
rect 2170 3013 2173 3136
rect 2186 3133 2193 3136
rect 2162 2923 2165 2946
rect 2170 2866 2173 3006
rect 2178 2963 2181 3126
rect 2190 3046 2193 3133
rect 2186 3043 2193 3046
rect 2186 3023 2189 3043
rect 2178 2876 2181 2926
rect 2186 2923 2189 3006
rect 2178 2873 2189 2876
rect 2170 2863 2181 2866
rect 2154 2853 2165 2856
rect 2154 2523 2157 2736
rect 2142 2453 2149 2456
rect 2162 2453 2165 2853
rect 2178 2813 2181 2863
rect 2170 2706 2173 2786
rect 2186 2723 2189 2873
rect 2194 2763 2197 2986
rect 2202 2933 2205 3126
rect 2226 3116 2229 3136
rect 2218 3113 2229 3116
rect 2218 3036 2221 3113
rect 2234 3046 2237 3163
rect 2242 3133 2245 3156
rect 2254 3146 2257 3463
rect 2274 3436 2277 3636
rect 2314 3606 2317 3726
rect 2322 3723 2325 3826
rect 2354 3746 2357 3843
rect 2382 3826 2385 3883
rect 2378 3823 2385 3826
rect 2354 3743 2365 3746
rect 2338 3613 2341 3726
rect 2362 3673 2365 3743
rect 2370 3733 2373 3816
rect 2378 3803 2381 3823
rect 2394 3766 2397 3903
rect 2426 3856 2429 3876
rect 2482 3863 2485 3956
rect 2498 3933 2501 3966
rect 2530 3933 2533 3993
rect 2498 3903 2501 3926
rect 2554 3923 2557 3996
rect 2426 3853 2433 3856
rect 2386 3763 2397 3766
rect 2386 3746 2389 3763
rect 2378 3723 2381 3746
rect 2386 3743 2397 3746
rect 2354 3613 2365 3616
rect 2290 3593 2293 3606
rect 2314 3603 2325 3606
rect 2314 3533 2317 3556
rect 2266 3433 2277 3436
rect 2266 3196 2269 3433
rect 2322 3426 2325 3603
rect 2346 3533 2349 3606
rect 2314 3423 2325 3426
rect 2282 3343 2285 3406
rect 2314 3356 2317 3423
rect 2330 3383 2333 3416
rect 2346 3403 2349 3526
rect 2370 3513 2373 3696
rect 2386 3626 2389 3736
rect 2394 3656 2397 3743
rect 2402 3733 2405 3746
rect 2410 3673 2413 3736
rect 2418 3656 2421 3776
rect 2430 3756 2433 3853
rect 2426 3753 2433 3756
rect 2426 3723 2429 3753
rect 2442 3723 2445 3816
rect 2426 3686 2429 3706
rect 2458 3703 2461 3726
rect 2426 3683 2437 3686
rect 2394 3653 2405 3656
rect 2378 3623 2389 3626
rect 2378 3563 2381 3623
rect 2386 3603 2389 3616
rect 2386 3543 2389 3586
rect 2402 3576 2405 3653
rect 2394 3573 2405 3576
rect 2414 3653 2421 3656
rect 2394 3526 2397 3573
rect 2414 3546 2417 3653
rect 2434 3636 2437 3683
rect 2474 3676 2477 3836
rect 2490 3733 2493 3816
rect 2530 3813 2533 3896
rect 2506 3733 2509 3806
rect 2538 3796 2541 3816
rect 2546 3803 2549 3816
rect 2554 3796 2557 3806
rect 2538 3793 2557 3796
rect 2522 3726 2525 3746
rect 2514 3706 2517 3726
rect 2522 3723 2533 3726
rect 2562 3723 2565 3906
rect 2426 3633 2437 3636
rect 2458 3673 2477 3676
rect 2506 3703 2517 3706
rect 2414 3543 2421 3546
rect 2386 3523 2397 3526
rect 2386 3456 2389 3523
rect 2386 3453 2393 3456
rect 2370 3396 2373 3416
rect 2378 3413 2381 3436
rect 2370 3393 2377 3396
rect 2282 3316 2285 3336
rect 2278 3313 2285 3316
rect 2278 3246 2281 3313
rect 2278 3243 2285 3246
rect 2274 3203 2277 3226
rect 2266 3193 2277 3196
rect 2254 3143 2261 3146
rect 2250 3073 2253 3126
rect 2258 3056 2261 3143
rect 2266 3133 2269 3146
rect 2254 3053 2261 3056
rect 2234 3043 2245 3046
rect 2218 3033 2229 3036
rect 2218 2933 2221 3016
rect 2226 3003 2229 3033
rect 2226 2926 2229 2996
rect 2242 2976 2245 3043
rect 2218 2923 2229 2926
rect 2234 2973 2245 2976
rect 2254 2976 2257 3053
rect 2266 3013 2269 3066
rect 2274 2976 2277 3193
rect 2282 3166 2285 3243
rect 2290 3183 2293 3336
rect 2282 3163 2289 3166
rect 2286 3016 2289 3163
rect 2282 3013 2289 3016
rect 2282 2993 2285 3013
rect 2254 2973 2261 2976
rect 2274 2973 2281 2976
rect 2202 2746 2205 2896
rect 2210 2766 2213 2806
rect 2218 2786 2221 2923
rect 2234 2893 2237 2973
rect 2234 2803 2237 2886
rect 2258 2786 2261 2973
rect 2266 2923 2269 2966
rect 2278 2916 2281 2973
rect 2298 2963 2301 3356
rect 2314 3353 2325 3356
rect 2322 3333 2325 3353
rect 2306 3243 2309 3326
rect 2314 3323 2325 3326
rect 2306 3213 2309 3236
rect 2314 3223 2317 3323
rect 2330 3313 2333 3336
rect 2346 3316 2349 3336
rect 2338 3313 2349 3316
rect 2314 3063 2317 3216
rect 2322 3183 2325 3216
rect 2338 3213 2341 3313
rect 2330 3203 2341 3206
rect 2338 3166 2341 3203
rect 2330 3163 2341 3166
rect 2330 3066 2333 3163
rect 2346 3146 2349 3226
rect 2354 3186 2357 3326
rect 2362 3323 2365 3386
rect 2374 3336 2377 3393
rect 2390 3366 2393 3453
rect 2402 3433 2405 3486
rect 2402 3373 2405 3426
rect 2390 3363 2397 3366
rect 2370 3333 2377 3336
rect 2394 3336 2397 3363
rect 2410 3353 2413 3526
rect 2394 3333 2401 3336
rect 2370 3226 2373 3333
rect 2386 3296 2389 3326
rect 2362 3223 2373 3226
rect 2382 3293 2389 3296
rect 2382 3226 2385 3293
rect 2398 3286 2401 3333
rect 2394 3283 2401 3286
rect 2382 3223 2389 3226
rect 2362 3203 2365 3223
rect 2354 3183 2361 3186
rect 2342 3143 2349 3146
rect 2342 3086 2345 3143
rect 2358 3136 2361 3183
rect 2354 3133 2361 3136
rect 2342 3083 2349 3086
rect 2330 3063 2341 3066
rect 2322 3013 2325 3046
rect 2278 2913 2285 2916
rect 2282 2856 2285 2913
rect 2306 2886 2309 2986
rect 2314 2973 2317 3006
rect 2298 2883 2309 2886
rect 2298 2866 2301 2883
rect 2298 2863 2305 2866
rect 2278 2853 2285 2856
rect 2218 2783 2229 2786
rect 2210 2763 2217 2766
rect 2198 2743 2205 2746
rect 2170 2703 2181 2706
rect 2178 2576 2181 2703
rect 2198 2686 2201 2743
rect 2214 2696 2217 2763
rect 2214 2693 2221 2696
rect 2198 2683 2205 2686
rect 2202 2626 2205 2683
rect 2170 2573 2181 2576
rect 2194 2623 2205 2626
rect 2194 2576 2197 2623
rect 2194 2573 2201 2576
rect 2170 2553 2173 2573
rect 2198 2516 2201 2573
rect 2210 2523 2213 2616
rect 2218 2613 2221 2693
rect 2226 2606 2229 2783
rect 2254 2783 2261 2786
rect 2234 2613 2237 2736
rect 2242 2686 2245 2726
rect 2254 2706 2257 2783
rect 2266 2733 2269 2816
rect 2278 2776 2281 2853
rect 2302 2776 2305 2863
rect 2278 2773 2285 2776
rect 2254 2703 2261 2706
rect 2242 2683 2253 2686
rect 2250 2613 2253 2683
rect 2218 2603 2229 2606
rect 2198 2513 2205 2516
rect 2142 2356 2145 2453
rect 2154 2413 2157 2446
rect 2202 2416 2205 2513
rect 2218 2486 2221 2603
rect 2258 2553 2261 2703
rect 2266 2643 2269 2706
rect 2282 2626 2285 2773
rect 2298 2773 2305 2776
rect 2298 2756 2301 2773
rect 2294 2753 2301 2756
rect 2294 2646 2297 2753
rect 2314 2746 2317 2816
rect 2322 2786 2325 2966
rect 2330 2903 2333 2976
rect 2330 2803 2333 2816
rect 2338 2803 2341 3063
rect 2346 3046 2349 3083
rect 2354 3063 2357 3133
rect 2346 3043 2357 3046
rect 2354 2946 2357 3043
rect 2370 3026 2373 3146
rect 2378 3093 2381 3206
rect 2386 3183 2389 3223
rect 2366 3023 2373 3026
rect 2366 2966 2369 3023
rect 2366 2963 2373 2966
rect 2346 2943 2357 2946
rect 2346 2906 2349 2943
rect 2370 2933 2373 2963
rect 2362 2923 2373 2926
rect 2378 2923 2381 3016
rect 2386 3013 2389 3136
rect 2394 3003 2397 3283
rect 2402 3166 2405 3216
rect 2410 3203 2413 3336
rect 2418 3203 2421 3543
rect 2426 3213 2429 3633
rect 2434 3523 2437 3616
rect 2458 3533 2461 3673
rect 2506 3626 2509 3703
rect 2530 3656 2533 3723
rect 2570 3706 2573 4133
rect 2602 4113 2605 4136
rect 2610 4123 2613 4143
rect 2618 4123 2621 4146
rect 2626 4133 2629 4356
rect 2650 4343 2669 4346
rect 2650 4323 2653 4343
rect 2658 4323 2661 4336
rect 2666 4333 2669 4343
rect 2634 4196 2637 4216
rect 2642 4203 2645 4246
rect 2650 4196 2653 4206
rect 2634 4193 2653 4196
rect 2658 4146 2661 4216
rect 2674 4213 2677 4366
rect 2682 4353 2685 4536
rect 2690 4523 2693 4573
rect 2714 4533 2717 4546
rect 2778 4533 2781 4556
rect 2802 4553 2805 4616
rect 2834 4613 2853 4616
rect 2810 4583 2813 4606
rect 2794 4543 2805 4546
rect 2690 4413 2693 4436
rect 2714 4396 2717 4416
rect 2722 4403 2725 4436
rect 2730 4396 2733 4406
rect 2714 4393 2733 4396
rect 2738 4363 2741 4526
rect 2826 4463 2829 4536
rect 2834 4523 2837 4536
rect 2842 4483 2845 4536
rect 2850 4523 2853 4606
rect 2858 4603 2861 4626
rect 2866 4593 2869 4606
rect 2858 4436 2861 4536
rect 2874 4523 2877 4616
rect 2898 4606 2901 4626
rect 2890 4533 2893 4606
rect 2898 4603 2909 4606
rect 2906 4546 2909 4603
rect 2922 4593 2925 4626
rect 3026 4623 3037 4626
rect 2898 4543 2909 4546
rect 2898 4516 2901 4543
rect 2890 4513 2901 4516
rect 2890 4446 2893 4513
rect 2890 4443 2901 4446
rect 2842 4433 2861 4436
rect 2746 4413 2749 4426
rect 2786 4413 2789 4426
rect 2834 4406 2837 4426
rect 2842 4413 2845 4433
rect 2866 4426 2869 4436
rect 2866 4423 2877 4426
rect 2706 4323 2709 4336
rect 2706 4213 2709 4226
rect 2722 4156 2725 4356
rect 2762 4353 2765 4406
rect 2834 4403 2845 4406
rect 2746 4323 2749 4336
rect 2802 4326 2805 4396
rect 2794 4323 2805 4326
rect 2746 4213 2749 4226
rect 2802 4213 2805 4246
rect 2810 4233 2813 4346
rect 2834 4333 2837 4366
rect 2842 4323 2845 4403
rect 2850 4393 2853 4406
rect 2850 4303 2853 4336
rect 2738 4176 2741 4196
rect 2650 4143 2661 4146
rect 2706 4153 2725 4156
rect 2730 4173 2741 4176
rect 2626 4056 2629 4116
rect 2578 3976 2581 4006
rect 2594 3986 2597 4056
rect 2622 4053 2629 4056
rect 2602 4003 2605 4016
rect 2594 3983 2601 3986
rect 2578 3973 2589 3976
rect 2578 3906 2581 3946
rect 2586 3923 2589 3973
rect 2598 3906 2601 3983
rect 2610 3933 2613 4016
rect 2622 3996 2625 4053
rect 2650 4046 2653 4143
rect 2658 4063 2661 4126
rect 2666 4113 2669 4136
rect 2674 4116 2677 4126
rect 2682 4123 2685 4136
rect 2690 4116 2693 4136
rect 2698 4123 2701 4136
rect 2674 4113 2693 4116
rect 2650 4043 2657 4046
rect 2642 4003 2645 4016
rect 2654 3996 2657 4043
rect 2706 4036 2709 4153
rect 2714 4113 2717 4126
rect 2622 3993 2629 3996
rect 2578 3903 2585 3906
rect 2582 3816 2585 3903
rect 2594 3903 2601 3906
rect 2610 3903 2613 3926
rect 2618 3923 2621 3976
rect 2626 3933 2629 3993
rect 2650 3993 2657 3996
rect 2690 4033 2709 4036
rect 2650 3903 2653 3993
rect 2690 3976 2693 4033
rect 2690 3973 2701 3976
rect 2658 3943 2677 3946
rect 2658 3923 2661 3943
rect 2666 3923 2669 3936
rect 2674 3933 2677 3943
rect 2674 3903 2677 3926
rect 2594 3823 2597 3903
rect 2698 3896 2701 3973
rect 2730 3936 2733 4173
rect 2754 4113 2757 4126
rect 2690 3893 2701 3896
rect 2722 3933 2733 3936
rect 2578 3813 2585 3816
rect 2642 3813 2645 3826
rect 2682 3813 2685 3826
rect 2578 3743 2581 3813
rect 2586 3723 2589 3796
rect 2594 3723 2597 3736
rect 2602 3733 2605 3746
rect 2526 3653 2533 3656
rect 2562 3703 2573 3706
rect 2562 3656 2565 3703
rect 2562 3653 2573 3656
rect 2506 3623 2517 3626
rect 2514 3603 2517 3623
rect 2526 3596 2529 3653
rect 2522 3593 2529 3596
rect 2474 3523 2477 3566
rect 2434 3383 2437 3516
rect 2442 3276 2445 3426
rect 2450 3413 2453 3486
rect 2506 3446 2509 3526
rect 2514 3523 2517 3546
rect 2490 3443 2509 3446
rect 2490 3433 2493 3443
rect 2474 3393 2477 3406
rect 2498 3363 2501 3443
rect 2506 3413 2509 3436
rect 2514 3383 2517 3416
rect 2522 3403 2525 3593
rect 2538 3576 2541 3636
rect 2570 3633 2573 3653
rect 2570 3613 2573 3626
rect 2534 3573 2541 3576
rect 2534 3516 2537 3573
rect 2546 3523 2549 3566
rect 2534 3513 2541 3516
rect 2530 3393 2533 3416
rect 2490 3333 2493 3346
rect 2438 3273 2445 3276
rect 2438 3226 2441 3273
rect 2450 3233 2453 3326
rect 2438 3223 2445 3226
rect 2402 3163 2413 3166
rect 2402 3093 2405 3136
rect 2410 3073 2413 3163
rect 2418 3133 2421 3186
rect 2426 3143 2429 3206
rect 2410 3046 2413 3066
rect 2426 3056 2429 3136
rect 2406 3043 2413 3046
rect 2418 3053 2429 3056
rect 2418 3043 2421 3053
rect 2406 2956 2409 3043
rect 2406 2953 2413 2956
rect 2402 2923 2405 2936
rect 2410 2906 2413 2953
rect 2346 2903 2357 2906
rect 2354 2826 2357 2903
rect 2402 2903 2413 2906
rect 2402 2836 2405 2903
rect 2402 2833 2413 2836
rect 2346 2823 2357 2826
rect 2322 2783 2329 2786
rect 2346 2783 2349 2823
rect 2378 2813 2405 2816
rect 2306 2743 2317 2746
rect 2294 2643 2301 2646
rect 2282 2623 2289 2626
rect 2242 2533 2245 2546
rect 2274 2543 2277 2616
rect 2286 2566 2289 2623
rect 2282 2563 2289 2566
rect 2258 2533 2277 2536
rect 2266 2513 2269 2526
rect 2218 2483 2237 2486
rect 2218 2426 2221 2446
rect 2218 2423 2225 2426
rect 2142 2353 2149 2356
rect 2138 2323 2141 2336
rect 2130 2303 2137 2306
rect 2134 2206 2137 2303
rect 2130 2203 2137 2206
rect 2106 2163 2117 2166
rect 2098 2143 2105 2146
rect 2102 1956 2105 2143
rect 2098 1953 2105 1956
rect 2098 1813 2101 1953
rect 2114 1936 2117 2163
rect 2106 1933 2117 1936
rect 2106 1863 2109 1933
rect 2130 1926 2133 2203
rect 2146 2146 2149 2353
rect 2154 2333 2157 2406
rect 2170 2403 2173 2416
rect 2178 2413 2189 2416
rect 2198 2413 2205 2416
rect 2154 2323 2165 2326
rect 2178 2323 2181 2413
rect 2186 2306 2189 2406
rect 2198 2356 2201 2413
rect 2198 2353 2205 2356
rect 2178 2303 2189 2306
rect 2178 2256 2181 2303
rect 2178 2253 2189 2256
rect 2186 2213 2189 2253
rect 2194 2206 2197 2336
rect 2202 2243 2205 2353
rect 2210 2333 2213 2406
rect 2222 2326 2225 2423
rect 2218 2323 2225 2326
rect 2170 2193 2173 2206
rect 2186 2203 2197 2206
rect 2146 2143 2165 2146
rect 2146 2053 2149 2126
rect 2146 2013 2149 2026
rect 2154 2003 2157 2136
rect 2162 2066 2165 2143
rect 2170 2133 2173 2156
rect 2178 2123 2181 2136
rect 2186 2133 2189 2203
rect 2218 2183 2221 2323
rect 2226 2133 2229 2236
rect 2234 2133 2237 2483
rect 2250 2343 2253 2496
rect 2274 2493 2277 2533
rect 2282 2496 2285 2563
rect 2298 2533 2301 2643
rect 2306 2603 2309 2743
rect 2314 2623 2317 2736
rect 2326 2716 2329 2783
rect 2338 2733 2341 2766
rect 2326 2713 2333 2716
rect 2330 2646 2333 2713
rect 2322 2643 2333 2646
rect 2282 2493 2289 2496
rect 2274 2413 2277 2486
rect 2286 2416 2289 2493
rect 2282 2413 2289 2416
rect 2282 2396 2285 2413
rect 2274 2393 2285 2396
rect 2242 2213 2245 2326
rect 2274 2266 2277 2393
rect 2274 2263 2285 2266
rect 2266 2193 2269 2206
rect 2282 2186 2285 2263
rect 2250 2116 2253 2186
rect 2274 2183 2285 2186
rect 2258 2123 2261 2136
rect 2242 2113 2253 2116
rect 2162 2063 2181 2066
rect 2162 1933 2165 2016
rect 2170 2003 2173 2036
rect 2178 1996 2181 2063
rect 2186 2013 2189 2026
rect 2218 1996 2221 2076
rect 2242 2016 2245 2113
rect 2242 2013 2253 2016
rect 2178 1993 2189 1996
rect 2218 1993 2229 1996
rect 2186 1926 2189 1993
rect 2130 1923 2141 1926
rect 2106 1733 2109 1806
rect 2114 1756 2117 1816
rect 2122 1813 2125 1916
rect 2138 1866 2141 1923
rect 2130 1863 2141 1866
rect 2178 1923 2189 1926
rect 2130 1843 2133 1863
rect 2178 1836 2181 1923
rect 2210 1906 2213 1986
rect 2162 1833 2181 1836
rect 2202 1903 2213 1906
rect 2202 1836 2205 1903
rect 2226 1836 2229 1993
rect 2242 1933 2245 1946
rect 2202 1833 2213 1836
rect 2138 1813 2141 1826
rect 2122 1793 2125 1806
rect 2138 1773 2141 1806
rect 2146 1803 2149 1816
rect 2114 1753 2125 1756
rect 2098 1713 2101 1726
rect 2122 1706 2125 1753
rect 2154 1723 2157 1816
rect 2114 1703 2125 1706
rect 2162 1703 2165 1833
rect 2170 1723 2173 1806
rect 2178 1733 2181 1826
rect 2202 1803 2205 1816
rect 2202 1706 2205 1726
rect 2210 1723 2213 1833
rect 2218 1833 2229 1836
rect 2218 1753 2221 1833
rect 2226 1793 2229 1806
rect 2242 1793 2245 1806
rect 2194 1703 2205 1706
rect 2114 1656 2117 1703
rect 2090 1606 2093 1636
rect 2098 1613 2101 1656
rect 2110 1653 2117 1656
rect 2090 1603 2101 1606
rect 2082 1543 2089 1546
rect 2066 1533 2077 1536
rect 2058 1513 2065 1516
rect 2062 1386 2065 1513
rect 2058 1383 2065 1386
rect 2058 1366 2061 1383
rect 2050 1363 2061 1366
rect 2050 1276 2053 1363
rect 2074 1303 2077 1486
rect 2086 1466 2089 1543
rect 2082 1463 2089 1466
rect 2082 1376 2085 1463
rect 2082 1373 2093 1376
rect 2090 1286 2093 1373
rect 2098 1313 2101 1603
rect 2110 1436 2113 1653
rect 2194 1646 2197 1703
rect 2218 1656 2221 1746
rect 2242 1743 2245 1756
rect 2242 1713 2245 1736
rect 2250 1716 2253 2013
rect 2266 2003 2269 2136
rect 2274 2083 2277 2183
rect 2274 2013 2277 2026
rect 2266 1913 2269 1926
rect 2274 1923 2277 2006
rect 2282 2003 2285 2126
rect 2290 2073 2293 2246
rect 2298 2233 2301 2456
rect 2314 2413 2317 2496
rect 2306 2283 2309 2406
rect 2290 1943 2293 2016
rect 2298 2003 2301 2126
rect 2314 2033 2317 2406
rect 2322 2386 2325 2643
rect 2346 2613 2349 2626
rect 2354 2606 2357 2806
rect 2386 2776 2389 2806
rect 2402 2803 2405 2813
rect 2386 2773 2405 2776
rect 2362 2723 2365 2736
rect 2330 2543 2333 2606
rect 2338 2603 2357 2606
rect 2330 2513 2333 2526
rect 2338 2453 2341 2603
rect 2330 2393 2333 2416
rect 2346 2403 2349 2556
rect 2362 2463 2365 2576
rect 2370 2406 2373 2616
rect 2378 2603 2381 2746
rect 2386 2733 2389 2756
rect 2402 2733 2405 2773
rect 2394 2703 2397 2726
rect 2410 2613 2413 2833
rect 2418 2663 2421 3006
rect 2442 2946 2445 3223
rect 2474 3213 2477 3296
rect 2506 3293 2509 3336
rect 2538 3223 2541 3513
rect 2554 3423 2557 3536
rect 2562 3493 2565 3526
rect 2570 3513 2573 3536
rect 2586 3466 2589 3696
rect 2602 3646 2605 3726
rect 2618 3723 2621 3746
rect 2634 3656 2637 3736
rect 2642 3703 2645 3736
rect 2650 3683 2653 3726
rect 2658 3693 2661 3806
rect 2690 3756 2693 3893
rect 2722 3793 2725 3933
rect 2754 3923 2757 4016
rect 2794 4003 2797 4156
rect 2802 4123 2813 4126
rect 2802 4106 2805 4123
rect 2802 4103 2809 4106
rect 2806 4036 2809 4103
rect 2802 4033 2809 4036
rect 2802 4013 2805 4033
rect 2730 3813 2741 3816
rect 2738 3803 2749 3806
rect 2746 3793 2749 3803
rect 2674 3753 2693 3756
rect 2674 3733 2677 3753
rect 2682 3733 2685 3746
rect 2630 3653 2637 3656
rect 2602 3643 2613 3646
rect 2610 3536 2613 3643
rect 2618 3613 2621 3626
rect 2630 3546 2633 3653
rect 2666 3613 2669 3726
rect 2714 3723 2717 3736
rect 2722 3703 2725 3726
rect 2730 3623 2733 3726
rect 2754 3723 2757 3736
rect 2770 3716 2773 3926
rect 2786 3923 2789 3936
rect 2810 3923 2813 4016
rect 2818 4013 2821 4226
rect 2826 4143 2829 4166
rect 2842 4163 2845 4296
rect 2858 4223 2861 4416
rect 2882 4413 2885 4426
rect 2874 4336 2877 4396
rect 2882 4383 2885 4406
rect 2874 4333 2881 4336
rect 2866 4293 2869 4326
rect 2878 4286 2881 4333
rect 2890 4293 2893 4416
rect 2898 4343 2901 4443
rect 2906 4393 2909 4526
rect 2914 4413 2917 4426
rect 2922 4416 2925 4536
rect 2930 4533 2933 4606
rect 2930 4513 2933 4526
rect 2938 4456 2941 4596
rect 2954 4523 2957 4616
rect 3026 4566 3029 4623
rect 3042 4573 3045 4606
rect 3058 4603 3061 4616
rect 3026 4563 3037 4566
rect 2962 4533 2965 4556
rect 3034 4546 3037 4563
rect 3034 4543 3045 4546
rect 2970 4523 2973 4536
rect 3018 4533 3029 4536
rect 2978 4523 2997 4526
rect 2938 4453 2949 4456
rect 2946 4423 2949 4453
rect 2922 4413 2941 4416
rect 2914 4356 2917 4406
rect 2922 4393 2925 4406
rect 2938 4383 2941 4406
rect 2946 4403 2949 4416
rect 2970 4413 2973 4516
rect 2978 4506 2981 4516
rect 3026 4506 3029 4526
rect 2978 4503 2989 4506
rect 2978 4413 2981 4436
rect 2986 4416 2989 4503
rect 3018 4503 3029 4506
rect 3018 4446 3021 4503
rect 3034 4453 3037 4536
rect 3042 4533 3045 4543
rect 3058 4533 3061 4596
rect 3082 4593 3085 4616
rect 3066 4526 3069 4556
rect 3018 4443 3029 4446
rect 2986 4413 2997 4416
rect 2978 4403 2989 4406
rect 2994 4396 2997 4413
rect 2986 4393 2997 4396
rect 3002 4396 3005 4426
rect 3002 4393 3013 4396
rect 2914 4353 2925 4356
rect 2906 4323 2909 4336
rect 2922 4323 2925 4353
rect 2930 4343 2933 4376
rect 2898 4303 2901 4316
rect 2874 4283 2881 4286
rect 2866 4213 2869 4226
rect 2858 4173 2861 4196
rect 2866 4193 2869 4206
rect 2834 4083 2837 4136
rect 2842 4133 2845 4146
rect 2858 4106 2861 4126
rect 2850 4103 2861 4106
rect 2850 4036 2853 4103
rect 2850 4033 2861 4036
rect 2818 3943 2821 4006
rect 2826 4003 2829 4016
rect 2842 4013 2853 4016
rect 2818 3906 2821 3936
rect 2826 3913 2829 3926
rect 2814 3903 2821 3906
rect 2802 3803 2805 3866
rect 2814 3836 2817 3903
rect 2826 3846 2829 3876
rect 2842 3866 2845 4013
rect 2858 4003 2861 4033
rect 2866 3956 2869 4166
rect 2858 3953 2869 3956
rect 2858 3873 2861 3953
rect 2866 3893 2869 3946
rect 2842 3863 2853 3866
rect 2826 3843 2837 3846
rect 2814 3833 2821 3836
rect 2810 3803 2813 3816
rect 2818 3813 2821 3833
rect 2802 3733 2805 3796
rect 2818 3743 2821 3766
rect 2834 3756 2837 3843
rect 2826 3753 2837 3756
rect 2770 3713 2781 3716
rect 2630 3543 2637 3546
rect 2578 3463 2589 3466
rect 2602 3533 2613 3536
rect 2562 3413 2565 3456
rect 2562 3393 2565 3406
rect 2578 3383 2581 3463
rect 2602 3456 2605 3533
rect 2602 3453 2613 3456
rect 2602 3413 2605 3436
rect 2554 3313 2557 3326
rect 2466 3133 2469 3206
rect 2498 3166 2501 3186
rect 2514 3173 2517 3216
rect 2522 3203 2525 3216
rect 2562 3213 2565 3326
rect 2594 3313 2597 3326
rect 2538 3183 2541 3206
rect 2490 3163 2501 3166
rect 2458 3106 2461 3126
rect 2454 3103 2461 3106
rect 2454 3036 2457 3103
rect 2466 3053 2469 3126
rect 2490 3086 2493 3163
rect 2506 3133 2509 3146
rect 2514 3143 2533 3146
rect 2514 3123 2517 3143
rect 2522 3116 2525 3136
rect 2530 3133 2533 3143
rect 2538 3116 2541 3136
rect 2546 3123 2549 3176
rect 2570 3123 2573 3216
rect 2578 3133 2581 3146
rect 2602 3143 2605 3186
rect 2610 3126 2613 3453
rect 2618 3413 2621 3526
rect 2634 3453 2637 3543
rect 2642 3443 2645 3546
rect 2658 3393 2661 3526
rect 2674 3513 2677 3536
rect 2690 3533 2693 3546
rect 2698 3496 2701 3526
rect 2690 3493 2701 3496
rect 2666 3403 2669 3416
rect 2690 3376 2693 3493
rect 2690 3373 2701 3376
rect 2642 3266 2645 3336
rect 2658 3303 2661 3336
rect 2682 3323 2685 3356
rect 2698 3333 2701 3373
rect 2706 3353 2709 3616
rect 2714 3453 2717 3536
rect 2722 3483 2725 3536
rect 2730 3523 2733 3606
rect 2738 3533 2741 3706
rect 2746 3593 2749 3676
rect 2762 3603 2765 3636
rect 2778 3526 2781 3713
rect 2826 3696 2829 3753
rect 2818 3693 2829 3696
rect 2818 3626 2821 3693
rect 2834 3663 2837 3736
rect 2818 3623 2829 3626
rect 2842 3623 2845 3646
rect 2794 3533 2797 3606
rect 2778 3523 2797 3526
rect 2802 3523 2805 3536
rect 2730 3413 2733 3436
rect 2770 3413 2773 3436
rect 2746 3383 2749 3406
rect 2642 3263 2661 3266
rect 2618 3133 2621 3216
rect 2626 3213 2629 3226
rect 2522 3113 2541 3116
rect 2578 3103 2581 3126
rect 2602 3123 2613 3126
rect 2490 3083 2509 3086
rect 2454 3033 2461 3036
rect 2458 3013 2461 3033
rect 2482 2983 2485 3006
rect 2506 3003 2509 3083
rect 2602 3036 2605 3123
rect 2602 3033 2613 3036
rect 2426 2943 2445 2946
rect 2426 2646 2429 2943
rect 2434 2923 2437 2936
rect 2450 2926 2453 2946
rect 2442 2923 2453 2926
rect 2474 2923 2477 2936
rect 2522 2933 2525 2986
rect 2538 2923 2541 3016
rect 2578 2943 2597 2946
rect 2434 2846 2437 2866
rect 2434 2843 2441 2846
rect 2438 2746 2441 2843
rect 2450 2813 2453 2826
rect 2458 2763 2461 2816
rect 2490 2813 2493 2826
rect 2538 2766 2541 2806
rect 2554 2803 2557 2816
rect 2530 2763 2541 2766
rect 2422 2643 2429 2646
rect 2434 2743 2441 2746
rect 2378 2553 2389 2556
rect 2378 2413 2381 2553
rect 2386 2503 2389 2536
rect 2402 2523 2405 2606
rect 2422 2546 2425 2643
rect 2418 2543 2425 2546
rect 2418 2503 2421 2543
rect 2434 2536 2437 2743
rect 2442 2603 2445 2726
rect 2482 2723 2485 2736
rect 2430 2533 2437 2536
rect 2442 2533 2445 2566
rect 2370 2403 2381 2406
rect 2322 2383 2333 2386
rect 2330 2046 2333 2383
rect 2354 2313 2357 2386
rect 2346 2123 2349 2286
rect 2362 2053 2365 2126
rect 2370 2116 2373 2326
rect 2378 2306 2381 2403
rect 2386 2323 2389 2446
rect 2418 2436 2421 2456
rect 2410 2433 2421 2436
rect 2394 2393 2397 2426
rect 2410 2356 2413 2433
rect 2430 2426 2433 2533
rect 2450 2523 2453 2706
rect 2530 2676 2533 2763
rect 2522 2673 2533 2676
rect 2530 2623 2533 2673
rect 2538 2646 2541 2676
rect 2554 2663 2557 2726
rect 2538 2643 2549 2646
rect 2458 2583 2461 2606
rect 2466 2603 2469 2616
rect 2474 2553 2477 2606
rect 2530 2596 2533 2616
rect 2522 2593 2533 2596
rect 2458 2506 2461 2536
rect 2466 2523 2469 2546
rect 2426 2423 2433 2426
rect 2410 2353 2421 2356
rect 2402 2333 2413 2336
rect 2418 2333 2421 2353
rect 2426 2326 2429 2423
rect 2434 2373 2437 2396
rect 2378 2303 2385 2306
rect 2382 2236 2385 2303
rect 2378 2233 2385 2236
rect 2378 2213 2381 2233
rect 2394 2213 2397 2306
rect 2410 2283 2413 2326
rect 2422 2323 2429 2326
rect 2422 2276 2425 2323
rect 2434 2303 2437 2336
rect 2418 2273 2425 2276
rect 2386 2203 2397 2206
rect 2402 2203 2405 2236
rect 2418 2226 2421 2273
rect 2414 2223 2421 2226
rect 2370 2113 2381 2116
rect 2378 2046 2381 2113
rect 2326 2043 2333 2046
rect 2370 2043 2381 2046
rect 2314 2013 2317 2026
rect 2306 1993 2309 2006
rect 2326 1996 2329 2043
rect 2322 1993 2329 1996
rect 2322 1936 2325 1993
rect 2338 1983 2341 2036
rect 2322 1933 2333 1936
rect 2354 1933 2357 1976
rect 2370 1943 2373 2043
rect 2386 1933 2389 2006
rect 2402 1933 2405 2126
rect 2414 2036 2417 2223
rect 2426 2203 2429 2216
rect 2414 2033 2421 2036
rect 2410 2003 2413 2016
rect 2306 1913 2309 1926
rect 2330 1913 2333 1933
rect 2258 1723 2261 1816
rect 2266 1733 2269 1756
rect 2290 1723 2293 1806
rect 2250 1713 2261 1716
rect 2214 1653 2221 1656
rect 2194 1643 2205 1646
rect 2130 1556 2133 1616
rect 2202 1613 2205 1643
rect 2122 1553 2133 1556
rect 2110 1433 2117 1436
rect 2106 1313 2109 1416
rect 2114 1386 2117 1433
rect 2122 1393 2125 1553
rect 2138 1456 2141 1586
rect 2178 1583 2181 1606
rect 2214 1576 2217 1653
rect 2258 1646 2261 1713
rect 2298 1706 2301 1846
rect 2250 1643 2261 1646
rect 2290 1703 2301 1706
rect 2290 1646 2293 1703
rect 2290 1643 2301 1646
rect 2214 1573 2221 1576
rect 2138 1453 2149 1456
rect 2114 1383 2125 1386
rect 2114 1306 2117 1336
rect 2122 1323 2125 1383
rect 2138 1313 2141 1366
rect 2146 1343 2149 1453
rect 2170 1436 2173 1526
rect 2218 1523 2221 1573
rect 2166 1433 2173 1436
rect 2166 1356 2169 1433
rect 2186 1393 2189 1406
rect 2162 1353 2169 1356
rect 2162 1336 2165 1353
rect 2146 1333 2165 1336
rect 2178 1333 2181 1346
rect 2210 1333 2213 1416
rect 2082 1283 2093 1286
rect 2050 1273 2069 1276
rect 2034 1113 2037 1126
rect 2010 1103 2021 1106
rect 2018 1036 2021 1103
rect 2010 1033 2021 1036
rect 2010 986 2013 1033
rect 2018 996 2021 1006
rect 2026 1003 2029 1016
rect 2034 996 2037 1016
rect 2042 1003 2045 1196
rect 2066 1156 2069 1273
rect 2050 1153 2069 1156
rect 2082 1156 2085 1283
rect 2098 1166 2101 1306
rect 2106 1303 2125 1306
rect 2122 1233 2125 1303
rect 2130 1226 2133 1306
rect 2106 1223 2133 1226
rect 2106 1206 2109 1223
rect 2106 1203 2117 1206
rect 2098 1163 2105 1166
rect 2082 1153 2093 1156
rect 2050 1043 2053 1153
rect 2058 1123 2061 1136
rect 2082 1113 2085 1136
rect 2090 1096 2093 1153
rect 2082 1093 2093 1096
rect 2018 993 2037 996
rect 2010 983 2029 986
rect 1990 893 1997 896
rect 1962 783 1965 806
rect 1874 723 1885 726
rect 1898 703 1901 726
rect 1914 723 1925 726
rect 1874 596 1877 616
rect 1874 593 1881 596
rect 1878 506 1881 593
rect 1890 523 1893 616
rect 1914 603 1917 723
rect 1946 713 1949 726
rect 1914 533 1917 596
rect 1878 503 1885 506
rect 1882 446 1885 503
rect 1874 443 1885 446
rect 1842 383 1845 406
rect 1874 386 1877 443
rect 1898 413 1901 426
rect 1890 393 1893 406
rect 1874 383 1885 386
rect 1770 333 1773 346
rect 1746 293 1757 296
rect 1746 226 1749 293
rect 1738 223 1749 226
rect 1714 133 1717 146
rect 1730 133 1733 216
rect 1738 206 1741 223
rect 1738 203 1749 206
rect 1754 203 1757 226
rect 1762 213 1765 326
rect 1778 276 1781 326
rect 1770 273 1781 276
rect 1770 203 1773 273
rect 1746 193 1749 203
rect 1778 173 1781 236
rect 1690 113 1693 126
rect 1730 113 1733 126
rect 1786 123 1789 206
rect 1802 203 1805 216
rect 1818 213 1821 246
rect 1810 193 1813 206
rect 1826 203 1829 216
rect 1858 213 1861 326
rect 1882 216 1885 383
rect 1906 323 1909 436
rect 1922 426 1925 526
rect 1930 523 1933 706
rect 1954 606 1957 766
rect 1970 703 1973 816
rect 1994 743 1997 893
rect 2018 876 2021 976
rect 2010 873 2021 876
rect 2010 806 2013 873
rect 2026 813 2029 983
rect 2042 933 2045 976
rect 2034 896 2037 926
rect 2042 913 2045 926
rect 2034 893 2041 896
rect 2038 826 2041 893
rect 2034 823 2041 826
rect 2010 803 2021 806
rect 2034 803 2037 823
rect 1994 723 1997 736
rect 2010 716 2013 746
rect 2018 723 2021 803
rect 2010 713 2021 716
rect 2018 696 2021 713
rect 2010 693 2021 696
rect 2010 636 2013 693
rect 2034 656 2037 726
rect 2034 653 2045 656
rect 2010 633 2021 636
rect 1946 603 1957 606
rect 1914 403 1917 426
rect 1922 423 1933 426
rect 1922 413 1925 423
rect 1874 213 1885 216
rect 1922 213 1925 226
rect 1866 183 1869 206
rect 1874 176 1877 213
rect 1866 173 1877 176
rect 1866 133 1869 173
rect 1882 133 1885 206
rect 1842 113 1845 126
rect 1882 113 1885 126
rect 1930 123 1933 206
rect 1938 196 1941 216
rect 1946 203 1949 603
rect 1962 593 1965 616
rect 1954 543 1973 546
rect 1954 523 1957 543
rect 1962 523 1965 536
rect 1970 533 1973 543
rect 1970 483 1973 526
rect 1954 323 1957 416
rect 1962 393 1965 406
rect 1970 383 1973 416
rect 1986 266 1989 566
rect 2010 523 2013 616
rect 2018 596 2021 633
rect 2018 593 2029 596
rect 1994 473 2005 476
rect 1994 396 1997 416
rect 2002 403 2005 473
rect 2026 436 2029 593
rect 2042 563 2045 653
rect 2050 633 2053 1016
rect 2058 1013 2061 1036
rect 2082 1026 2085 1093
rect 2102 1086 2105 1163
rect 2098 1083 2105 1086
rect 2082 1023 2093 1026
rect 2058 803 2061 926
rect 2066 833 2069 1006
rect 2090 1003 2093 1023
rect 2098 986 2101 1083
rect 2114 1036 2117 1203
rect 2094 983 2101 986
rect 2106 1033 2117 1036
rect 2074 876 2077 936
rect 2082 903 2085 916
rect 2074 873 2085 876
rect 2058 706 2061 796
rect 2066 723 2069 816
rect 2058 703 2065 706
rect 2062 636 2065 703
rect 2058 633 2065 636
rect 2058 613 2061 633
rect 2050 556 2053 586
rect 2074 563 2077 826
rect 2082 803 2085 873
rect 2094 816 2097 983
rect 2106 823 2109 1033
rect 2114 886 2117 1016
rect 2130 933 2133 1206
rect 2138 1183 2141 1236
rect 2138 1013 2141 1126
rect 2146 1106 2149 1333
rect 2154 1113 2157 1326
rect 2146 1103 2157 1106
rect 2162 1086 2165 1316
rect 2170 1153 2173 1216
rect 2158 1083 2165 1086
rect 2114 883 2133 886
rect 2130 826 2133 883
rect 2146 873 2149 1046
rect 2158 946 2161 1083
rect 2158 943 2165 946
rect 2154 836 2157 926
rect 2162 923 2165 943
rect 2170 916 2173 1116
rect 2138 833 2157 836
rect 2162 913 2173 916
rect 2130 823 2141 826
rect 2094 813 2101 816
rect 2130 813 2133 823
rect 2098 723 2101 813
rect 2146 783 2149 826
rect 2162 813 2165 913
rect 2170 813 2173 826
rect 2162 746 2165 806
rect 2162 743 2169 746
rect 2138 686 2141 736
rect 2166 696 2169 743
rect 2162 693 2169 696
rect 2138 683 2149 686
rect 2042 553 2053 556
rect 2042 523 2045 553
rect 2098 536 2101 616
rect 2082 533 2101 536
rect 2122 533 2125 546
rect 2082 516 2085 533
rect 2078 513 2085 516
rect 2078 456 2081 513
rect 2078 453 2085 456
rect 2026 433 2037 436
rect 2010 416 2013 426
rect 2010 413 2021 416
rect 2010 396 2013 406
rect 1994 393 2013 396
rect 2002 323 2005 336
rect 2018 326 2021 413
rect 2034 376 2037 433
rect 2066 413 2069 426
rect 2074 413 2077 436
rect 2082 396 2085 453
rect 2010 323 2021 326
rect 2026 373 2037 376
rect 2074 393 2085 396
rect 1986 263 1997 266
rect 1954 216 1957 236
rect 1954 213 1965 216
rect 1954 196 1957 206
rect 1938 193 1957 196
rect 1962 153 1965 213
rect 1986 123 1989 216
rect 1994 196 1997 263
rect 2002 203 2005 296
rect 2010 213 2013 323
rect 2026 306 2029 373
rect 2042 323 2045 346
rect 2050 333 2053 356
rect 2058 313 2061 326
rect 2026 303 2037 306
rect 2034 236 2037 303
rect 2074 266 2077 393
rect 2074 263 2085 266
rect 2026 233 2037 236
rect 1994 193 2013 196
rect 2010 133 2013 193
rect 2026 156 2029 233
rect 2050 213 2061 216
rect 2026 153 2033 156
rect 2030 106 2033 153
rect 2042 123 2045 206
rect 2050 203 2061 206
rect 2066 183 2069 246
rect 2074 203 2077 216
rect 2026 103 2033 106
rect 2026 83 2029 103
rect 2082 86 2085 263
rect 2090 216 2093 526
rect 2138 506 2141 576
rect 2146 543 2149 683
rect 2162 613 2165 693
rect 2178 676 2181 1316
rect 2202 1276 2205 1316
rect 2194 1273 2205 1276
rect 2194 1226 2197 1273
rect 2194 1223 2205 1226
rect 2202 1203 2205 1223
rect 2210 1186 2213 1326
rect 2218 1313 2221 1456
rect 2226 1413 2229 1506
rect 2234 1363 2237 1616
rect 2250 1596 2253 1643
rect 2250 1593 2261 1596
rect 2242 1503 2245 1526
rect 2250 1366 2253 1446
rect 2258 1436 2261 1593
rect 2282 1583 2285 1606
rect 2266 1513 2269 1526
rect 2274 1513 2277 1576
rect 2274 1456 2277 1506
rect 2298 1503 2301 1643
rect 2306 1613 2309 1806
rect 2314 1803 2317 1816
rect 2322 1813 2325 1856
rect 2314 1573 2317 1736
rect 2322 1566 2325 1756
rect 2338 1723 2341 1816
rect 2346 1813 2349 1826
rect 2362 1763 2365 1816
rect 2378 1813 2381 1916
rect 2410 1913 2413 1926
rect 2418 1826 2421 2033
rect 2426 1843 2429 2196
rect 2442 2183 2445 2506
rect 2454 2503 2461 2506
rect 2522 2506 2525 2593
rect 2546 2586 2549 2643
rect 2538 2583 2549 2586
rect 2538 2523 2541 2583
rect 2562 2553 2565 2926
rect 2570 2916 2573 2936
rect 2578 2933 2581 2943
rect 2570 2913 2577 2916
rect 2574 2636 2577 2913
rect 2570 2633 2577 2636
rect 2570 2613 2573 2633
rect 2554 2543 2573 2546
rect 2546 2513 2549 2536
rect 2554 2523 2557 2543
rect 2562 2523 2565 2536
rect 2570 2533 2573 2543
rect 2522 2503 2533 2506
rect 2454 2426 2457 2503
rect 2454 2423 2461 2426
rect 2450 2283 2453 2406
rect 2458 2333 2461 2423
rect 2466 2323 2469 2476
rect 2474 2383 2477 2456
rect 2434 2136 2437 2166
rect 2434 2133 2445 2136
rect 2434 2083 2437 2126
rect 2450 2123 2453 2136
rect 2458 2133 2461 2206
rect 2434 2003 2437 2036
rect 2434 1926 2437 1946
rect 2434 1923 2441 1926
rect 2438 1836 2441 1923
rect 2458 1913 2461 1926
rect 2466 1883 2469 2186
rect 2490 1973 2493 2256
rect 2498 2213 2501 2326
rect 2506 2323 2509 2336
rect 2530 2323 2533 2503
rect 2554 2376 2557 2416
rect 2570 2403 2573 2526
rect 2578 2393 2581 2416
rect 2554 2373 2573 2376
rect 2570 2323 2573 2373
rect 2530 2193 2533 2316
rect 2578 2276 2581 2326
rect 2546 2213 2549 2276
rect 2570 2273 2581 2276
rect 2554 2206 2557 2246
rect 2546 2203 2557 2206
rect 2506 2053 2509 2136
rect 2506 2003 2509 2026
rect 2506 1933 2509 1976
rect 2522 1896 2525 2136
rect 2530 2106 2533 2186
rect 2546 2123 2549 2203
rect 2570 2196 2573 2273
rect 2586 2203 2589 2936
rect 2594 2923 2597 2943
rect 2602 2933 2605 3016
rect 2610 2933 2613 3033
rect 2618 3013 2621 3026
rect 2610 2903 2613 2926
rect 2618 2863 2621 2926
rect 2626 2923 2629 3206
rect 2658 3196 2661 3263
rect 2674 3196 2677 3216
rect 2682 3203 2685 3316
rect 2698 3313 2701 3326
rect 2714 3246 2717 3336
rect 2714 3243 2725 3246
rect 2690 3196 2693 3206
rect 2658 3193 2669 3196
rect 2674 3193 2693 3196
rect 2634 3143 2653 3146
rect 2634 3123 2637 3143
rect 2642 3103 2645 3136
rect 2650 3133 2653 3143
rect 2634 2996 2637 3016
rect 2642 3003 2645 3046
rect 2650 2996 2653 3006
rect 2634 2993 2653 2996
rect 2618 2823 2637 2826
rect 2618 2816 2621 2823
rect 2610 2813 2621 2816
rect 2626 2783 2629 2806
rect 2634 2803 2637 2823
rect 2602 2733 2605 2746
rect 2594 2723 2605 2726
rect 2594 2506 2597 2556
rect 2610 2523 2613 2726
rect 2618 2723 2621 2736
rect 2642 2723 2645 2906
rect 2650 2886 2653 2986
rect 2658 2903 2661 3176
rect 2666 3156 2669 3193
rect 2698 3173 2701 3216
rect 2666 3153 2685 3156
rect 2682 3046 2685 3153
rect 2706 3123 2709 3136
rect 2722 3056 2725 3243
rect 2738 3213 2741 3326
rect 2738 3183 2741 3206
rect 2786 3166 2789 3523
rect 2810 3516 2813 3606
rect 2826 3526 2829 3623
rect 2834 3543 2837 3556
rect 2850 3536 2853 3863
rect 2874 3816 2877 4283
rect 2882 4203 2885 4246
rect 2890 4193 2893 4216
rect 2898 4146 2901 4206
rect 2882 4143 2901 4146
rect 2882 4023 2885 4143
rect 2890 4116 2893 4136
rect 2890 4113 2901 4116
rect 2922 4113 2925 4226
rect 2898 4036 2901 4113
rect 2930 4096 2933 4316
rect 2954 4263 2957 4336
rect 2962 4323 2973 4326
rect 2978 4303 2981 4336
rect 2986 4226 2989 4393
rect 2994 4306 2997 4346
rect 3010 4326 3013 4393
rect 3018 4333 3021 4406
rect 3026 4403 3029 4443
rect 3010 4323 3021 4326
rect 2994 4303 3005 4306
rect 2938 4213 2941 4226
rect 2954 4203 2957 4216
rect 2890 4033 2901 4036
rect 2922 4093 2933 4096
rect 2890 4016 2893 4033
rect 2922 4026 2925 4093
rect 2922 4023 2933 4026
rect 2882 4013 2893 4016
rect 2882 3923 2885 4013
rect 2890 3983 2893 4006
rect 2890 3933 2893 3946
rect 2898 3873 2901 3936
rect 2906 3923 2909 3936
rect 2914 3923 2917 4006
rect 2866 3813 2877 3816
rect 2866 3736 2869 3813
rect 2922 3806 2925 3916
rect 2930 3896 2933 4023
rect 2938 4006 2941 4116
rect 2938 4003 2949 4006
rect 2946 3946 2949 4003
rect 2938 3943 2949 3946
rect 2938 3913 2941 3943
rect 2962 3936 2965 4226
rect 2970 4193 2973 4226
rect 2978 4223 2989 4226
rect 2978 4123 2981 4216
rect 2994 4213 2997 4226
rect 3002 4163 3005 4303
rect 3018 4223 3021 4323
rect 3034 4293 3037 4406
rect 3042 4376 3045 4526
rect 3066 4523 3085 4526
rect 3050 4393 3053 4406
rect 3058 4403 3061 4416
rect 3066 4376 3069 4506
rect 3090 4503 3093 4536
rect 3138 4533 3141 4616
rect 3146 4533 3149 4666
rect 3250 4656 3253 4736
rect 3242 4653 3253 4656
rect 3186 4596 3189 4616
rect 3202 4603 3205 4616
rect 3178 4593 3189 4596
rect 3178 4526 3181 4593
rect 3202 4533 3205 4596
rect 3226 4593 3229 4616
rect 3242 4576 3245 4653
rect 3146 4493 3149 4526
rect 3178 4523 3189 4526
rect 3210 4523 3213 4576
rect 3242 4573 3253 4576
rect 3074 4413 3077 4456
rect 3106 4393 3109 4416
rect 3042 4373 3053 4376
rect 3066 4373 3077 4376
rect 3050 4326 3053 4373
rect 3042 4323 3053 4326
rect 3066 4326 3069 4336
rect 3074 4333 3077 4373
rect 3066 4323 3085 4326
rect 3026 4203 3029 4216
rect 3034 4186 3037 4236
rect 3030 4183 3037 4186
rect 3018 4123 3021 4136
rect 3030 4116 3033 4183
rect 3042 4123 3045 4323
rect 3082 4306 3085 4323
rect 3074 4303 3085 4306
rect 3074 4236 3077 4303
rect 3074 4233 3085 4236
rect 3050 4186 3053 4206
rect 3058 4203 3061 4216
rect 3082 4213 3085 4233
rect 3090 4223 3093 4336
rect 3098 4303 3101 4326
rect 3106 4286 3109 4336
rect 3114 4316 3117 4356
rect 3154 4323 3157 4416
rect 3186 4403 3189 4523
rect 3218 4503 3221 4536
rect 3250 4456 3253 4573
rect 3274 4523 3277 4536
rect 3282 4533 3285 4606
rect 3314 4573 3317 4616
rect 3346 4603 3349 4616
rect 3370 4603 3373 4616
rect 3306 4533 3309 4546
rect 3290 4493 3293 4526
rect 3314 4523 3317 4536
rect 3330 4533 3333 4596
rect 3426 4593 3429 4616
rect 3250 4453 3257 4456
rect 3178 4323 3181 4336
rect 3186 4333 3189 4396
rect 3210 4393 3213 4416
rect 3254 4376 3257 4453
rect 3250 4373 3257 4376
rect 3202 4333 3205 4346
rect 3114 4313 3125 4316
rect 3102 4283 3109 4286
rect 3082 4193 3085 4206
rect 3102 4186 3105 4283
rect 3122 4266 3125 4313
rect 3114 4263 3125 4266
rect 3114 4193 3117 4263
rect 3146 4213 3149 4226
rect 3050 4183 3061 4186
rect 3102 4183 3109 4186
rect 3030 4113 3037 4116
rect 2962 3933 2973 3936
rect 2930 3893 2937 3896
rect 2866 3733 2877 3736
rect 2882 3733 2885 3806
rect 2914 3803 2925 3806
rect 2914 3756 2917 3803
rect 2914 3753 2925 3756
rect 2866 3696 2869 3716
rect 2862 3693 2869 3696
rect 2862 3606 2865 3693
rect 2862 3603 2869 3606
rect 2866 3583 2869 3603
rect 2874 3566 2877 3733
rect 2914 3716 2917 3736
rect 2906 3713 2917 3716
rect 2906 3666 2909 3713
rect 2906 3663 2917 3666
rect 2890 3596 2893 3646
rect 2898 3603 2901 3616
rect 2914 3613 2917 3663
rect 2922 3623 2925 3753
rect 2934 3656 2937 3893
rect 2954 3816 2957 3926
rect 2970 3846 2973 3933
rect 2930 3653 2937 3656
rect 2946 3813 2957 3816
rect 2962 3843 2973 3846
rect 2890 3593 2901 3596
rect 2906 3593 2909 3606
rect 2870 3563 2877 3566
rect 2794 3513 2813 3516
rect 2818 3523 2829 3526
rect 2818 3496 2821 3523
rect 2814 3493 2821 3496
rect 2814 3426 2817 3493
rect 2826 3426 2829 3516
rect 2834 3513 2837 3526
rect 2842 3513 2845 3536
rect 2850 3533 2861 3536
rect 2814 3423 2821 3426
rect 2818 3406 2821 3423
rect 2826 3423 2845 3426
rect 2826 3413 2829 3423
rect 2818 3403 2825 3406
rect 2802 3333 2805 3346
rect 2794 3313 2797 3326
rect 2802 3203 2805 3216
rect 2786 3163 2793 3166
rect 2746 3123 2749 3136
rect 2790 3086 2793 3163
rect 2802 3103 2805 3126
rect 2786 3083 2793 3086
rect 2786 3056 2789 3083
rect 2666 3043 2685 3046
rect 2714 3053 2725 3056
rect 2782 3053 2789 3056
rect 2666 2983 2669 3043
rect 2698 3013 2701 3026
rect 2714 2956 2717 3053
rect 2738 3013 2741 3026
rect 2782 2986 2785 3053
rect 2794 3013 2797 3046
rect 2810 2986 2813 3346
rect 2822 3266 2825 3403
rect 2834 3343 2837 3416
rect 2842 3403 2845 3423
rect 2858 3413 2861 3533
rect 2870 3336 2873 3563
rect 2882 3533 2885 3556
rect 2882 3513 2885 3526
rect 2890 3523 2893 3536
rect 2898 3513 2901 3593
rect 2914 3566 2917 3586
rect 2910 3563 2917 3566
rect 2910 3486 2913 3563
rect 2910 3483 2917 3486
rect 2822 3263 2829 3266
rect 2826 3246 2829 3263
rect 2834 3253 2837 3336
rect 2842 3323 2845 3336
rect 2870 3333 2877 3336
rect 2826 3243 2837 3246
rect 2834 3106 2837 3243
rect 2826 3103 2837 3106
rect 2826 3036 2829 3103
rect 2826 3033 2837 3036
rect 2826 2993 2829 3016
rect 2706 2953 2717 2956
rect 2650 2883 2661 2886
rect 2658 2716 2661 2883
rect 2674 2823 2677 2926
rect 2690 2903 2693 2926
rect 2698 2803 2701 2826
rect 2642 2713 2661 2716
rect 2642 2556 2645 2713
rect 2690 2683 2693 2726
rect 2706 2656 2709 2953
rect 2714 2933 2717 2946
rect 2730 2933 2733 2986
rect 2782 2983 2789 2986
rect 2810 2983 2829 2986
rect 2786 2966 2789 2983
rect 2786 2963 2797 2966
rect 2794 2946 2797 2963
rect 2794 2943 2801 2946
rect 2730 2816 2733 2906
rect 2714 2803 2717 2816
rect 2726 2813 2733 2816
rect 2754 2813 2757 2926
rect 2798 2886 2801 2943
rect 2810 2923 2813 2946
rect 2818 2933 2821 2966
rect 2826 2906 2829 2983
rect 2834 2923 2837 3033
rect 2842 3013 2845 3206
rect 2842 2983 2845 3006
rect 2850 2936 2853 3236
rect 2858 3213 2861 3226
rect 2858 3076 2861 3206
rect 2866 3203 2869 3316
rect 2874 3213 2877 3333
rect 2882 3216 2885 3466
rect 2914 3463 2917 3483
rect 2898 3423 2901 3436
rect 2922 3433 2925 3606
rect 2930 3583 2933 3653
rect 2946 3636 2949 3813
rect 2954 3723 2957 3736
rect 2962 3723 2965 3843
rect 2970 3803 2973 3826
rect 2986 3793 2989 4036
rect 3002 3983 3005 4006
rect 3002 3893 3005 3936
rect 3018 3736 3021 4106
rect 3034 4043 3037 4113
rect 3058 4066 3061 4183
rect 3098 4116 3101 4136
rect 3050 4063 3061 4066
rect 3090 4113 3101 4116
rect 3090 4066 3093 4113
rect 3106 4093 3109 4183
rect 3186 4173 3189 4326
rect 3194 4276 3197 4326
rect 3210 4323 3213 4336
rect 3234 4306 3237 4326
rect 3226 4303 3237 4306
rect 3194 4273 3205 4276
rect 3202 4213 3205 4273
rect 3226 4236 3229 4303
rect 3226 4233 3237 4236
rect 3234 4216 3237 4233
rect 3226 4213 3237 4216
rect 3114 4116 3117 4136
rect 3154 4133 3157 4146
rect 3146 4116 3149 4126
rect 3154 4123 3165 4126
rect 3114 4113 3125 4116
rect 3146 4113 3157 4116
rect 3090 4063 3101 4066
rect 3050 4013 3053 4063
rect 3098 4013 3101 4063
rect 3122 4006 3125 4113
rect 3114 4003 3125 4006
rect 3066 3923 3069 3956
rect 3018 3733 3029 3736
rect 3034 3733 3037 3816
rect 3066 3766 3069 3916
rect 3114 3913 3117 4003
rect 3154 3976 3157 4113
rect 3178 4036 3181 4136
rect 3202 4133 3205 4206
rect 3218 4193 3221 4206
rect 3242 4193 3245 4206
rect 3250 4196 3253 4373
rect 3266 4336 3269 4416
rect 3258 4333 3269 4336
rect 3274 4316 3277 4336
rect 3266 4313 3277 4316
rect 3266 4246 3269 4313
rect 3282 4256 3285 4446
rect 3306 4266 3309 4456
rect 3338 4453 3341 4516
rect 3330 4393 3333 4416
rect 3346 4383 3349 4506
rect 3354 4443 3357 4526
rect 3394 4523 3397 4536
rect 3442 4533 3445 4616
rect 3458 4533 3461 4566
rect 3498 4533 3501 4616
rect 3530 4593 3533 4606
rect 3578 4593 3581 4606
rect 3538 4533 3541 4556
rect 3370 4503 3373 4516
rect 3362 4386 3365 4416
rect 3354 4383 3365 4386
rect 3354 4333 3357 4383
rect 3298 4263 3309 4266
rect 3282 4253 3289 4256
rect 3266 4243 3277 4246
rect 3258 4213 3261 4226
rect 3274 4213 3277 4243
rect 3250 4193 3261 4196
rect 3218 4076 3221 4176
rect 3242 4123 3245 4146
rect 3258 4116 3261 4193
rect 3274 4183 3277 4206
rect 3286 4196 3289 4253
rect 3282 4193 3289 4196
rect 3282 4173 3285 4193
rect 3210 4073 3221 4076
rect 3250 4113 3261 4116
rect 3178 4033 3189 4036
rect 3154 3973 3165 3976
rect 3122 3893 3125 3926
rect 3130 3836 3133 3936
rect 3154 3933 3157 3956
rect 3146 3893 3149 3926
rect 3122 3833 3133 3836
rect 3058 3763 3069 3766
rect 3002 3723 3021 3726
rect 2970 3703 2973 3716
rect 2938 3633 2949 3636
rect 2938 3536 2941 3633
rect 2946 3603 2949 3626
rect 2930 3533 2941 3536
rect 2930 3506 2933 3533
rect 2962 3523 2965 3676
rect 3026 3673 3029 3733
rect 3058 3636 3061 3763
rect 3082 3746 3085 3826
rect 3074 3733 3077 3746
rect 3082 3743 3093 3746
rect 3058 3633 3069 3636
rect 3066 3616 3069 3633
rect 3010 3593 3013 3616
rect 3050 3613 3061 3616
rect 3066 3613 3077 3616
rect 2930 3503 2949 3506
rect 2906 3413 2925 3416
rect 2890 3393 2893 3406
rect 2906 3403 2909 3413
rect 2946 3406 2949 3503
rect 2978 3413 2981 3536
rect 3002 3533 3005 3566
rect 3018 3536 3021 3576
rect 3010 3533 3021 3536
rect 3010 3493 3013 3533
rect 3018 3513 3021 3526
rect 3026 3523 3029 3566
rect 3034 3413 3037 3536
rect 3066 3533 3069 3606
rect 3042 3513 3045 3526
rect 2930 3403 2949 3406
rect 2930 3326 2933 3403
rect 2970 3393 2973 3406
rect 2962 3333 2965 3346
rect 2890 3223 2893 3326
rect 2882 3213 2893 3216
rect 2882 3143 2885 3156
rect 2858 3073 2869 3076
rect 2858 3003 2861 3046
rect 2866 3013 2869 3073
rect 2850 2933 2857 2936
rect 2794 2883 2801 2886
rect 2818 2903 2829 2906
rect 2726 2756 2729 2813
rect 2726 2753 2733 2756
rect 2690 2653 2709 2656
rect 2690 2586 2693 2653
rect 2714 2613 2717 2686
rect 2634 2553 2645 2556
rect 2666 2583 2693 2586
rect 2634 2506 2637 2553
rect 2666 2533 2669 2583
rect 2650 2513 2653 2526
rect 2690 2513 2693 2526
rect 2594 2503 2613 2506
rect 2634 2503 2653 2506
rect 2610 2376 2613 2503
rect 2642 2413 2645 2426
rect 2594 2373 2613 2376
rect 2570 2193 2581 2196
rect 2578 2146 2581 2193
rect 2594 2186 2597 2373
rect 2634 2356 2637 2406
rect 2650 2396 2653 2503
rect 2658 2403 2661 2416
rect 2650 2393 2661 2396
rect 2634 2353 2641 2356
rect 2618 2313 2621 2336
rect 2638 2306 2641 2353
rect 2562 2143 2581 2146
rect 2590 2183 2597 2186
rect 2554 2113 2557 2126
rect 2530 2103 2541 2106
rect 2538 1916 2541 2103
rect 2554 2013 2557 2036
rect 2562 1996 2565 2143
rect 2554 1993 2565 1996
rect 2554 1946 2557 1993
rect 2554 1943 2565 1946
rect 2562 1923 2565 1943
rect 2518 1893 2525 1896
rect 2530 1913 2541 1916
rect 2518 1836 2521 1893
rect 2530 1866 2533 1913
rect 2530 1863 2541 1866
rect 2434 1833 2441 1836
rect 2418 1823 2429 1826
rect 2410 1813 2421 1816
rect 2410 1723 2413 1806
rect 2426 1756 2429 1823
rect 2434 1813 2437 1833
rect 2482 1813 2485 1826
rect 2450 1793 2453 1806
rect 2418 1753 2429 1756
rect 2386 1623 2389 1666
rect 2362 1603 2365 1616
rect 2322 1563 2329 1566
rect 2314 1486 2317 1526
rect 2306 1483 2317 1486
rect 2274 1453 2285 1456
rect 2258 1433 2269 1436
rect 2266 1376 2269 1433
rect 2246 1363 2253 1366
rect 2258 1373 2269 1376
rect 2246 1316 2249 1363
rect 2258 1323 2261 1373
rect 2282 1356 2285 1453
rect 2306 1406 2309 1483
rect 2326 1476 2329 1563
rect 2338 1533 2341 1596
rect 2386 1583 2389 1606
rect 2338 1506 2341 1526
rect 2378 1523 2381 1566
rect 2338 1503 2349 1506
rect 2322 1473 2329 1476
rect 2322 1413 2325 1473
rect 2346 1406 2349 1503
rect 2306 1403 2317 1406
rect 2314 1366 2317 1403
rect 2338 1403 2349 1406
rect 2314 1363 2325 1366
rect 2274 1353 2285 1356
rect 2274 1323 2277 1353
rect 2246 1313 2253 1316
rect 2250 1263 2253 1313
rect 2274 1213 2277 1226
rect 2206 1183 2213 1186
rect 2186 943 2189 1166
rect 2194 1013 2197 1106
rect 2206 976 2209 1183
rect 2218 1126 2221 1186
rect 2226 1143 2229 1206
rect 2218 1123 2237 1126
rect 2218 1003 2221 1123
rect 2206 973 2213 976
rect 2210 953 2213 973
rect 2194 923 2197 936
rect 2210 896 2213 946
rect 2202 893 2213 896
rect 2186 823 2189 866
rect 2194 813 2197 836
rect 2202 743 2205 893
rect 2234 886 2237 956
rect 2210 883 2237 886
rect 2174 673 2181 676
rect 2174 596 2177 673
rect 2174 593 2181 596
rect 2178 573 2181 593
rect 2162 533 2165 546
rect 2130 503 2141 506
rect 2106 413 2109 426
rect 2098 323 2109 326
rect 2090 213 2097 216
rect 2094 116 2097 213
rect 2106 123 2109 216
rect 2114 213 2117 486
rect 2130 446 2133 503
rect 2186 486 2189 726
rect 2210 566 2213 883
rect 2218 723 2221 876
rect 2242 856 2245 1166
rect 2274 1113 2277 1196
rect 2290 1176 2293 1276
rect 2282 1173 2293 1176
rect 2282 1096 2285 1173
rect 2298 1156 2301 1336
rect 2322 1286 2325 1363
rect 2338 1333 2341 1403
rect 2386 1346 2389 1496
rect 2402 1453 2405 1676
rect 2410 1613 2413 1626
rect 2418 1596 2421 1753
rect 2414 1593 2421 1596
rect 2426 1743 2445 1746
rect 2414 1516 2417 1593
rect 2426 1523 2429 1743
rect 2434 1623 2437 1736
rect 2442 1733 2445 1743
rect 2482 1733 2485 1766
rect 2490 1713 2493 1726
rect 2506 1713 2509 1836
rect 2518 1833 2525 1836
rect 2522 1813 2525 1833
rect 2530 1803 2533 1826
rect 2538 1773 2541 1863
rect 2546 1763 2549 1816
rect 2554 1796 2557 1896
rect 2562 1813 2565 1886
rect 2570 1876 2573 2136
rect 2590 2126 2593 2183
rect 2602 2133 2605 2206
rect 2610 2196 2613 2216
rect 2618 2203 2621 2306
rect 2634 2303 2641 2306
rect 2634 2213 2637 2303
rect 2658 2226 2661 2393
rect 2682 2333 2685 2366
rect 2706 2363 2709 2406
rect 2714 2403 2717 2426
rect 2658 2223 2669 2226
rect 2626 2196 2629 2206
rect 2610 2193 2629 2196
rect 2626 2143 2645 2146
rect 2590 2123 2597 2126
rect 2626 2123 2629 2143
rect 2578 2013 2581 2066
rect 2578 1923 2581 1946
rect 2586 1923 2589 1936
rect 2594 1906 2597 2123
rect 2634 2116 2637 2136
rect 2642 2133 2645 2143
rect 2650 2116 2653 2206
rect 2634 2113 2653 2116
rect 2602 2013 2605 2026
rect 2602 1933 2605 1946
rect 2618 1923 2621 2066
rect 2658 2063 2661 2216
rect 2666 2176 2669 2223
rect 2690 2213 2693 2326
rect 2730 2236 2733 2753
rect 2738 2723 2741 2806
rect 2746 2783 2749 2806
rect 2778 2756 2781 2816
rect 2778 2753 2785 2756
rect 2738 2526 2741 2596
rect 2754 2543 2757 2586
rect 2762 2533 2765 2686
rect 2770 2613 2773 2746
rect 2782 2676 2785 2753
rect 2794 2706 2797 2883
rect 2818 2806 2821 2903
rect 2842 2886 2845 2926
rect 2834 2883 2845 2886
rect 2834 2836 2837 2883
rect 2854 2846 2857 2933
rect 2866 2896 2869 2946
rect 2874 2943 2877 2996
rect 2890 2953 2893 3213
rect 2906 3203 2909 3326
rect 2922 3323 2933 3326
rect 2970 3323 2973 3336
rect 2994 3323 3013 3326
rect 2922 3256 2925 3323
rect 2922 3253 2933 3256
rect 2930 3233 2933 3253
rect 2914 3203 2917 3226
rect 2938 3223 2941 3316
rect 2906 3093 2909 3196
rect 2922 3133 2925 3216
rect 2930 3203 2933 3216
rect 2930 3113 2933 3126
rect 2946 3096 2949 3216
rect 2930 3093 2949 3096
rect 2930 2996 2933 3093
rect 2954 3003 2957 3126
rect 2930 2993 2949 2996
rect 2890 2913 2893 2926
rect 2866 2893 2877 2896
rect 2850 2843 2857 2846
rect 2834 2833 2845 2836
rect 2842 2813 2845 2833
rect 2818 2803 2829 2806
rect 2802 2743 2805 2756
rect 2810 2723 2813 2786
rect 2826 2753 2829 2803
rect 2834 2723 2837 2736
rect 2842 2723 2845 2806
rect 2794 2703 2805 2706
rect 2778 2673 2785 2676
rect 2738 2523 2749 2526
rect 2778 2523 2781 2673
rect 2802 2626 2805 2703
rect 2794 2623 2805 2626
rect 2746 2413 2749 2426
rect 2762 2403 2765 2476
rect 2786 2413 2789 2426
rect 2738 2303 2741 2326
rect 2714 2233 2733 2236
rect 2666 2173 2677 2176
rect 2674 2056 2677 2173
rect 2706 2143 2709 2166
rect 2658 2053 2677 2056
rect 2714 2056 2717 2233
rect 2762 2226 2765 2396
rect 2762 2223 2769 2226
rect 2730 2193 2733 2206
rect 2722 2133 2725 2166
rect 2754 2156 2757 2216
rect 2746 2153 2757 2156
rect 2746 2123 2749 2153
rect 2766 2146 2769 2223
rect 2778 2203 2781 2336
rect 2786 2323 2789 2336
rect 2794 2256 2797 2623
rect 2802 2593 2805 2606
rect 2810 2393 2813 2556
rect 2826 2546 2829 2606
rect 2834 2593 2837 2606
rect 2842 2593 2845 2626
rect 2850 2576 2853 2843
rect 2874 2826 2877 2893
rect 2858 2803 2861 2826
rect 2866 2823 2877 2826
rect 2866 2803 2869 2823
rect 2898 2806 2901 2966
rect 2906 2926 2909 2936
rect 2906 2923 2925 2926
rect 2930 2923 2933 2936
rect 2946 2903 2949 2993
rect 2962 2863 2965 2946
rect 2922 2823 2925 2836
rect 2930 2813 2949 2816
rect 2890 2803 2901 2806
rect 2858 2733 2861 2746
rect 2866 2666 2869 2756
rect 2890 2736 2893 2803
rect 2906 2773 2909 2796
rect 2890 2733 2901 2736
rect 2890 2696 2893 2716
rect 2862 2663 2869 2666
rect 2886 2693 2893 2696
rect 2862 2606 2865 2663
rect 2818 2543 2829 2546
rect 2842 2573 2853 2576
rect 2858 2603 2865 2606
rect 2874 2603 2877 2656
rect 2886 2626 2889 2693
rect 2886 2623 2893 2626
rect 2826 2416 2829 2536
rect 2842 2526 2845 2573
rect 2858 2536 2861 2603
rect 2882 2593 2885 2606
rect 2890 2603 2893 2623
rect 2874 2543 2877 2566
rect 2858 2533 2869 2536
rect 2842 2523 2853 2526
rect 2826 2413 2845 2416
rect 2842 2363 2845 2413
rect 2818 2303 2821 2336
rect 2842 2306 2845 2326
rect 2834 2303 2845 2306
rect 2834 2256 2837 2303
rect 2794 2253 2801 2256
rect 2834 2253 2845 2256
rect 2798 2196 2801 2253
rect 2810 2203 2813 2216
rect 2798 2193 2805 2196
rect 2818 2193 2821 2226
rect 2762 2143 2769 2146
rect 2714 2053 2729 2056
rect 2642 2003 2645 2026
rect 2658 1973 2661 2053
rect 2682 2013 2685 2036
rect 2726 2006 2729 2053
rect 2738 2013 2741 2026
rect 2726 2003 2733 2006
rect 2594 1903 2605 1906
rect 2570 1873 2581 1876
rect 2570 1813 2573 1866
rect 2578 1803 2581 1873
rect 2602 1836 2605 1903
rect 2594 1833 2605 1836
rect 2554 1793 2565 1796
rect 2562 1736 2565 1793
rect 2554 1733 2565 1736
rect 2414 1513 2421 1516
rect 2418 1426 2421 1513
rect 2458 1476 2461 1526
rect 2454 1473 2461 1476
rect 2418 1423 2429 1426
rect 2314 1283 2325 1286
rect 2314 1226 2317 1283
rect 2306 1223 2317 1226
rect 2306 1193 2309 1223
rect 2314 1213 2325 1216
rect 2274 1093 2285 1096
rect 2294 1153 2301 1156
rect 2274 1026 2277 1093
rect 2294 1086 2297 1153
rect 2330 1136 2333 1236
rect 2322 1133 2333 1136
rect 2294 1083 2301 1086
rect 2274 1023 2285 1026
rect 2250 963 2253 1006
rect 2258 956 2261 1006
rect 2250 953 2261 956
rect 2250 863 2253 953
rect 2258 923 2261 946
rect 2274 933 2277 1006
rect 2234 853 2245 856
rect 2226 723 2229 816
rect 2234 766 2237 853
rect 2242 783 2245 846
rect 2266 836 2269 856
rect 2262 833 2269 836
rect 2250 773 2253 806
rect 2262 776 2265 833
rect 2274 796 2277 816
rect 2282 813 2285 1023
rect 2298 1013 2301 1083
rect 2322 1066 2325 1133
rect 2330 1113 2333 1126
rect 2314 1063 2325 1066
rect 2314 1023 2317 1063
rect 2338 1036 2341 1326
rect 2362 1323 2365 1346
rect 2378 1343 2389 1346
rect 2346 1203 2349 1226
rect 2354 1213 2357 1246
rect 2362 1133 2365 1146
rect 2378 1143 2381 1343
rect 2386 1333 2397 1336
rect 2410 1333 2413 1416
rect 2426 1336 2429 1423
rect 2454 1386 2457 1473
rect 2454 1383 2461 1386
rect 2418 1333 2429 1336
rect 2386 1096 2389 1116
rect 2378 1093 2389 1096
rect 2378 1036 2381 1093
rect 2394 1086 2397 1326
rect 2410 1203 2413 1226
rect 2418 1216 2421 1333
rect 2434 1233 2437 1316
rect 2418 1213 2429 1216
rect 2402 1093 2405 1156
rect 2410 1133 2413 1186
rect 2426 1146 2429 1213
rect 2458 1163 2461 1383
rect 2466 1333 2469 1626
rect 2530 1623 2533 1726
rect 2538 1613 2541 1726
rect 2546 1613 2549 1716
rect 2554 1713 2557 1733
rect 2586 1713 2589 1726
rect 2578 1693 2581 1706
rect 2594 1626 2597 1833
rect 2618 1796 2621 1816
rect 2626 1803 2629 1836
rect 2634 1813 2637 1926
rect 2674 1913 2677 1926
rect 2690 1886 2693 1976
rect 2714 1913 2717 1926
rect 2690 1883 2709 1886
rect 2690 1813 2693 1826
rect 2634 1796 2637 1806
rect 2706 1803 2709 1883
rect 2618 1793 2637 1796
rect 2602 1703 2605 1736
rect 2586 1623 2597 1626
rect 2498 1566 2501 1606
rect 2498 1563 2509 1566
rect 2474 1323 2477 1536
rect 2482 1523 2485 1546
rect 2506 1533 2509 1563
rect 2522 1543 2525 1606
rect 2546 1603 2557 1606
rect 2586 1566 2589 1623
rect 2586 1563 2597 1566
rect 2482 1403 2485 1516
rect 2538 1433 2541 1546
rect 2546 1533 2549 1546
rect 2594 1543 2597 1563
rect 2602 1523 2605 1616
rect 2634 1513 2637 1526
rect 2594 1416 2597 1436
rect 2490 1306 2493 1396
rect 2498 1316 2501 1336
rect 2554 1323 2557 1336
rect 2498 1313 2509 1316
rect 2482 1303 2493 1306
rect 2482 1213 2485 1303
rect 2506 1256 2509 1313
rect 2578 1306 2581 1416
rect 2498 1253 2509 1256
rect 2570 1303 2581 1306
rect 2590 1413 2597 1416
rect 2590 1306 2593 1413
rect 2602 1383 2605 1456
rect 2642 1453 2645 1706
rect 2650 1533 2653 1706
rect 2658 1613 2661 1726
rect 2690 1713 2693 1726
rect 2706 1713 2709 1776
rect 2698 1693 2701 1706
rect 2714 1703 2717 1716
rect 2722 1693 2725 1706
rect 2698 1636 2701 1656
rect 2730 1653 2733 2003
rect 2762 1936 2765 2143
rect 2778 2063 2781 2136
rect 2778 2013 2781 2026
rect 2778 1943 2781 1996
rect 2754 1933 2765 1936
rect 2754 1886 2757 1933
rect 2762 1923 2773 1926
rect 2786 1906 2789 2136
rect 2794 2003 2797 2126
rect 2802 2106 2805 2193
rect 2826 2183 2829 2236
rect 2842 2213 2845 2253
rect 2842 2183 2845 2206
rect 2802 2103 2813 2106
rect 2810 2046 2813 2103
rect 2802 2043 2813 2046
rect 2802 2006 2805 2043
rect 2802 2003 2813 2006
rect 2746 1883 2757 1886
rect 2778 1903 2789 1906
rect 2738 1813 2741 1826
rect 2746 1696 2749 1883
rect 2778 1856 2781 1903
rect 2778 1853 2789 1856
rect 2786 1813 2789 1853
rect 2794 1803 2797 1926
rect 2810 1836 2813 2003
rect 2834 1893 2837 1936
rect 2802 1833 2813 1836
rect 2802 1813 2805 1833
rect 2834 1816 2837 1846
rect 2842 1823 2845 1926
rect 2826 1813 2837 1816
rect 2754 1713 2757 1726
rect 2794 1723 2797 1796
rect 2826 1756 2829 1813
rect 2842 1793 2845 1806
rect 2850 1773 2853 2523
rect 2866 2406 2869 2533
rect 2890 2523 2893 2536
rect 2890 2503 2893 2516
rect 2898 2486 2901 2733
rect 2906 2716 2909 2736
rect 2914 2733 2917 2806
rect 2930 2803 2933 2813
rect 2946 2763 2949 2806
rect 2954 2803 2957 2836
rect 2970 2823 2973 3316
rect 2994 3256 2997 3323
rect 2986 3253 2997 3256
rect 2986 3203 2989 3253
rect 2978 3063 2981 3136
rect 2986 3116 2989 3136
rect 2986 3113 2997 3116
rect 2994 3046 2997 3113
rect 2986 3043 2997 3046
rect 2986 3023 2989 3043
rect 3018 2996 3021 3206
rect 3034 3203 3037 3326
rect 3050 3313 3053 3336
rect 3026 3133 3029 3146
rect 3034 3123 3037 3136
rect 3034 3093 3037 3116
rect 3010 2993 3021 2996
rect 2906 2713 2913 2716
rect 2910 2636 2913 2713
rect 2906 2633 2913 2636
rect 2906 2613 2909 2633
rect 2914 2533 2917 2586
rect 2922 2546 2925 2726
rect 2930 2713 2933 2726
rect 2922 2543 2933 2546
rect 2906 2523 2917 2526
rect 2922 2503 2925 2536
rect 2930 2513 2933 2543
rect 2954 2526 2957 2746
rect 2962 2733 2965 2806
rect 2970 2723 2973 2736
rect 2970 2703 2973 2716
rect 2994 2713 2997 2826
rect 3010 2723 3013 2993
rect 3034 2923 3037 3016
rect 3058 2963 3061 3526
rect 3074 3516 3077 3613
rect 3082 3603 3085 3736
rect 3090 3726 3093 3743
rect 3098 3733 3101 3806
rect 3122 3803 3125 3833
rect 3122 3736 3125 3756
rect 3130 3743 3133 3826
rect 3138 3803 3149 3806
rect 3162 3796 3165 3973
rect 3170 3933 3173 4026
rect 3186 3956 3189 4033
rect 3210 3976 3213 4073
rect 3178 3953 3189 3956
rect 3202 3973 3213 3976
rect 3178 3923 3181 3953
rect 3202 3916 3205 3973
rect 3226 3923 3229 3986
rect 3234 3933 3237 4016
rect 3202 3913 3213 3916
rect 3210 3856 3213 3913
rect 3242 3903 3245 3926
rect 3250 3856 3253 4113
rect 3258 3933 3261 3966
rect 3298 3946 3301 4263
rect 3314 4193 3317 4216
rect 3338 4123 3349 4126
rect 3330 3983 3333 4016
rect 3298 3943 3309 3946
rect 3274 3903 3277 3936
rect 3306 3896 3309 3943
rect 3322 3923 3325 3956
rect 3202 3853 3213 3856
rect 3242 3853 3253 3856
rect 3298 3893 3309 3896
rect 3146 3793 3165 3796
rect 3106 3733 3117 3736
rect 3122 3733 3133 3736
rect 3090 3723 3109 3726
rect 3090 3613 3101 3616
rect 3070 3513 3077 3516
rect 3070 3446 3073 3513
rect 3070 3443 3077 3446
rect 3074 3376 3077 3443
rect 3070 3373 3077 3376
rect 3082 3376 3085 3516
rect 3098 3513 3101 3606
rect 3106 3593 3109 3606
rect 3122 3603 3125 3716
rect 3130 3603 3133 3636
rect 3146 3563 3149 3793
rect 3170 3733 3173 3796
rect 3186 3746 3189 3806
rect 3202 3793 3205 3853
rect 3226 3803 3229 3816
rect 3242 3776 3245 3853
rect 3242 3773 3253 3776
rect 3186 3743 3205 3746
rect 3194 3686 3197 3726
rect 3186 3683 3197 3686
rect 3178 3613 3181 3676
rect 3186 3603 3189 3683
rect 3194 3613 3197 3636
rect 3202 3596 3205 3743
rect 3186 3593 3205 3596
rect 3234 3593 3237 3606
rect 3106 3533 3109 3546
rect 3098 3383 3101 3406
rect 3146 3403 3149 3416
rect 3082 3373 3101 3376
rect 3070 3316 3073 3373
rect 3098 3356 3101 3373
rect 3098 3353 3109 3356
rect 3070 3313 3077 3316
rect 3074 3293 3077 3313
rect 3066 3213 3085 3216
rect 3074 3006 3077 3206
rect 3090 3203 3093 3326
rect 3106 3296 3109 3353
rect 3138 3333 3141 3386
rect 3098 3293 3109 3296
rect 3090 3123 3093 3136
rect 3074 3003 3085 3006
rect 3042 2873 3045 2956
rect 3050 2906 3053 2936
rect 3058 2933 3061 2946
rect 3058 2923 3069 2926
rect 3050 2903 3061 2906
rect 3058 2836 3061 2903
rect 3034 2723 3037 2816
rect 3042 2803 3045 2836
rect 3050 2833 3061 2836
rect 3050 2813 3053 2833
rect 3058 2806 3061 2816
rect 3050 2803 3061 2806
rect 3066 2793 3069 2806
rect 3074 2803 3077 2826
rect 3082 2803 3085 3003
rect 3098 2816 3101 3293
rect 3106 3166 3109 3276
rect 3114 3203 3117 3216
rect 3122 3183 3125 3206
rect 3106 3163 3125 3166
rect 3122 3026 3125 3163
rect 3114 3023 3125 3026
rect 3114 2906 3117 3023
rect 3138 2923 3141 3006
rect 3106 2903 3117 2906
rect 3106 2883 3109 2903
rect 3146 2853 3149 3286
rect 3154 3276 3157 3346
rect 3162 3283 3165 3536
rect 3186 3486 3189 3593
rect 3178 3483 3189 3486
rect 3178 3436 3181 3483
rect 3178 3433 3189 3436
rect 3154 3273 3165 3276
rect 3162 3213 3165 3273
rect 3162 3173 3165 3206
rect 3170 3203 3173 3406
rect 3178 3333 3181 3416
rect 3178 3203 3181 3266
rect 3186 3203 3189 3433
rect 3194 3376 3197 3516
rect 3202 3503 3205 3526
rect 3218 3503 3221 3556
rect 3226 3523 3237 3526
rect 3242 3433 3245 3626
rect 3210 3383 3213 3406
rect 3194 3373 3201 3376
rect 3198 3256 3201 3373
rect 3242 3336 3245 3416
rect 3194 3253 3201 3256
rect 3194 3233 3197 3253
rect 3194 3196 3197 3216
rect 3178 3193 3197 3196
rect 3178 3133 3181 3193
rect 3186 3133 3189 3186
rect 3202 3133 3205 3206
rect 3210 3183 3213 3336
rect 3234 3333 3245 3336
rect 3250 3333 3253 3773
rect 3298 3756 3301 3893
rect 3338 3836 3341 3926
rect 3330 3833 3341 3836
rect 3314 3813 3317 3826
rect 3330 3786 3333 3833
rect 3330 3783 3341 3786
rect 3338 3766 3341 3783
rect 3338 3763 3345 3766
rect 3294 3753 3301 3756
rect 3282 3673 3285 3726
rect 3294 3706 3297 3753
rect 3294 3703 3301 3706
rect 3258 3633 3261 3646
rect 3258 3613 3261 3626
rect 3274 3623 3277 3646
rect 3258 3423 3261 3536
rect 3274 3456 3277 3616
rect 3282 3493 3285 3516
rect 3290 3513 3293 3526
rect 3274 3453 3281 3456
rect 3278 3406 3281 3453
rect 3298 3426 3301 3703
rect 3314 3566 3317 3746
rect 3342 3696 3345 3763
rect 3354 3743 3357 4176
rect 3362 4153 3365 4206
rect 3378 4136 3381 4516
rect 3434 4513 3437 4526
rect 3482 4513 3485 4526
rect 3490 4506 3493 4526
rect 3506 4513 3509 4526
rect 3522 4506 3525 4526
rect 3394 4483 3397 4506
rect 3490 4503 3525 4506
rect 3546 4483 3549 4546
rect 3570 4533 3573 4586
rect 3594 4576 3597 4596
rect 3602 4583 3605 4616
rect 3594 4573 3605 4576
rect 3562 4486 3565 4526
rect 3578 4523 3581 4546
rect 3562 4483 3573 4486
rect 3418 4433 3421 4466
rect 3402 4256 3405 4426
rect 3442 4423 3445 4456
rect 3426 4383 3429 4416
rect 3418 4333 3429 4336
rect 3434 4333 3437 4396
rect 3450 4346 3453 4416
rect 3506 4393 3509 4416
rect 3530 4346 3533 4436
rect 3450 4343 3461 4346
rect 3410 4323 3429 4326
rect 3398 4253 3405 4256
rect 3370 4133 3381 4136
rect 3370 3866 3373 4133
rect 3386 4036 3389 4226
rect 3398 4206 3401 4253
rect 3410 4233 3413 4246
rect 3426 4226 3429 4323
rect 3450 4233 3453 4336
rect 3458 4333 3461 4343
rect 3510 4343 3533 4346
rect 3458 4243 3469 4246
rect 3410 4213 3413 4226
rect 3426 4223 3437 4226
rect 3458 4223 3461 4243
rect 3398 4203 3405 4206
rect 3394 4103 3397 4126
rect 3382 4033 3389 4036
rect 3382 3916 3385 4033
rect 3394 4003 3397 4026
rect 3394 3923 3397 3976
rect 3402 3923 3405 4203
rect 3426 4123 3429 4216
rect 3434 4203 3437 4223
rect 3410 4013 3413 4116
rect 3418 4083 3421 4106
rect 3410 3916 3413 4006
rect 3418 3973 3421 4016
rect 3426 3953 3429 4006
rect 3418 3923 3421 3936
rect 3382 3913 3389 3916
rect 3370 3863 3381 3866
rect 3362 3713 3365 3726
rect 3338 3693 3345 3696
rect 3338 3613 3341 3693
rect 3378 3676 3381 3863
rect 3370 3673 3381 3676
rect 3370 3616 3373 3673
rect 3370 3613 3377 3616
rect 3314 3563 3325 3566
rect 3298 3423 3305 3426
rect 3274 3403 3281 3406
rect 3226 3313 3229 3326
rect 3242 3263 3245 3326
rect 3258 3313 3261 3326
rect 3178 3123 3197 3126
rect 3210 3123 3213 3176
rect 3218 3133 3221 3196
rect 3226 3106 3229 3186
rect 3234 3166 3237 3236
rect 3250 3203 3253 3216
rect 3258 3186 3261 3296
rect 3254 3183 3261 3186
rect 3234 3163 3245 3166
rect 3218 3103 3229 3106
rect 3218 3036 3221 3103
rect 3242 3096 3245 3163
rect 3254 3106 3257 3183
rect 3266 3113 3269 3336
rect 3254 3103 3261 3106
rect 3234 3093 3245 3096
rect 3234 3046 3237 3093
rect 3234 3043 3241 3046
rect 3218 3033 3229 3036
rect 3170 2923 3173 2946
rect 3170 2836 3173 2856
rect 3166 2833 3173 2836
rect 3094 2813 3101 2816
rect 3058 2733 3061 2746
rect 3066 2733 3069 2786
rect 3094 2746 3097 2813
rect 3094 2743 3101 2746
rect 2970 2593 2973 2606
rect 2986 2536 2989 2666
rect 3050 2656 3053 2726
rect 3074 2713 3077 2726
rect 3074 2686 3077 2706
rect 3070 2683 3077 2686
rect 3050 2653 3061 2656
rect 3034 2613 3037 2646
rect 3034 2576 3037 2606
rect 3034 2573 3045 2576
rect 2986 2533 2997 2536
rect 3034 2533 3037 2546
rect 3042 2533 3045 2573
rect 3058 2566 3061 2653
rect 3070 2636 3073 2683
rect 3082 2643 3085 2736
rect 3070 2633 3077 2636
rect 3050 2563 3061 2566
rect 2954 2523 2981 2526
rect 2898 2483 2917 2486
rect 2866 2403 2873 2406
rect 2858 2373 2861 2396
rect 2870 2356 2873 2403
rect 2882 2393 2885 2406
rect 2866 2353 2873 2356
rect 2866 2323 2869 2353
rect 2890 2333 2893 2416
rect 2914 2336 2917 2483
rect 2954 2456 2957 2516
rect 2950 2453 2957 2456
rect 2970 2456 2973 2523
rect 2994 2466 2997 2533
rect 2986 2463 2997 2466
rect 2970 2453 2977 2456
rect 2938 2393 2941 2416
rect 2950 2376 2953 2453
rect 2974 2376 2977 2453
rect 2950 2373 2957 2376
rect 2898 2333 2917 2336
rect 2898 2316 2901 2333
rect 2858 2296 2861 2316
rect 2890 2313 2901 2316
rect 2858 2293 2869 2296
rect 2866 2226 2869 2293
rect 2890 2246 2893 2313
rect 2890 2243 2901 2246
rect 2858 2223 2869 2226
rect 2858 2203 2861 2223
rect 2890 2206 2893 2226
rect 2882 2203 2893 2206
rect 2882 2156 2885 2203
rect 2882 2153 2893 2156
rect 2882 2113 2885 2136
rect 2890 2006 2893 2153
rect 2882 2003 2893 2006
rect 2882 1956 2885 2003
rect 2898 1996 2901 2243
rect 2906 2223 2909 2306
rect 2922 2143 2925 2156
rect 2906 2133 2917 2136
rect 2906 2106 2909 2126
rect 2930 2123 2933 2316
rect 2954 2303 2957 2373
rect 2970 2373 2977 2376
rect 2970 2313 2973 2373
rect 2986 2253 2989 2463
rect 2994 2413 2997 2426
rect 3018 2376 3021 2526
rect 3050 2473 3053 2563
rect 3058 2503 3061 2536
rect 3066 2493 3069 2546
rect 3074 2533 3077 2633
rect 3090 2593 3093 2726
rect 3034 2393 3037 2406
rect 3010 2373 3021 2376
rect 3010 2276 3013 2373
rect 3042 2346 3045 2416
rect 3050 2413 3069 2416
rect 3058 2346 3061 2406
rect 3074 2403 3077 2426
rect 3034 2343 3045 2346
rect 3050 2343 3061 2346
rect 3034 2333 3037 2343
rect 3050 2336 3053 2343
rect 3042 2333 3053 2336
rect 3002 2273 3013 2276
rect 2978 2226 2981 2246
rect 2970 2223 2981 2226
rect 2970 2156 2973 2223
rect 2986 2193 2989 2206
rect 2970 2153 2981 2156
rect 2906 2103 2917 2106
rect 2914 2036 2917 2103
rect 2970 2083 2973 2136
rect 2978 2133 2981 2153
rect 2978 2113 2981 2126
rect 2994 2066 2997 2146
rect 2906 2033 2917 2036
rect 2986 2063 2997 2066
rect 2906 2016 2909 2033
rect 2906 2013 2917 2016
rect 2898 1993 2905 1996
rect 2882 1953 2893 1956
rect 2858 1813 2861 1926
rect 2866 1923 2869 1936
rect 2866 1896 2869 1916
rect 2890 1913 2893 1953
rect 2902 1906 2905 1993
rect 2898 1903 2905 1906
rect 2914 1906 2917 2013
rect 2946 1933 2949 1976
rect 2954 1923 2957 2006
rect 2986 1976 2989 2063
rect 2986 1973 2997 1976
rect 2914 1903 2925 1906
rect 2866 1893 2877 1896
rect 2874 1836 2877 1893
rect 2866 1833 2877 1836
rect 2866 1813 2869 1833
rect 2874 1793 2877 1806
rect 2826 1753 2837 1756
rect 2802 1716 2805 1726
rect 2810 1723 2813 1736
rect 2802 1713 2829 1716
rect 2746 1693 2757 1696
rect 2754 1646 2757 1693
rect 2746 1643 2757 1646
rect 2698 1633 2705 1636
rect 2682 1583 2685 1606
rect 2702 1586 2705 1633
rect 2698 1583 2705 1586
rect 2682 1506 2685 1526
rect 2674 1503 2685 1506
rect 2674 1456 2677 1503
rect 2698 1456 2701 1583
rect 2714 1566 2717 1606
rect 2746 1593 2749 1643
rect 2802 1613 2805 1713
rect 2834 1696 2837 1753
rect 2842 1726 2845 1746
rect 2842 1723 2853 1726
rect 2826 1693 2837 1696
rect 2826 1596 2829 1693
rect 2850 1676 2853 1723
rect 2842 1673 2853 1676
rect 2842 1626 2845 1673
rect 2842 1623 2853 1626
rect 2850 1603 2853 1623
rect 2826 1593 2837 1596
rect 2710 1563 2717 1566
rect 2710 1486 2713 1563
rect 2746 1536 2749 1586
rect 2738 1533 2749 1536
rect 2778 1533 2781 1586
rect 2834 1563 2837 1593
rect 2710 1483 2717 1486
rect 2674 1453 2681 1456
rect 2698 1453 2705 1456
rect 2626 1413 2629 1426
rect 2634 1413 2637 1436
rect 2658 1413 2661 1426
rect 2602 1313 2605 1336
rect 2610 1323 2613 1406
rect 2658 1393 2661 1406
rect 2590 1303 2597 1306
rect 2498 1236 2501 1253
rect 2490 1233 2501 1236
rect 2570 1236 2573 1303
rect 2570 1233 2581 1236
rect 2490 1153 2493 1233
rect 2506 1213 2509 1226
rect 2418 1143 2429 1146
rect 2394 1083 2405 1086
rect 2418 1083 2421 1143
rect 2522 1126 2525 1146
rect 2538 1133 2541 1216
rect 2578 1213 2581 1233
rect 2546 1133 2549 1146
rect 2426 1113 2429 1126
rect 2434 1103 2437 1126
rect 2522 1123 2533 1126
rect 2330 1033 2341 1036
rect 2290 923 2293 966
rect 2314 946 2317 1006
rect 2330 966 2333 1033
rect 2330 963 2341 966
rect 2306 943 2317 946
rect 2306 906 2309 926
rect 2298 903 2309 906
rect 2298 846 2301 903
rect 2298 843 2309 846
rect 2314 843 2317 936
rect 2306 823 2309 843
rect 2274 793 2281 796
rect 2262 773 2269 776
rect 2234 763 2241 766
rect 2238 716 2241 763
rect 2234 713 2241 716
rect 2234 643 2237 713
rect 2266 686 2269 773
rect 2278 726 2281 793
rect 2274 723 2281 726
rect 2290 723 2293 806
rect 2322 756 2325 946
rect 2330 813 2333 916
rect 2338 853 2341 963
rect 2346 943 2349 1026
rect 2346 846 2349 936
rect 2354 913 2357 1036
rect 2378 1033 2389 1036
rect 2362 953 2365 1006
rect 2378 1005 2381 1016
rect 2386 1003 2389 1033
rect 2402 1013 2405 1083
rect 2450 1003 2453 1036
rect 2450 906 2453 926
rect 2338 843 2349 846
rect 2338 813 2341 843
rect 2354 836 2357 906
rect 2442 903 2453 906
rect 2442 846 2445 903
rect 2442 843 2453 846
rect 2346 833 2357 836
rect 2346 813 2349 833
rect 2450 816 2453 843
rect 2330 803 2341 806
rect 2354 756 2357 816
rect 2442 813 2453 816
rect 2442 793 2445 813
rect 2450 793 2453 806
rect 2322 753 2333 756
rect 2274 703 2277 723
rect 2206 563 2213 566
rect 2226 566 2229 616
rect 2226 563 2233 566
rect 2182 483 2189 486
rect 2126 443 2133 446
rect 2126 396 2129 443
rect 2170 413 2173 456
rect 2182 416 2185 483
rect 2182 413 2189 416
rect 2126 393 2133 396
rect 2154 393 2157 406
rect 2130 323 2133 393
rect 2146 276 2149 356
rect 2178 333 2181 396
rect 2186 353 2189 413
rect 2194 356 2197 526
rect 2206 486 2209 563
rect 2230 486 2233 563
rect 2242 523 2245 566
rect 2250 496 2253 686
rect 2266 683 2285 686
rect 2282 576 2285 683
rect 2314 616 2317 746
rect 2330 726 2333 753
rect 2346 753 2357 756
rect 2346 733 2349 753
rect 2354 743 2365 746
rect 2458 743 2461 816
rect 2466 803 2469 1096
rect 2474 1086 2477 1106
rect 2474 1083 2485 1086
rect 2482 976 2485 1083
rect 2498 1066 2501 1086
rect 2474 973 2485 976
rect 2494 1063 2501 1066
rect 2474 906 2477 973
rect 2482 923 2485 956
rect 2494 936 2497 1063
rect 2506 1013 2509 1106
rect 2530 1103 2533 1123
rect 2554 1036 2557 1126
rect 2570 1123 2573 1196
rect 2578 1183 2581 1206
rect 2586 1123 2589 1226
rect 2546 1033 2557 1036
rect 2522 1013 2541 1016
rect 2546 1013 2549 1033
rect 2506 946 2509 1006
rect 2514 963 2517 1006
rect 2506 943 2517 946
rect 2494 933 2501 936
rect 2474 903 2485 906
rect 2482 836 2485 903
rect 2474 833 2485 836
rect 2474 793 2477 833
rect 2482 803 2485 816
rect 2466 733 2469 786
rect 2474 726 2477 736
rect 2490 733 2493 816
rect 2330 723 2349 726
rect 2330 623 2333 636
rect 2314 613 2321 616
rect 2266 573 2285 576
rect 2266 556 2269 573
rect 2258 553 2269 556
rect 2258 506 2261 553
rect 2274 533 2277 546
rect 2306 523 2309 606
rect 2318 566 2321 613
rect 2346 603 2349 723
rect 2354 613 2357 636
rect 2378 623 2381 706
rect 2394 606 2397 646
rect 2354 593 2357 606
rect 2314 563 2321 566
rect 2314 543 2317 563
rect 2362 523 2365 606
rect 2370 523 2373 606
rect 2386 603 2397 606
rect 2258 503 2277 506
rect 2250 493 2261 496
rect 2206 483 2213 486
rect 2210 456 2213 483
rect 2226 483 2233 486
rect 2210 453 2217 456
rect 2194 353 2205 356
rect 2194 333 2197 346
rect 2154 313 2157 326
rect 2138 273 2149 276
rect 2138 176 2141 273
rect 2162 176 2165 296
rect 2138 173 2149 176
rect 2130 133 2133 146
rect 2090 113 2097 116
rect 2090 93 2093 113
rect 2146 106 2149 173
rect 2130 103 2149 106
rect 2154 173 2165 176
rect 2074 83 2085 86
rect 2074 0 2077 83
rect 2090 0 2093 86
rect 2114 0 2117 96
rect 2130 0 2133 103
rect 2154 0 2157 173
rect 2162 93 2165 156
rect 2170 33 2173 216
rect 2178 26 2181 326
rect 2194 313 2197 326
rect 2202 306 2205 353
rect 2214 316 2217 453
rect 2226 426 2229 483
rect 2226 423 2237 426
rect 2186 303 2205 306
rect 2210 313 2217 316
rect 2186 196 2189 303
rect 2210 293 2213 313
rect 2186 193 2197 196
rect 2210 193 2213 206
rect 2194 166 2197 193
rect 2194 163 2205 166
rect 2202 86 2205 163
rect 2226 143 2229 416
rect 2234 313 2237 423
rect 2258 393 2261 493
rect 2242 323 2245 386
rect 2274 366 2277 503
rect 2386 446 2389 603
rect 2402 583 2405 606
rect 2282 413 2285 446
rect 2386 443 2397 446
rect 2270 363 2277 366
rect 2234 213 2237 306
rect 2258 256 2261 316
rect 2270 286 2273 363
rect 2338 333 2341 396
rect 2346 356 2349 416
rect 2370 393 2373 406
rect 2370 366 2373 386
rect 2346 353 2357 356
rect 2270 283 2277 286
rect 2254 253 2261 256
rect 2242 133 2245 196
rect 2254 176 2257 253
rect 2274 203 2277 283
rect 2290 246 2293 326
rect 2354 296 2357 353
rect 2362 323 2365 366
rect 2370 363 2377 366
rect 2386 363 2389 396
rect 2286 243 2293 246
rect 2346 293 2357 296
rect 2254 173 2261 176
rect 2258 156 2261 173
rect 2286 166 2289 243
rect 2298 173 2301 216
rect 2322 193 2325 206
rect 2346 176 2349 293
rect 2362 213 2365 316
rect 2374 206 2377 363
rect 2394 256 2397 443
rect 2402 313 2405 536
rect 2410 413 2413 626
rect 2418 506 2421 706
rect 2426 583 2429 616
rect 2442 613 2445 726
rect 2466 723 2477 726
rect 2426 533 2429 576
rect 2450 556 2453 616
rect 2466 603 2469 723
rect 2498 703 2501 933
rect 2514 766 2517 943
rect 2530 913 2533 936
rect 2538 923 2541 1013
rect 2594 1003 2597 1303
rect 2602 1203 2605 1236
rect 2626 1233 2629 1326
rect 2626 1213 2629 1226
rect 2634 1213 2637 1386
rect 2666 1323 2669 1436
rect 2678 1356 2681 1453
rect 2702 1396 2705 1453
rect 2698 1393 2705 1396
rect 2698 1376 2701 1393
rect 2690 1373 2701 1376
rect 2678 1353 2685 1356
rect 2602 1116 2605 1196
rect 2610 1123 2613 1186
rect 2618 1123 2621 1176
rect 2626 1123 2629 1166
rect 2602 1113 2609 1116
rect 2634 1113 2637 1126
rect 2606 1036 2609 1113
rect 2618 1046 2621 1106
rect 2618 1043 2625 1046
rect 2606 1033 2613 1036
rect 2602 1003 2605 1016
rect 2586 933 2589 986
rect 2530 813 2533 836
rect 2538 803 2541 826
rect 2506 763 2517 766
rect 2554 766 2557 896
rect 2562 813 2565 826
rect 2554 763 2581 766
rect 2506 686 2509 763
rect 2522 736 2525 746
rect 2502 683 2509 686
rect 2514 733 2525 736
rect 2474 613 2485 616
rect 2474 593 2477 613
rect 2490 606 2493 616
rect 2482 603 2493 606
rect 2482 593 2485 603
rect 2434 553 2453 556
rect 2434 523 2437 553
rect 2490 533 2493 586
rect 2502 516 2505 683
rect 2514 523 2517 733
rect 2522 713 2525 726
rect 2554 703 2557 726
rect 2570 723 2573 736
rect 2502 513 2509 516
rect 2418 503 2429 506
rect 2426 446 2429 503
rect 2418 443 2429 446
rect 2410 303 2413 326
rect 2394 253 2401 256
rect 2286 163 2293 166
rect 2258 153 2265 156
rect 2170 23 2181 26
rect 2194 83 2205 86
rect 2170 0 2173 23
rect 2194 0 2197 83
rect 2218 66 2221 126
rect 2210 63 2221 66
rect 2210 0 2213 63
rect 2226 0 2229 36
rect 2242 0 2245 126
rect 2262 106 2265 153
rect 2290 143 2293 163
rect 2330 156 2333 176
rect 2346 173 2357 176
rect 2330 153 2337 156
rect 2290 123 2293 136
rect 2258 103 2265 106
rect 2258 0 2261 103
rect 2274 76 2277 116
rect 2314 113 2317 126
rect 2322 106 2325 146
rect 2314 103 2325 106
rect 2314 76 2317 103
rect 2334 96 2337 153
rect 2274 73 2285 76
rect 2282 16 2285 73
rect 2274 13 2285 16
rect 2306 73 2317 76
rect 2330 93 2337 96
rect 2306 16 2309 73
rect 2306 13 2317 16
rect 2274 0 2277 13
rect 2314 0 2317 13
rect 2330 0 2333 93
rect 2354 86 2357 173
rect 2362 106 2365 206
rect 2370 203 2377 206
rect 2370 123 2373 203
rect 2398 176 2401 253
rect 2410 213 2413 226
rect 2394 173 2401 176
rect 2394 113 2397 173
rect 2362 103 2373 106
rect 2346 83 2357 86
rect 2346 0 2349 83
rect 2370 16 2373 103
rect 2418 93 2421 443
rect 2434 376 2437 406
rect 2434 373 2445 376
rect 2442 193 2445 373
rect 2466 323 2469 416
rect 2506 383 2509 513
rect 2522 496 2525 616
rect 2538 603 2541 626
rect 2578 613 2581 763
rect 2586 723 2589 926
rect 2610 893 2613 1033
rect 2622 886 2625 1043
rect 2634 1003 2637 1016
rect 2634 913 2637 926
rect 2642 923 2645 1126
rect 2650 1103 2653 1226
rect 2658 1163 2661 1216
rect 2666 1166 2669 1256
rect 2674 1193 2677 1336
rect 2682 1253 2685 1353
rect 2690 1296 2693 1373
rect 2714 1346 2717 1483
rect 2738 1476 2741 1533
rect 2754 1486 2757 1526
rect 2754 1483 2765 1486
rect 2858 1483 2861 1766
rect 2866 1706 2869 1746
rect 2882 1733 2885 1816
rect 2898 1763 2901 1903
rect 2922 1856 2925 1903
rect 2914 1853 2925 1856
rect 2994 1853 2997 1973
rect 3002 1953 3005 2273
rect 3050 2266 3053 2326
rect 3042 2263 3053 2266
rect 3010 2106 3013 2126
rect 3018 2123 3021 2196
rect 3042 2193 3045 2263
rect 3058 2256 3061 2336
rect 3066 2306 3069 2326
rect 3082 2323 3085 2476
rect 3090 2403 3093 2516
rect 3090 2333 3093 2356
rect 3098 2306 3101 2743
rect 3106 2703 3109 2806
rect 3130 2746 3133 2806
rect 3154 2793 3157 2816
rect 3122 2743 3133 2746
rect 3106 2593 3109 2616
rect 3122 2593 3125 2743
rect 3138 2723 3141 2746
rect 3146 2613 3149 2736
rect 3166 2726 3169 2833
rect 3178 2733 3181 2896
rect 3218 2876 3221 3016
rect 3226 3003 3229 3033
rect 3238 2996 3241 3043
rect 3234 2993 3241 2996
rect 3234 2956 3237 2993
rect 3234 2953 3241 2956
rect 3238 2906 3241 2953
rect 3210 2873 3221 2876
rect 3234 2903 3241 2906
rect 3210 2796 3213 2873
rect 3210 2793 3221 2796
rect 3194 2756 3197 2776
rect 3218 2773 3221 2793
rect 3234 2766 3237 2903
rect 3190 2753 3197 2756
rect 3230 2763 3237 2766
rect 3250 2766 3253 3056
rect 3258 2943 3261 3103
rect 3274 3096 3277 3403
rect 3282 3316 3285 3386
rect 3290 3333 3293 3416
rect 3302 3376 3305 3423
rect 3322 3403 3325 3563
rect 3330 3533 3333 3546
rect 3338 3513 3341 3526
rect 3346 3413 3349 3536
rect 3354 3523 3357 3536
rect 3362 3533 3365 3596
rect 3302 3373 3309 3376
rect 3282 3313 3289 3316
rect 3286 3256 3289 3313
rect 3306 3306 3309 3373
rect 3298 3303 3309 3306
rect 3298 3263 3301 3303
rect 3322 3266 3325 3286
rect 3318 3263 3325 3266
rect 3286 3253 3301 3256
rect 3270 3093 3277 3096
rect 3270 3026 3273 3093
rect 3270 3023 3277 3026
rect 3266 2933 3269 3006
rect 3274 2973 3277 3023
rect 3282 3013 3285 3136
rect 3290 3133 3293 3166
rect 3298 3126 3301 3253
rect 3318 3136 3321 3263
rect 3290 3123 3301 3126
rect 3314 3133 3321 3136
rect 3290 3013 3293 3123
rect 3290 2993 3293 3006
rect 3274 2833 3277 2926
rect 3282 2846 3285 2936
rect 3298 2923 3301 3116
rect 3306 2923 3309 3006
rect 3282 2843 3293 2846
rect 3290 2826 3293 2843
rect 3298 2833 3301 2846
rect 3258 2813 3261 2826
rect 3250 2763 3257 2766
rect 3154 2713 3157 2726
rect 3162 2723 3169 2726
rect 3162 2606 3165 2723
rect 3190 2686 3193 2753
rect 3202 2706 3205 2736
rect 3210 2723 3213 2746
rect 3202 2703 3209 2706
rect 3190 2683 3197 2686
rect 3158 2603 3165 2606
rect 3158 2546 3161 2603
rect 3158 2543 3165 2546
rect 3106 2516 3109 2536
rect 3130 2523 3133 2536
rect 3106 2513 3113 2516
rect 3110 2426 3113 2513
rect 3154 2503 3157 2526
rect 3122 2456 3125 2476
rect 3162 2473 3165 2543
rect 3122 2453 3133 2456
rect 3106 2423 3113 2426
rect 3106 2376 3109 2423
rect 3106 2373 3117 2376
rect 3066 2303 3077 2306
rect 3050 2253 3061 2256
rect 3050 2213 3053 2253
rect 3074 2236 3077 2303
rect 3066 2233 3077 2236
rect 3090 2303 3101 2306
rect 3090 2236 3093 2303
rect 3106 2243 3109 2336
rect 3090 2233 3101 2236
rect 3066 2166 3069 2233
rect 3058 2163 3069 2166
rect 3010 2103 3021 2106
rect 3018 2036 3021 2103
rect 3058 2046 3061 2163
rect 3082 2133 3085 2216
rect 3098 2143 3101 2233
rect 3058 2043 3069 2046
rect 3010 2033 3021 2036
rect 3010 1993 3013 2033
rect 3066 2023 3069 2043
rect 3074 2016 3077 2096
rect 3026 2013 3045 2016
rect 3066 2013 3077 2016
rect 3082 2013 3085 2026
rect 3010 1923 3013 1946
rect 3034 1933 3037 1956
rect 3050 1943 3053 2006
rect 3066 2003 3069 2013
rect 3074 1993 3077 2006
rect 3074 1933 3077 1956
rect 2914 1823 2917 1853
rect 2906 1756 2909 1816
rect 2898 1753 2909 1756
rect 2874 1723 2893 1726
rect 2866 1703 2877 1706
rect 2874 1656 2877 1703
rect 2898 1696 2901 1753
rect 2922 1733 2925 1836
rect 2994 1823 2997 1836
rect 2978 1813 2997 1816
rect 2970 1793 2973 1806
rect 2930 1733 2933 1756
rect 2978 1733 2981 1746
rect 2986 1733 2989 1756
rect 2906 1723 2925 1726
rect 2906 1703 2909 1723
rect 2978 1713 2981 1726
rect 2994 1723 2997 1813
rect 3002 1713 3005 1746
rect 3010 1743 3013 1756
rect 2898 1693 2909 1696
rect 2866 1653 2877 1656
rect 2866 1633 2869 1653
rect 2898 1616 2901 1636
rect 2890 1613 2901 1616
rect 2890 1556 2893 1613
rect 2890 1553 2901 1556
rect 2898 1533 2901 1553
rect 2906 1523 2909 1693
rect 2738 1473 2749 1476
rect 2722 1413 2725 1426
rect 2746 1383 2749 1473
rect 2762 1413 2765 1483
rect 2762 1393 2765 1406
rect 2714 1343 2725 1346
rect 2698 1313 2701 1326
rect 2690 1293 2697 1296
rect 2694 1176 2697 1293
rect 2690 1173 2697 1176
rect 2706 1173 2709 1336
rect 2722 1266 2725 1343
rect 2714 1263 2725 1266
rect 2714 1223 2717 1263
rect 2714 1203 2717 1216
rect 2666 1163 2677 1166
rect 2674 1086 2677 1163
rect 2690 1113 2693 1173
rect 2738 1156 2741 1326
rect 2754 1203 2757 1246
rect 2770 1213 2773 1246
rect 2786 1233 2789 1416
rect 2826 1333 2829 1386
rect 2850 1366 2853 1396
rect 2874 1393 2877 1406
rect 2842 1363 2853 1366
rect 2802 1313 2805 1326
rect 2842 1243 2845 1363
rect 2882 1356 2885 1446
rect 2890 1403 2893 1506
rect 2922 1443 2925 1526
rect 2930 1513 2933 1626
rect 3010 1613 3013 1626
rect 3018 1613 3021 1716
rect 3026 1633 3029 1736
rect 3034 1723 3037 1746
rect 3042 1733 3045 1806
rect 3066 1803 3069 1836
rect 3098 1793 3101 2006
rect 3114 2003 3117 2373
rect 3130 2356 3133 2453
rect 3122 2353 3133 2356
rect 3122 2233 3125 2353
rect 3146 2323 3149 2336
rect 3162 2333 3165 2426
rect 3170 2403 3173 2596
rect 3186 2576 3189 2666
rect 3178 2573 3189 2576
rect 3178 2423 3181 2573
rect 3194 2523 3197 2683
rect 3206 2636 3209 2703
rect 3202 2633 3209 2636
rect 3202 2613 3205 2633
rect 3218 2613 3221 2716
rect 3230 2646 3233 2763
rect 3230 2643 3237 2646
rect 3210 2553 3213 2606
rect 3226 2603 3229 2626
rect 3234 2596 3237 2643
rect 3226 2593 3237 2596
rect 3226 2506 3229 2593
rect 3242 2536 3245 2756
rect 3254 2686 3257 2763
rect 3266 2753 3269 2826
rect 3282 2823 3293 2826
rect 3282 2806 3285 2823
rect 3290 2813 3301 2816
rect 3282 2803 3301 2806
rect 3274 2733 3277 2776
rect 3298 2723 3301 2803
rect 3314 2756 3317 3133
rect 3330 3036 3333 3316
rect 3338 3303 3341 3396
rect 3346 3313 3349 3326
rect 3362 3283 3365 3526
rect 3374 3476 3377 3613
rect 3374 3473 3381 3476
rect 3378 3456 3381 3473
rect 3386 3466 3389 3913
rect 3394 3793 3397 3816
rect 3394 3603 3397 3726
rect 3402 3516 3405 3916
rect 3410 3913 3421 3916
rect 3410 3863 3413 3906
rect 3418 3896 3421 3913
rect 3418 3893 3425 3896
rect 3422 3836 3425 3893
rect 3434 3863 3437 4136
rect 3442 4113 3445 4206
rect 3466 4193 3469 4216
rect 3474 4213 3485 4216
rect 3490 4206 3493 4326
rect 3498 4213 3501 4336
rect 3510 4236 3513 4343
rect 3530 4333 3541 4336
rect 3546 4333 3549 4396
rect 3506 4233 3513 4236
rect 3522 4323 3541 4326
rect 3482 4203 3493 4206
rect 3450 4053 3453 4146
rect 3482 4133 3485 4203
rect 3466 4103 3469 4126
rect 3482 4086 3485 4126
rect 3474 4083 3485 4086
rect 3490 4086 3493 4196
rect 3498 4153 3501 4206
rect 3506 4143 3509 4233
rect 3498 4126 3501 4136
rect 3498 4123 3509 4126
rect 3506 4103 3509 4123
rect 3490 4083 3501 4086
rect 3474 4036 3477 4083
rect 3474 4033 3485 4036
rect 3442 3993 3445 4006
rect 3450 3976 3453 4016
rect 3446 3973 3453 3976
rect 3446 3836 3449 3973
rect 3458 3883 3461 4016
rect 3482 4013 3485 4033
rect 3498 3996 3501 4083
rect 3514 4023 3517 4216
rect 3522 4203 3525 4323
rect 3522 4073 3525 4136
rect 3530 4123 3533 4236
rect 3538 4213 3541 4316
rect 3554 4213 3557 4226
rect 3538 4166 3541 4186
rect 3538 4163 3549 4166
rect 3546 4116 3549 4163
rect 3538 4113 3549 4116
rect 3562 4116 3565 4326
rect 3570 4323 3573 4483
rect 3586 4473 3589 4556
rect 3602 4346 3605 4573
rect 3618 4513 3621 4536
rect 3650 4533 3653 4556
rect 3658 4533 3661 4546
rect 3674 4533 3677 4616
rect 3626 4493 3629 4526
rect 3642 4503 3645 4526
rect 3626 4396 3629 4416
rect 3618 4393 3629 4396
rect 3594 4343 3605 4346
rect 3570 4193 3573 4216
rect 3578 4213 3581 4286
rect 3570 4133 3573 4146
rect 3578 4123 3581 4156
rect 3562 4113 3573 4116
rect 3538 4046 3541 4113
rect 3530 4043 3541 4046
rect 3570 4046 3573 4113
rect 3570 4043 3581 4046
rect 3482 3993 3501 3996
rect 3530 3996 3533 4043
rect 3546 4003 3549 4036
rect 3554 4003 3557 4016
rect 3530 3993 3541 3996
rect 3474 3933 3477 3976
rect 3474 3893 3477 3916
rect 3418 3833 3425 3836
rect 3434 3833 3449 3836
rect 3418 3736 3421 3833
rect 3434 3756 3437 3833
rect 3450 3813 3453 3826
rect 3434 3753 3441 3756
rect 3418 3733 3429 3736
rect 3410 3706 3413 3726
rect 3410 3703 3417 3706
rect 3414 3636 3417 3703
rect 3410 3633 3417 3636
rect 3410 3533 3413 3633
rect 3418 3533 3421 3616
rect 3426 3543 3429 3733
rect 3438 3606 3441 3753
rect 3450 3613 3453 3806
rect 3458 3726 3461 3866
rect 3482 3836 3485 3993
rect 3498 3923 3501 3936
rect 3482 3833 3501 3836
rect 3466 3793 3469 3806
rect 3474 3733 3477 3816
rect 3482 3803 3485 3816
rect 3490 3803 3493 3826
rect 3498 3736 3501 3833
rect 3514 3826 3517 3926
rect 3514 3823 3525 3826
rect 3506 3803 3509 3816
rect 3494 3733 3501 3736
rect 3458 3723 3485 3726
rect 3438 3603 3445 3606
rect 3458 3603 3461 3616
rect 3466 3603 3469 3716
rect 3482 3636 3485 3723
rect 3474 3633 3485 3636
rect 3418 3523 3429 3526
rect 3442 3516 3445 3603
rect 3450 3533 3453 3556
rect 3474 3533 3477 3633
rect 3494 3626 3497 3733
rect 3494 3623 3501 3626
rect 3506 3623 3509 3726
rect 3490 3573 3493 3606
rect 3498 3556 3501 3623
rect 3494 3553 3501 3556
rect 3402 3513 3421 3516
rect 3386 3463 3405 3466
rect 3378 3453 3389 3456
rect 3386 3333 3389 3453
rect 3402 3366 3405 3463
rect 3394 3363 3405 3366
rect 3418 3366 3421 3513
rect 3418 3363 3429 3366
rect 3394 3346 3397 3363
rect 3394 3343 3405 3346
rect 3338 3213 3341 3226
rect 3346 3166 3349 3236
rect 3354 3223 3357 3266
rect 3354 3213 3365 3216
rect 3342 3163 3349 3166
rect 3342 3056 3345 3163
rect 3378 3156 3381 3326
rect 3394 3303 3397 3316
rect 3402 3236 3405 3343
rect 3410 3333 3413 3346
rect 3418 3313 3421 3326
rect 3394 3233 3405 3236
rect 3418 3233 3421 3246
rect 3394 3176 3397 3233
rect 3394 3173 3405 3176
rect 3354 3153 3381 3156
rect 3354 3096 3357 3153
rect 3362 3123 3365 3136
rect 3354 3093 3365 3096
rect 3322 3033 3333 3036
rect 3338 3053 3345 3056
rect 3338 3033 3341 3053
rect 3362 3046 3365 3093
rect 3378 3053 3381 3146
rect 3402 3056 3405 3173
rect 3410 3133 3413 3226
rect 3410 3083 3413 3126
rect 3402 3053 3409 3056
rect 3362 3043 3381 3046
rect 3322 2986 3325 3033
rect 3338 3003 3341 3016
rect 3362 2993 3365 3016
rect 3322 2983 3341 2986
rect 3322 2933 3325 2946
rect 3330 2823 3333 2976
rect 3338 2966 3341 2983
rect 3338 2963 3349 2966
rect 3346 2856 3349 2963
rect 3338 2853 3349 2856
rect 3314 2753 3321 2756
rect 3306 2716 3309 2746
rect 3250 2683 3257 2686
rect 3298 2713 3309 2716
rect 3250 2663 3253 2683
rect 3250 2593 3253 2616
rect 3266 2603 3269 2626
rect 3298 2613 3301 2713
rect 3318 2706 3321 2753
rect 3314 2703 3321 2706
rect 3314 2656 3317 2703
rect 3310 2653 3317 2656
rect 3310 2596 3313 2653
rect 3338 2616 3341 2853
rect 3346 2683 3349 2826
rect 3354 2813 3357 2836
rect 3354 2723 3357 2806
rect 3362 2783 3365 2936
rect 3370 2766 3373 3036
rect 3378 3026 3381 3043
rect 3378 3023 3385 3026
rect 3382 2846 3385 3023
rect 3406 2996 3409 3053
rect 3418 3013 3421 3126
rect 3426 2996 3429 3363
rect 3434 3343 3437 3516
rect 3442 3513 3449 3516
rect 3434 3223 3437 3336
rect 3446 3246 3449 3513
rect 3458 3323 3461 3526
rect 3482 3503 3485 3536
rect 3494 3496 3497 3553
rect 3506 3533 3509 3586
rect 3522 3553 3525 3823
rect 3538 3803 3541 3993
rect 3554 3896 3557 3986
rect 3562 3923 3565 4016
rect 3570 4003 3573 4026
rect 3578 3983 3581 4043
rect 3586 4013 3589 4336
rect 3594 4253 3597 4343
rect 3610 4336 3613 4356
rect 3602 4333 3613 4336
rect 3618 4333 3621 4393
rect 3634 4333 3637 4476
rect 3666 4466 3669 4486
rect 3666 4463 3673 4466
rect 3670 4376 3673 4463
rect 3690 4436 3693 4526
rect 3698 4466 3701 4526
rect 3706 4523 3717 4526
rect 3698 4463 3709 4466
rect 3690 4433 3697 4436
rect 3666 4373 3673 4376
rect 3602 4316 3605 4333
rect 3626 4323 3645 4326
rect 3602 4313 3613 4316
rect 3610 4236 3613 4313
rect 3602 4233 3613 4236
rect 3594 4203 3597 4226
rect 3602 4193 3605 4233
rect 3610 4183 3613 4216
rect 3626 4213 3629 4226
rect 3618 4193 3621 4206
rect 3634 4203 3637 4216
rect 3642 4213 3645 4226
rect 3586 3993 3589 4006
rect 3594 3986 3597 4116
rect 3618 4113 3621 4136
rect 3642 4123 3645 4146
rect 3650 4133 3653 4206
rect 3666 4166 3669 4373
rect 3682 4333 3685 4416
rect 3694 4326 3697 4433
rect 3662 4163 3669 4166
rect 3690 4323 3697 4326
rect 3690 4166 3693 4323
rect 3706 4283 3709 4463
rect 3722 4346 3725 4606
rect 3770 4603 3773 4616
rect 3730 4513 3733 4526
rect 3754 4523 3765 4526
rect 3770 4513 3773 4536
rect 3778 4533 3781 4566
rect 3794 4533 3797 4606
rect 3786 4456 3789 4526
rect 3802 4523 3805 4556
rect 3818 4553 3821 4616
rect 3858 4593 3861 4606
rect 3882 4576 3885 4616
rect 3866 4573 3885 4576
rect 3786 4453 3793 4456
rect 3770 4393 3773 4416
rect 3790 4376 3793 4453
rect 3790 4373 3797 4376
rect 3718 4343 3725 4346
rect 3718 4266 3721 4343
rect 3730 4333 3741 4336
rect 3746 4333 3749 4356
rect 3718 4263 3725 4266
rect 3722 4233 3725 4263
rect 3730 4243 3733 4326
rect 3722 4193 3725 4216
rect 3690 4163 3701 4166
rect 3662 4056 3665 4163
rect 3698 4086 3701 4163
rect 3738 4123 3741 4156
rect 3746 4086 3749 4126
rect 3650 4053 3665 4056
rect 3690 4083 3701 4086
rect 3738 4083 3749 4086
rect 3586 3983 3597 3986
rect 3570 3933 3573 3956
rect 3586 3923 3589 3983
rect 3602 3953 3605 4016
rect 3618 3996 3621 4016
rect 3618 3993 3629 3996
rect 3610 3963 3613 3986
rect 3554 3893 3565 3896
rect 3562 3836 3565 3893
rect 3554 3833 3565 3836
rect 3554 3816 3557 3833
rect 3586 3816 3589 3906
rect 3610 3903 3613 3926
rect 3626 3896 3629 3993
rect 3650 3976 3653 4053
rect 3690 4036 3693 4083
rect 3690 4033 3697 4036
rect 3682 4013 3685 4026
rect 3694 3986 3697 4033
rect 3722 4003 3725 4046
rect 3738 4013 3741 4083
rect 3770 4066 3773 4246
rect 3762 4063 3773 4066
rect 3694 3983 3701 3986
rect 3650 3973 3661 3976
rect 3618 3893 3629 3896
rect 3550 3813 3557 3816
rect 3538 3706 3541 3786
rect 3550 3746 3553 3813
rect 3550 3743 3557 3746
rect 3554 3723 3557 3743
rect 3562 3733 3565 3816
rect 3586 3813 3597 3816
rect 3570 3733 3573 3796
rect 3538 3703 3549 3706
rect 3546 3586 3549 3703
rect 3538 3583 3549 3586
rect 3538 3536 3541 3583
rect 3530 3533 3541 3536
rect 3546 3533 3549 3546
rect 3562 3533 3565 3566
rect 3506 3506 3509 3526
rect 3506 3503 3517 3506
rect 3494 3493 3501 3496
rect 3474 3333 3477 3406
rect 3482 3333 3485 3426
rect 3490 3373 3493 3416
rect 3482 3266 3485 3326
rect 3490 3323 3493 3366
rect 3498 3323 3501 3493
rect 3514 3436 3517 3503
rect 3506 3433 3517 3436
rect 3506 3413 3509 3433
rect 3530 3416 3533 3533
rect 3538 3506 3541 3526
rect 3570 3523 3573 3726
rect 3578 3716 3581 3806
rect 3594 3766 3597 3813
rect 3586 3763 3597 3766
rect 3618 3776 3621 3893
rect 3618 3773 3637 3776
rect 3586 3733 3589 3763
rect 3594 3723 3597 3746
rect 3610 3716 3613 3726
rect 3578 3713 3585 3716
rect 3582 3646 3585 3713
rect 3578 3643 3585 3646
rect 3594 3713 3613 3716
rect 3578 3586 3581 3643
rect 3586 3603 3589 3626
rect 3578 3583 3585 3586
rect 3582 3526 3585 3583
rect 3594 3553 3597 3713
rect 3602 3583 3605 3606
rect 3618 3603 3621 3773
rect 3642 3766 3645 3846
rect 3634 3763 3645 3766
rect 3634 3636 3637 3763
rect 3650 3746 3653 3926
rect 3658 3843 3661 3973
rect 3698 3966 3701 3983
rect 3762 3976 3765 4063
rect 3786 4016 3789 4326
rect 3794 4263 3797 4373
rect 3802 4333 3805 4396
rect 3810 4323 3813 4336
rect 3818 4333 3821 4536
rect 3866 4533 3869 4573
rect 3858 4513 3861 4526
rect 3874 4503 3877 4526
rect 3882 4483 3885 4536
rect 3898 4533 3901 4546
rect 3954 4536 3957 4616
rect 3970 4573 3973 4606
rect 4018 4576 4021 4616
rect 4018 4573 4029 4576
rect 3890 4523 3901 4526
rect 3834 4333 3837 4416
rect 3890 4413 3893 4523
rect 3906 4453 3909 4526
rect 3842 4326 3845 4376
rect 3834 4323 3845 4326
rect 3810 4203 3813 4226
rect 3834 4216 3837 4323
rect 3818 4203 3821 4216
rect 3826 4213 3837 4216
rect 3842 4133 3845 4236
rect 3850 4193 3853 4206
rect 3858 4186 3861 4356
rect 3882 4286 3885 4316
rect 3890 4303 3893 4366
rect 3898 4333 3901 4406
rect 3866 4213 3869 4226
rect 3874 4203 3877 4286
rect 3882 4283 3893 4286
rect 3882 4213 3885 4276
rect 3890 4236 3893 4283
rect 3898 4263 3901 4326
rect 3906 4313 3909 4416
rect 3922 4373 3925 4526
rect 3930 4513 3933 4526
rect 3946 4513 3949 4536
rect 3954 4533 3973 4536
rect 3930 4403 3933 4426
rect 3938 4403 3941 4416
rect 4002 4413 4005 4426
rect 3946 4343 3949 4406
rect 3994 4393 3997 4406
rect 3914 4236 3917 4326
rect 3946 4283 3949 4326
rect 3978 4266 3981 4286
rect 3970 4263 3981 4266
rect 3890 4233 3909 4236
rect 3914 4233 3925 4236
rect 3890 4213 3893 4226
rect 3858 4183 3865 4186
rect 3802 4103 3805 4126
rect 3850 4123 3853 4176
rect 3862 4126 3865 4183
rect 3890 4173 3893 4206
rect 3890 4133 3893 4146
rect 3858 4123 3865 4126
rect 3858 4106 3861 4123
rect 3850 4103 3861 4106
rect 3850 4026 3853 4103
rect 3874 4036 3877 4126
rect 3898 4123 3901 4196
rect 3906 4186 3909 4233
rect 3922 4203 3925 4233
rect 3930 4193 3933 4216
rect 3970 4186 3973 4263
rect 3994 4243 3997 4376
rect 4010 4283 4013 4536
rect 4026 4533 4029 4573
rect 4042 4533 4045 4626
rect 4050 4526 4053 4576
rect 4058 4533 4061 4616
rect 4018 4513 4021 4526
rect 4018 4243 4021 4406
rect 4034 4403 4037 4526
rect 4042 4513 4045 4526
rect 4050 4523 4061 4526
rect 4058 4363 4061 4523
rect 4074 4513 4077 4606
rect 4122 4603 4125 4616
rect 4082 4423 4085 4526
rect 4138 4516 4141 4536
rect 4130 4513 4141 4516
rect 4130 4466 4133 4513
rect 4130 4463 4141 4466
rect 4082 4393 4085 4416
rect 4138 4413 4141 4463
rect 4146 4393 4149 4556
rect 4162 4533 4165 4606
rect 4154 4506 4157 4526
rect 4170 4523 4173 4616
rect 4154 4503 4161 4506
rect 4158 4446 4161 4503
rect 4154 4443 4161 4446
rect 4026 4333 4029 4356
rect 4026 4273 4029 4326
rect 3986 4193 3989 4206
rect 3906 4183 3917 4186
rect 3970 4183 3981 4186
rect 3914 4116 3917 4183
rect 3930 4133 3933 4156
rect 3906 4113 3917 4116
rect 3906 4046 3909 4113
rect 3946 4076 3949 4176
rect 3978 4153 3981 4183
rect 4002 4173 4005 4206
rect 3970 4123 3973 4146
rect 4026 4123 4029 4196
rect 4050 4193 4053 4216
rect 4074 4173 4077 4296
rect 4082 4273 4085 4366
rect 4082 4143 4085 4216
rect 4090 4213 4093 4246
rect 4090 4173 4093 4206
rect 4090 4093 4093 4136
rect 3946 4073 3965 4076
rect 3906 4043 3917 4046
rect 3870 4033 3877 4036
rect 3850 4023 3861 4026
rect 3778 4013 3789 4016
rect 3762 3973 3773 3976
rect 3698 3963 3705 3966
rect 3666 3836 3669 3926
rect 3690 3923 3693 3956
rect 3702 3916 3705 3963
rect 3746 3923 3749 3936
rect 3770 3933 3773 3973
rect 3778 3956 3781 4013
rect 3786 3973 3789 4006
rect 3778 3953 3789 3956
rect 3794 3953 3797 4006
rect 3802 3996 3805 4016
rect 3802 3993 3813 3996
rect 3698 3913 3705 3916
rect 3698 3846 3701 3913
rect 3698 3843 3709 3846
rect 3658 3833 3669 3836
rect 3658 3803 3661 3833
rect 3674 3763 3677 3806
rect 3706 3796 3709 3843
rect 3698 3793 3709 3796
rect 3722 3793 3725 3816
rect 3698 3746 3701 3793
rect 3650 3743 3661 3746
rect 3658 3666 3661 3743
rect 3630 3633 3637 3636
rect 3650 3663 3661 3666
rect 3690 3743 3701 3746
rect 3630 3566 3633 3633
rect 3650 3576 3653 3663
rect 3674 3613 3677 3626
rect 3690 3586 3693 3743
rect 3714 3616 3717 3736
rect 3722 3733 3725 3746
rect 3754 3743 3757 3816
rect 3714 3613 3733 3616
rect 3690 3583 3701 3586
rect 3650 3573 3677 3576
rect 3630 3563 3637 3566
rect 3578 3523 3585 3526
rect 3578 3506 3581 3523
rect 3538 3503 3549 3506
rect 3546 3446 3549 3503
rect 3538 3443 3549 3446
rect 3570 3503 3581 3506
rect 3538 3423 3541 3443
rect 3514 3403 3517 3416
rect 3530 3413 3541 3416
rect 3522 3323 3525 3336
rect 3538 3333 3541 3413
rect 3570 3396 3573 3503
rect 3594 3403 3597 3526
rect 3626 3523 3629 3546
rect 3570 3393 3577 3396
rect 3478 3263 3485 3266
rect 3442 3243 3449 3246
rect 3442 3196 3445 3243
rect 3466 3233 3469 3246
rect 3450 3213 3453 3226
rect 3478 3206 3481 3263
rect 3490 3233 3493 3256
rect 3498 3223 3501 3236
rect 3506 3216 3509 3316
rect 3574 3296 3577 3393
rect 3586 3323 3589 3346
rect 3618 3336 3621 3436
rect 3610 3333 3621 3336
rect 3574 3293 3581 3296
rect 3578 3276 3581 3293
rect 3538 3223 3541 3246
rect 3562 3223 3565 3236
rect 3490 3213 3509 3216
rect 3570 3213 3573 3276
rect 3578 3273 3589 3276
rect 3586 3206 3589 3273
rect 3610 3246 3613 3333
rect 3610 3243 3621 3246
rect 3602 3223 3613 3226
rect 3478 3203 3485 3206
rect 3442 3193 3461 3196
rect 3458 3046 3461 3193
rect 3482 3136 3485 3203
rect 3578 3203 3589 3206
rect 3610 3203 3613 3216
rect 3578 3166 3581 3203
rect 3618 3186 3621 3243
rect 3626 3213 3629 3326
rect 3610 3183 3621 3186
rect 3578 3163 3589 3166
rect 3446 3043 3461 3046
rect 3474 3133 3485 3136
rect 3474 3046 3477 3133
rect 3474 3043 3485 3046
rect 3402 2993 3409 2996
rect 3418 2993 3429 2996
rect 3402 2896 3405 2993
rect 3366 2763 3373 2766
rect 3378 2843 3385 2846
rect 3394 2893 3405 2896
rect 3418 2896 3421 2993
rect 3434 2976 3437 3026
rect 3430 2973 3437 2976
rect 3430 2916 3433 2973
rect 3446 2966 3449 3043
rect 3474 3013 3477 3026
rect 3482 3016 3485 3043
rect 3490 3023 3493 3126
rect 3506 3033 3509 3136
rect 3482 3013 3493 3016
rect 3442 2963 3449 2966
rect 3442 2926 3445 2963
rect 3442 2923 3449 2926
rect 3430 2913 3437 2916
rect 3418 2893 3429 2896
rect 3366 2676 3369 2763
rect 3366 2673 3373 2676
rect 3370 2656 3373 2673
rect 3378 2663 3381 2843
rect 3394 2836 3397 2893
rect 3418 2856 3421 2876
rect 3414 2853 3421 2856
rect 3394 2833 3405 2836
rect 3386 2703 3389 2826
rect 3402 2736 3405 2833
rect 3414 2776 3417 2853
rect 3414 2773 3421 2776
rect 3418 2753 3421 2773
rect 3394 2733 3405 2736
rect 3394 2713 3397 2733
rect 3370 2653 3381 2656
rect 3334 2613 3341 2616
rect 3210 2503 3229 2506
rect 3178 2413 3189 2416
rect 3154 2323 3165 2326
rect 3178 2323 3181 2413
rect 3210 2396 3213 2503
rect 3234 2416 3237 2536
rect 3242 2533 3253 2536
rect 3282 2533 3285 2596
rect 3310 2593 3317 2596
rect 3242 2493 3245 2526
rect 3250 2503 3253 2533
rect 3266 2523 3293 2526
rect 3274 2486 3277 2506
rect 3266 2483 3277 2486
rect 3266 2416 3269 2483
rect 3234 2413 3253 2416
rect 3266 2413 3273 2416
rect 3234 2403 3237 2413
rect 3210 2393 3237 2396
rect 3242 2393 3245 2406
rect 3250 2396 3253 2413
rect 3250 2393 3261 2396
rect 3226 2333 3229 2346
rect 3194 2313 3197 2326
rect 3186 2206 3189 2256
rect 3218 2213 3221 2226
rect 3226 2213 3229 2316
rect 3234 2296 3237 2393
rect 3250 2333 3253 2393
rect 3270 2356 3273 2413
rect 3270 2353 3277 2356
rect 3234 2293 3245 2296
rect 3242 2236 3245 2293
rect 3234 2233 3245 2236
rect 3186 2203 3205 2206
rect 3130 2123 3133 2136
rect 3138 2133 3141 2146
rect 3146 2106 3149 2126
rect 3154 2123 3157 2136
rect 3202 2133 3205 2203
rect 3226 2123 3229 2146
rect 3234 2116 3237 2233
rect 3242 2213 3253 2216
rect 3242 2203 3245 2213
rect 3266 2203 3269 2226
rect 3242 2176 3245 2196
rect 3274 2186 3277 2353
rect 3282 2343 3285 2523
rect 3314 2476 3317 2593
rect 3334 2556 3337 2613
rect 3330 2553 3337 2556
rect 3330 2496 3333 2553
rect 3330 2493 3337 2496
rect 3314 2473 3325 2476
rect 3306 2433 3317 2436
rect 3290 2256 3293 2426
rect 3298 2323 3301 2346
rect 3290 2253 3301 2256
rect 3270 2183 3277 2186
rect 3242 2173 3249 2176
rect 3138 2103 3149 2106
rect 3226 2113 3237 2116
rect 3122 1973 3125 2016
rect 3138 2013 3141 2103
rect 3226 2096 3229 2113
rect 3246 2106 3249 2173
rect 3218 2093 3229 2096
rect 3242 2103 3249 2106
rect 3130 1966 3133 2006
rect 3154 2003 3157 2026
rect 3122 1963 3133 1966
rect 3122 1923 3125 1963
rect 3138 1956 3141 1976
rect 3138 1953 3145 1956
rect 3142 1886 3145 1953
rect 3186 1933 3189 2006
rect 3202 1963 3205 2036
rect 3218 2023 3221 2093
rect 3242 2046 3245 2103
rect 3234 2043 3245 2046
rect 3234 1946 3237 2043
rect 3234 1943 3245 1946
rect 3090 1746 3093 1776
rect 3074 1743 3093 1746
rect 3074 1733 3077 1743
rect 3106 1736 3109 1886
rect 3138 1883 3145 1886
rect 3090 1733 3109 1736
rect 3114 1733 3117 1796
rect 3122 1793 3125 1806
rect 3042 1713 3045 1726
rect 3090 1646 3093 1733
rect 3074 1643 3093 1646
rect 3018 1543 3021 1556
rect 3002 1533 3029 1536
rect 3034 1533 3037 1626
rect 3042 1603 3045 1616
rect 2994 1436 2997 1526
rect 3018 1506 3021 1526
rect 3010 1503 3021 1506
rect 3026 1506 3029 1533
rect 3026 1503 3037 1506
rect 3010 1456 3013 1503
rect 3010 1453 3021 1456
rect 2994 1433 3005 1436
rect 2898 1413 2901 1426
rect 3002 1416 3005 1433
rect 2850 1323 2853 1356
rect 2866 1353 2885 1356
rect 2866 1336 2869 1353
rect 2862 1333 2869 1336
rect 2906 1333 2909 1416
rect 2994 1413 3005 1416
rect 2994 1393 2997 1413
rect 3010 1403 3013 1416
rect 3018 1413 3021 1453
rect 3034 1406 3037 1503
rect 3026 1403 3037 1406
rect 3050 1403 3053 1566
rect 3074 1556 3077 1643
rect 3098 1613 3101 1636
rect 3106 1606 3109 1656
rect 3130 1633 3133 1816
rect 3138 1813 3141 1883
rect 3154 1803 3157 1926
rect 3162 1833 3165 1916
rect 3226 1913 3229 1926
rect 3218 1873 3221 1906
rect 3242 1843 3245 1943
rect 3250 1913 3253 2036
rect 3258 2033 3261 2066
rect 3270 2046 3273 2183
rect 3270 2043 3277 2046
rect 3266 2013 3269 2026
rect 3274 1996 3277 2043
rect 3266 1993 3277 1996
rect 3266 1926 3269 1993
rect 3282 1933 3285 2246
rect 3298 2156 3301 2253
rect 3322 2243 3325 2473
rect 3334 2426 3337 2493
rect 3346 2433 3349 2606
rect 3370 2603 3373 2626
rect 3378 2533 3381 2653
rect 3394 2613 3397 2686
rect 3410 2673 3413 2706
rect 3426 2676 3429 2893
rect 3434 2813 3437 2913
rect 3446 2856 3449 2923
rect 3442 2853 3449 2856
rect 3434 2683 3437 2736
rect 3442 2706 3445 2853
rect 3450 2823 3453 2836
rect 3458 2713 3461 3006
rect 3466 3003 3477 3006
rect 3466 2816 3469 2836
rect 3474 2823 3477 2876
rect 3482 2833 3485 3013
rect 3490 2993 3493 3006
rect 3498 2933 3501 3006
rect 3506 2916 3509 3016
rect 3514 3003 3517 3086
rect 3522 3013 3541 3016
rect 3522 3003 3525 3013
rect 3530 2946 3533 3006
rect 3522 2943 3533 2946
rect 3498 2913 3509 2916
rect 3498 2836 3501 2913
rect 3498 2833 3509 2836
rect 3466 2813 3477 2816
rect 3474 2726 3477 2813
rect 3482 2803 3485 2826
rect 3490 2733 3493 2816
rect 3498 2743 3501 2806
rect 3506 2783 3509 2833
rect 3474 2723 3485 2726
rect 3442 2703 3453 2706
rect 3426 2673 3433 2676
rect 3410 2583 3413 2636
rect 3418 2613 3421 2626
rect 3354 2523 3381 2526
rect 3334 2423 3341 2426
rect 3362 2423 3365 2506
rect 3338 2226 3341 2423
rect 3370 2413 3373 2426
rect 3314 2203 3317 2226
rect 3322 2223 3341 2226
rect 3322 2196 3325 2223
rect 3322 2193 3333 2196
rect 3294 2153 3301 2156
rect 3294 1956 3297 2153
rect 3330 2136 3333 2193
rect 3306 2123 3309 2136
rect 3330 2133 3341 2136
rect 3306 2013 3309 2026
rect 3290 1953 3297 1956
rect 3266 1923 3277 1926
rect 3274 1883 3277 1923
rect 3154 1773 3157 1796
rect 3154 1723 3157 1736
rect 3138 1653 3141 1716
rect 3170 1703 3173 1806
rect 3178 1743 3181 1806
rect 3186 1753 3189 1816
rect 3234 1793 3237 1836
rect 3226 1746 3229 1766
rect 3222 1743 3229 1746
rect 3178 1713 3181 1726
rect 3186 1703 3189 1716
rect 3098 1603 3109 1606
rect 3074 1553 3093 1556
rect 3082 1523 3085 1536
rect 3090 1506 3093 1553
rect 3098 1536 3101 1603
rect 3106 1543 3109 1556
rect 3098 1533 3109 1536
rect 3114 1533 3117 1596
rect 3202 1563 3205 1616
rect 3146 1533 3149 1556
rect 3082 1503 3093 1506
rect 3082 1456 3085 1503
rect 3082 1453 3093 1456
rect 3090 1433 3093 1453
rect 3026 1356 3029 1403
rect 3018 1353 3029 1356
rect 2962 1343 2981 1346
rect 2962 1333 2973 1336
rect 2978 1333 2981 1343
rect 2862 1276 2865 1333
rect 2874 1296 2877 1326
rect 3018 1313 3021 1353
rect 3026 1296 3029 1346
rect 3058 1343 3061 1406
rect 3082 1386 3085 1416
rect 3074 1383 3085 1386
rect 3090 1383 3093 1396
rect 3034 1323 3061 1326
rect 2874 1293 2881 1296
rect 2862 1273 2869 1276
rect 2866 1253 2869 1273
rect 2878 1216 2881 1293
rect 3018 1293 3029 1296
rect 2714 1153 2741 1156
rect 2666 1083 2677 1086
rect 2650 913 2653 926
rect 2658 903 2661 926
rect 2618 883 2625 886
rect 2602 713 2605 726
rect 2618 706 2621 883
rect 2594 603 2597 706
rect 2602 703 2621 706
rect 2554 533 2557 546
rect 2602 523 2605 703
rect 2610 573 2613 676
rect 2634 613 2637 626
rect 2642 603 2645 716
rect 2666 703 2669 1083
rect 2674 1013 2677 1026
rect 2682 1013 2685 1036
rect 2690 1013 2693 1026
rect 2674 1003 2693 1006
rect 2714 963 2717 1153
rect 2730 1133 2733 1146
rect 2778 1143 2781 1216
rect 2866 1206 2869 1216
rect 2878 1213 2885 1216
rect 2866 1203 2877 1206
rect 2882 1203 2885 1213
rect 2890 1196 2893 1236
rect 2866 1193 2893 1196
rect 2850 1143 2853 1156
rect 2858 1133 2861 1146
rect 2730 1113 2733 1126
rect 2762 1063 2765 1126
rect 2770 1013 2773 1036
rect 2866 1033 2869 1136
rect 2890 1133 2893 1146
rect 2874 1113 2877 1126
rect 2898 1103 2901 1256
rect 2906 1183 2909 1196
rect 2994 1166 2997 1216
rect 3002 1213 3005 1246
rect 3018 1236 3021 1293
rect 3018 1233 3029 1236
rect 3026 1216 3029 1233
rect 3034 1223 3037 1316
rect 3026 1213 3033 1216
rect 3002 1203 3013 1206
rect 3018 1183 3021 1206
rect 2994 1163 3005 1166
rect 2906 1036 2909 1126
rect 2994 1123 2997 1146
rect 3002 1133 3005 1163
rect 3010 1133 3013 1156
rect 3030 1136 3033 1213
rect 3030 1133 3037 1136
rect 3010 1086 3013 1106
rect 3002 1083 3013 1086
rect 2906 1033 2917 1036
rect 2714 923 2717 956
rect 2674 813 2677 826
rect 2698 773 2701 806
rect 2714 783 2717 806
rect 2730 723 2733 836
rect 2738 773 2741 966
rect 2794 963 2797 1006
rect 2810 983 2813 1006
rect 2754 913 2757 926
rect 2818 913 2821 1016
rect 2842 963 2845 1016
rect 2826 923 2829 936
rect 2850 933 2853 976
rect 2746 763 2749 816
rect 2850 813 2853 836
rect 2866 803 2869 966
rect 2874 933 2877 1016
rect 2938 1003 2941 1066
rect 2946 996 2949 1006
rect 2930 993 2949 996
rect 3002 976 3005 1083
rect 3018 1016 3021 1126
rect 3018 1013 3029 1016
rect 3026 1003 3029 1013
rect 3034 996 3037 1133
rect 3042 1053 3045 1316
rect 3066 1303 3069 1316
rect 3074 1303 3077 1383
rect 3082 1333 3085 1346
rect 3098 1343 3101 1416
rect 3106 1403 3109 1533
rect 3114 1513 3117 1526
rect 3122 1506 3125 1526
rect 3186 1516 3189 1536
rect 3122 1503 3133 1506
rect 3130 1436 3133 1503
rect 3114 1403 3117 1436
rect 3122 1433 3133 1436
rect 3122 1413 3125 1433
rect 3130 1403 3133 1416
rect 3154 1396 3157 1516
rect 3178 1513 3189 1516
rect 3178 1416 3181 1513
rect 3194 1423 3197 1536
rect 3202 1513 3205 1536
rect 3210 1533 3213 1716
rect 3222 1646 3225 1743
rect 3222 1643 3229 1646
rect 3226 1626 3229 1643
rect 3234 1633 3237 1726
rect 3242 1713 3245 1816
rect 3250 1713 3253 1876
rect 3290 1873 3293 1953
rect 3314 1936 3317 2026
rect 3322 2003 3325 2036
rect 3330 2006 3333 2116
rect 3338 2023 3341 2133
rect 3346 2023 3349 2216
rect 3354 2203 3357 2326
rect 3362 2323 3365 2336
rect 3378 2293 3381 2436
rect 3394 2423 3397 2536
rect 3418 2533 3421 2606
rect 3430 2586 3433 2673
rect 3442 2593 3445 2646
rect 3430 2583 3437 2586
rect 3402 2523 3429 2526
rect 3434 2516 3437 2583
rect 3426 2513 3437 2516
rect 3426 2446 3429 2513
rect 3450 2503 3453 2703
rect 3458 2613 3461 2626
rect 3458 2533 3461 2576
rect 3458 2513 3461 2526
rect 3466 2496 3469 2716
rect 3418 2443 3429 2446
rect 3462 2493 3469 2496
rect 3354 2053 3357 2136
rect 3362 2113 3365 2236
rect 3370 2133 3373 2206
rect 3378 2193 3381 2276
rect 3378 2123 3381 2166
rect 3386 2116 3389 2156
rect 3378 2113 3389 2116
rect 3330 2003 3341 2006
rect 3338 1946 3341 2003
rect 3330 1943 3341 1946
rect 3282 1833 3301 1836
rect 3282 1823 3293 1826
rect 3298 1816 3301 1826
rect 3258 1813 3301 1816
rect 3306 1796 3309 1936
rect 3314 1933 3325 1936
rect 3298 1793 3309 1796
rect 3258 1656 3261 1746
rect 3298 1706 3301 1793
rect 3314 1743 3317 1926
rect 3322 1846 3325 1933
rect 3330 1923 3333 1943
rect 3330 1913 3341 1916
rect 3322 1843 3333 1846
rect 3322 1713 3325 1836
rect 3298 1703 3309 1706
rect 3250 1653 3261 1656
rect 3226 1623 3237 1626
rect 3234 1596 3237 1623
rect 3242 1603 3245 1636
rect 3250 1623 3253 1653
rect 3306 1643 3309 1703
rect 3330 1656 3333 1843
rect 3338 1813 3341 1826
rect 3322 1653 3333 1656
rect 3258 1613 3261 1626
rect 3274 1623 3293 1626
rect 3234 1593 3245 1596
rect 3210 1506 3213 1526
rect 3242 1523 3245 1593
rect 3266 1513 3269 1606
rect 3210 1503 3221 1506
rect 3218 1436 3221 1503
rect 3210 1433 3221 1436
rect 3178 1413 3189 1416
rect 3154 1393 3165 1396
rect 3042 1013 3045 1036
rect 3026 976 3029 996
rect 3034 993 3041 996
rect 3050 993 3053 1226
rect 3058 1116 3061 1246
rect 3082 1233 3085 1326
rect 3074 1213 3077 1226
rect 3066 1133 3069 1146
rect 3058 1113 3065 1116
rect 3062 1046 3065 1113
rect 3082 1103 3085 1126
rect 3058 1043 3065 1046
rect 3002 973 3013 976
rect 2882 943 2885 956
rect 2978 933 2989 936
rect 2994 933 2997 956
rect 2970 836 2973 926
rect 2978 913 2981 926
rect 3010 916 3013 973
rect 3002 913 3013 916
rect 3022 973 3029 976
rect 3002 856 3005 913
rect 3002 853 3013 856
rect 2970 833 2989 836
rect 2834 783 2837 796
rect 2754 706 2757 776
rect 2874 773 2877 826
rect 2770 723 2773 766
rect 2810 733 2813 746
rect 2818 726 2821 736
rect 2802 723 2821 726
rect 2754 703 2765 706
rect 2762 626 2765 703
rect 2802 673 2805 723
rect 2850 713 2853 726
rect 2762 623 2773 626
rect 2522 493 2533 496
rect 2530 436 2533 493
rect 2522 433 2533 436
rect 2522 413 2525 433
rect 2554 413 2557 426
rect 2562 413 2565 426
rect 2578 413 2581 426
rect 2602 413 2605 426
rect 2522 393 2525 406
rect 2546 366 2549 406
rect 2530 363 2549 366
rect 2530 323 2533 363
rect 2554 333 2557 346
rect 2570 303 2573 336
rect 2586 323 2589 406
rect 2618 393 2621 416
rect 2362 13 2373 16
rect 2466 13 2469 196
rect 2490 193 2493 206
rect 2362 0 2365 13
rect 2490 0 2493 126
rect 2514 123 2517 226
rect 2578 213 2581 286
rect 2578 123 2581 206
rect 2586 153 2589 216
rect 2618 213 2621 316
rect 2626 296 2629 436
rect 2634 423 2637 526
rect 2650 523 2653 616
rect 2754 583 2757 616
rect 2770 576 2773 623
rect 2818 593 2821 616
rect 2874 613 2877 746
rect 2890 723 2893 816
rect 2986 803 2989 833
rect 2922 733 2925 746
rect 2914 676 2917 726
rect 2914 673 2925 676
rect 2762 573 2773 576
rect 2658 366 2661 546
rect 2706 523 2709 536
rect 2730 533 2733 546
rect 2762 543 2765 573
rect 2842 543 2845 606
rect 2858 593 2861 606
rect 2898 543 2901 556
rect 2706 413 2709 426
rect 2650 363 2661 366
rect 2650 333 2653 363
rect 2626 293 2637 296
rect 2634 236 2637 293
rect 2626 233 2637 236
rect 2602 196 2605 206
rect 2626 203 2629 233
rect 2602 193 2621 196
rect 2586 133 2589 146
rect 2514 0 2517 116
rect 2602 113 2605 126
rect 2610 123 2613 146
rect 2618 116 2621 156
rect 2634 143 2637 206
rect 2650 203 2653 216
rect 2674 213 2677 326
rect 2682 213 2685 226
rect 2698 223 2701 236
rect 2714 213 2717 236
rect 2722 213 2725 226
rect 2746 213 2749 416
rect 2786 413 2789 426
rect 2762 393 2765 406
rect 2770 283 2773 346
rect 2794 323 2797 336
rect 2802 313 2805 406
rect 2842 403 2845 416
rect 2906 413 2909 536
rect 2922 533 2925 673
rect 2930 423 2933 526
rect 2946 423 2949 536
rect 2954 513 2957 796
rect 2978 736 2981 796
rect 2994 783 2997 806
rect 3010 793 3013 853
rect 3022 746 3025 973
rect 3038 926 3041 993
rect 3058 966 3061 1043
rect 3050 963 3061 966
rect 3038 923 3045 926
rect 3042 906 3045 923
rect 3034 903 3045 906
rect 3022 743 3029 746
rect 2970 733 2981 736
rect 2986 623 2989 726
rect 2994 713 2997 736
rect 3018 713 3021 726
rect 2994 613 2997 626
rect 2970 533 2973 556
rect 2866 393 2869 406
rect 2818 313 2821 346
rect 2706 203 2725 206
rect 2722 183 2725 203
rect 2762 193 2765 206
rect 2770 203 2773 216
rect 2778 203 2781 226
rect 2794 203 2797 216
rect 2802 193 2805 216
rect 2818 183 2821 216
rect 2834 203 2837 216
rect 2842 193 2845 206
rect 2698 133 2701 146
rect 2722 133 2725 176
rect 2610 113 2621 116
rect 2650 113 2653 126
rect 2770 123 2773 146
rect 2826 133 2829 146
rect 2834 123 2837 146
rect 2850 133 2853 206
rect 2858 203 2861 326
rect 2858 123 2861 186
rect 2866 123 2869 236
rect 2874 223 2893 226
rect 2874 203 2877 223
rect 2882 193 2885 216
rect 2890 213 2893 223
rect 2898 153 2901 326
rect 2914 306 2917 326
rect 2914 303 2925 306
rect 2922 246 2925 303
rect 2914 243 2925 246
rect 2914 203 2917 243
rect 2922 193 2925 206
rect 2882 123 2885 136
rect 2866 113 2877 116
rect 2890 103 2893 136
rect 2898 133 2901 146
rect 2906 123 2909 186
rect 2914 133 2925 136
rect 2930 133 2933 216
rect 2938 213 2941 226
rect 2946 193 2949 416
rect 2970 413 2973 526
rect 2994 436 2997 516
rect 3010 513 3013 616
rect 3026 593 3029 743
rect 3034 713 3037 903
rect 3050 826 3053 963
rect 3046 823 3053 826
rect 3046 756 3049 823
rect 3058 763 3061 816
rect 3066 783 3069 806
rect 3046 753 3053 756
rect 3042 703 3045 736
rect 3050 723 3053 753
rect 3066 733 3069 746
rect 3066 703 3069 726
rect 3074 693 3077 1056
rect 3082 1023 3085 1046
rect 3082 903 3085 916
rect 3082 813 3085 826
rect 3090 813 3093 1266
rect 3106 1233 3109 1326
rect 3114 1256 3117 1346
rect 3122 1263 3125 1326
rect 3138 1323 3141 1336
rect 3146 1333 3149 1386
rect 3162 1336 3165 1393
rect 3154 1333 3165 1336
rect 3114 1253 3125 1256
rect 3098 1213 3101 1226
rect 3114 1223 3117 1246
rect 3122 1203 3125 1253
rect 3154 1223 3157 1333
rect 3186 1293 3189 1413
rect 3210 1346 3213 1433
rect 3250 1423 3269 1426
rect 3202 1343 3213 1346
rect 3202 1326 3205 1343
rect 3198 1323 3205 1326
rect 3186 1203 3189 1236
rect 3198 1226 3201 1323
rect 3210 1313 3213 1336
rect 3218 1333 3221 1356
rect 3198 1223 3205 1226
rect 3194 1193 3197 1206
rect 3106 1133 3109 1156
rect 3146 1143 3149 1156
rect 3202 1146 3205 1223
rect 3210 1203 3213 1296
rect 3234 1253 3237 1416
rect 3242 1396 3245 1416
rect 3266 1413 3269 1423
rect 3274 1396 3277 1596
rect 3242 1393 3253 1396
rect 3250 1286 3253 1393
rect 3242 1283 3253 1286
rect 3266 1393 3277 1396
rect 3226 1213 3229 1226
rect 3234 1183 3237 1216
rect 3242 1213 3245 1283
rect 3202 1143 3213 1146
rect 3106 1123 3125 1126
rect 3098 1103 3101 1116
rect 3098 1033 3101 1096
rect 3130 1093 3133 1126
rect 3138 1113 3141 1136
rect 3178 1123 3181 1136
rect 3186 1106 3189 1136
rect 3178 1103 3189 1106
rect 3194 1103 3197 1126
rect 3178 1036 3181 1103
rect 3210 1096 3213 1143
rect 3202 1093 3213 1096
rect 3106 923 3109 1026
rect 3114 1023 3117 1036
rect 3178 1033 3189 1036
rect 3154 943 3157 1006
rect 3178 933 3181 1016
rect 3186 926 3189 1033
rect 3194 1003 3197 1026
rect 3114 906 3117 926
rect 3098 903 3117 906
rect 3138 893 3141 916
rect 3082 803 3093 806
rect 3098 803 3101 816
rect 3082 793 3085 803
rect 3098 783 3101 796
rect 3034 623 3037 636
rect 3050 633 3069 636
rect 3042 613 3045 626
rect 3018 503 3021 516
rect 2994 433 3005 436
rect 2986 323 2989 406
rect 2994 393 2997 426
rect 3002 393 3005 433
rect 3050 426 3053 616
rect 3066 613 3069 633
rect 3074 573 3077 626
rect 3082 613 3085 716
rect 3082 583 3085 596
rect 3074 533 3077 546
rect 3082 516 3085 556
rect 3078 513 3085 516
rect 3078 446 3081 513
rect 3078 443 3085 446
rect 3042 423 3053 426
rect 3066 423 3069 436
rect 3026 333 3029 396
rect 3042 366 3045 423
rect 3042 363 3053 366
rect 3050 343 3053 363
rect 3058 346 3061 416
rect 3058 343 3069 346
rect 2978 213 2989 216
rect 2914 123 2925 126
rect 2938 123 2941 146
rect 2954 123 2957 156
rect 2970 133 2973 146
rect 2978 133 2981 206
rect 2994 133 2997 206
rect 3002 193 3005 216
rect 3026 203 3029 316
rect 3042 283 3045 336
rect 3058 293 3061 326
rect 3066 323 3069 343
rect 3074 326 3077 426
rect 3082 423 3085 443
rect 3074 323 3085 326
rect 3066 213 3069 246
rect 3090 213 3093 766
rect 3098 603 3101 726
rect 3106 613 3109 816
rect 3114 803 3117 826
rect 3122 813 3133 816
rect 3114 623 3117 706
rect 3122 703 3125 806
rect 3146 796 3149 926
rect 3178 923 3189 926
rect 3154 876 3157 896
rect 3154 873 3165 876
rect 3142 793 3149 796
rect 3130 713 3133 726
rect 3142 646 3145 793
rect 3162 786 3165 873
rect 3178 813 3181 923
rect 3154 783 3165 786
rect 3142 643 3149 646
rect 3138 613 3141 626
rect 3146 606 3149 643
rect 3106 583 3109 606
rect 3130 603 3149 606
rect 3098 423 3101 536
rect 3106 426 3109 576
rect 3130 546 3133 603
rect 3154 586 3157 783
rect 3178 773 3181 806
rect 3162 713 3165 766
rect 3186 753 3189 816
rect 3202 753 3205 1093
rect 3218 933 3221 1006
rect 3234 933 3237 1176
rect 3242 1133 3245 1206
rect 3250 1203 3253 1226
rect 3258 1213 3261 1246
rect 3258 1133 3261 1156
rect 3242 1113 3245 1126
rect 3266 1096 3269 1393
rect 3274 1263 3277 1326
rect 3282 1286 3285 1616
rect 3290 1603 3293 1623
rect 3298 1603 3301 1616
rect 3322 1593 3325 1653
rect 3330 1603 3333 1646
rect 3338 1623 3341 1746
rect 3346 1703 3349 1826
rect 3354 1683 3357 1836
rect 3362 1813 3365 2106
rect 3378 1923 3381 2113
rect 3370 1893 3373 1906
rect 3386 1823 3389 1946
rect 3394 1916 3397 2416
rect 3418 2366 3421 2443
rect 3442 2403 3445 2436
rect 3450 2413 3453 2426
rect 3462 2396 3465 2493
rect 3458 2393 3465 2396
rect 3418 2363 3429 2366
rect 3402 2333 3413 2336
rect 3418 2333 3421 2346
rect 3410 2313 3413 2326
rect 3426 2316 3429 2363
rect 3422 2313 3429 2316
rect 3422 2236 3425 2313
rect 3422 2233 3429 2236
rect 3418 2203 3421 2216
rect 3426 2186 3429 2233
rect 3418 2183 3429 2186
rect 3402 2103 3405 2116
rect 3418 2086 3421 2183
rect 3434 2093 3437 2336
rect 3442 2333 3445 2356
rect 3458 2346 3461 2393
rect 3474 2356 3477 2666
rect 3482 2523 3485 2676
rect 3490 2603 3493 2686
rect 3498 2623 3501 2726
rect 3506 2696 3509 2776
rect 3514 2733 3517 2926
rect 3522 2816 3525 2943
rect 3530 2833 3533 2936
rect 3538 2903 3541 2996
rect 3546 2856 3549 3136
rect 3554 3113 3557 3126
rect 3586 3086 3589 3163
rect 3610 3116 3613 3183
rect 3626 3133 3629 3206
rect 3634 3163 3637 3563
rect 3642 3476 3645 3556
rect 3674 3533 3677 3573
rect 3642 3473 3653 3476
rect 3650 3376 3653 3473
rect 3690 3436 3693 3566
rect 3698 3463 3701 3583
rect 3690 3433 3697 3436
rect 3642 3373 3653 3376
rect 3642 3193 3645 3373
rect 3658 3336 3661 3356
rect 3650 3333 3661 3336
rect 3666 3333 3669 3346
rect 3650 3213 3653 3256
rect 3658 3203 3661 3326
rect 3682 3323 3685 3416
rect 3694 3356 3697 3433
rect 3706 3403 3709 3576
rect 3722 3533 3725 3546
rect 3714 3513 3717 3526
rect 3730 3503 3733 3526
rect 3738 3523 3741 3536
rect 3746 3506 3749 3616
rect 3754 3533 3757 3576
rect 3754 3513 3757 3526
rect 3762 3523 3765 3566
rect 3770 3553 3773 3816
rect 3786 3813 3789 3953
rect 3810 3946 3813 3993
rect 3802 3943 3813 3946
rect 3802 3803 3805 3943
rect 3810 3813 3813 3896
rect 3826 3836 3829 4006
rect 3858 4003 3861 4023
rect 3858 3936 3861 3996
rect 3870 3986 3873 4033
rect 3870 3983 3877 3986
rect 3834 3933 3845 3936
rect 3858 3933 3869 3936
rect 3834 3903 3837 3926
rect 3826 3833 3845 3836
rect 3826 3796 3829 3816
rect 3786 3733 3789 3746
rect 3802 3733 3805 3796
rect 3810 3793 3829 3796
rect 3778 3723 3797 3726
rect 3794 3646 3797 3723
rect 3786 3636 3789 3646
rect 3794 3643 3805 3646
rect 3786 3633 3797 3636
rect 3786 3603 3789 3626
rect 3794 3613 3797 3633
rect 3802 3603 3805 3643
rect 3810 3613 3813 3793
rect 3818 3733 3821 3786
rect 3810 3576 3813 3606
rect 3770 3513 3773 3536
rect 3746 3503 3765 3506
rect 3722 3376 3725 3466
rect 3690 3353 3697 3356
rect 3714 3373 3725 3376
rect 3690 3333 3693 3353
rect 3714 3326 3717 3373
rect 3730 3333 3733 3366
rect 3738 3333 3741 3346
rect 3666 3213 3669 3306
rect 3690 3253 3693 3326
rect 3714 3323 3725 3326
rect 3746 3323 3749 3496
rect 3762 3323 3765 3503
rect 3778 3333 3781 3526
rect 3786 3523 3789 3536
rect 3794 3413 3797 3576
rect 3802 3573 3813 3576
rect 3818 3573 3821 3726
rect 3826 3706 3829 3746
rect 3834 3723 3837 3816
rect 3826 3703 3833 3706
rect 3830 3636 3833 3703
rect 3826 3633 3833 3636
rect 3802 3533 3805 3573
rect 3826 3566 3829 3633
rect 3834 3573 3837 3616
rect 3842 3603 3845 3833
rect 3810 3563 3829 3566
rect 3850 3563 3853 3926
rect 3866 3916 3869 3933
rect 3862 3913 3869 3916
rect 3862 3846 3865 3913
rect 3862 3843 3869 3846
rect 3858 3803 3861 3826
rect 3866 3803 3869 3843
rect 3874 3813 3877 3983
rect 3890 3973 3893 4006
rect 3914 3956 3917 4043
rect 3938 3963 3941 4016
rect 3962 3976 3965 4073
rect 4098 4056 4101 4216
rect 4106 4203 4109 4326
rect 4114 4213 4133 4216
rect 4106 4133 4109 4196
rect 4122 4133 4125 4206
rect 4154 4166 4157 4443
rect 4170 4356 4173 4516
rect 4194 4456 4197 4536
rect 4202 4483 4205 4536
rect 4194 4453 4201 4456
rect 4198 4376 4201 4453
rect 4218 4433 4221 4606
rect 4242 4533 4245 4556
rect 4258 4533 4261 4616
rect 4274 4533 4277 4546
rect 4298 4533 4301 4616
rect 4338 4593 4341 4606
rect 4386 4603 4389 4616
rect 4250 4523 4261 4526
rect 4266 4523 4285 4526
rect 4322 4446 4325 4526
rect 4330 4503 4333 4526
rect 4346 4523 4349 4536
rect 4322 4443 4329 4446
rect 4194 4373 4201 4376
rect 4170 4353 4189 4356
rect 4194 4353 4197 4373
rect 4178 4333 4181 4346
rect 4170 4203 4173 4326
rect 4178 4283 4181 4326
rect 4186 4293 4189 4353
rect 4210 4333 4213 4416
rect 4218 4326 4221 4336
rect 4226 4333 4229 4356
rect 4250 4333 4253 4416
rect 4218 4323 4237 4326
rect 4250 4283 4253 4326
rect 4202 4213 4213 4216
rect 4154 4163 4173 4166
rect 4130 4133 4133 4146
rect 4114 4123 4133 4126
rect 4098 4053 4117 4056
rect 4026 4003 4029 4016
rect 3954 3973 3965 3976
rect 3906 3953 3917 3956
rect 3882 3923 3885 3936
rect 3906 3906 3909 3953
rect 3882 3803 3885 3906
rect 3906 3903 3917 3906
rect 3914 3836 3917 3903
rect 3914 3833 3925 3836
rect 3890 3813 3893 3826
rect 3906 3813 3909 3826
rect 3898 3803 3909 3806
rect 3898 3743 3901 3803
rect 3866 3646 3869 3736
rect 3906 3726 3909 3796
rect 3922 3776 3925 3833
rect 3890 3676 3893 3726
rect 3858 3643 3869 3646
rect 3874 3673 3893 3676
rect 3902 3723 3909 3726
rect 3914 3773 3925 3776
rect 3858 3606 3861 3643
rect 3866 3613 3869 3626
rect 3858 3603 3869 3606
rect 3874 3603 3877 3673
rect 3902 3666 3905 3723
rect 3914 3676 3917 3773
rect 3938 3763 3941 3956
rect 3954 3953 3957 3973
rect 3962 3903 3965 3926
rect 3914 3673 3925 3676
rect 3902 3663 3909 3666
rect 3810 3446 3813 3563
rect 3826 3533 3829 3556
rect 3850 3523 3853 3546
rect 3810 3443 3821 3446
rect 3802 3393 3805 3406
rect 3810 3343 3813 3426
rect 3818 3353 3821 3443
rect 3826 3326 3829 3506
rect 3834 3446 3837 3466
rect 3834 3443 3845 3446
rect 3674 3203 3677 3246
rect 3634 3123 3637 3136
rect 3610 3113 3621 3116
rect 3578 3083 3589 3086
rect 3554 3003 3557 3026
rect 3578 2973 3581 3083
rect 3554 2916 3557 2936
rect 3554 2913 3565 2916
rect 3542 2853 3549 2856
rect 3522 2813 3533 2816
rect 3514 2713 3517 2726
rect 3506 2693 3513 2696
rect 3510 2636 3513 2693
rect 3522 2643 3525 2806
rect 3530 2636 3533 2813
rect 3542 2806 3545 2853
rect 3562 2846 3565 2913
rect 3602 2903 3605 2926
rect 3554 2843 3565 2846
rect 3542 2803 3549 2806
rect 3538 2673 3541 2786
rect 3506 2633 3513 2636
rect 3522 2633 3533 2636
rect 3506 2616 3509 2633
rect 3498 2613 3509 2616
rect 3506 2533 3509 2606
rect 3522 2536 3525 2633
rect 3530 2576 3533 2626
rect 3546 2623 3549 2803
rect 3554 2776 3557 2843
rect 3602 2813 3605 2836
rect 3618 2806 3621 3113
rect 3642 3003 3645 3016
rect 3650 2923 3653 3016
rect 3666 3013 3669 3126
rect 3674 3113 3677 3136
rect 3682 3123 3685 3206
rect 3690 3013 3693 3156
rect 3698 3133 3701 3166
rect 3714 3163 3717 3216
rect 3722 3203 3725 3323
rect 3738 3213 3741 3236
rect 3770 3213 3773 3236
rect 3706 3103 3709 3126
rect 3722 3056 3725 3196
rect 3762 3193 3765 3206
rect 3730 3123 3733 3136
rect 3746 3113 3749 3136
rect 3762 3133 3765 3156
rect 3770 3126 3773 3206
rect 3754 3123 3773 3126
rect 3718 3053 3725 3056
rect 3658 2993 3661 3006
rect 3674 2973 3677 3006
rect 3658 2916 3661 2936
rect 3706 2933 3709 3016
rect 3718 2996 3721 3053
rect 3718 2993 3725 2996
rect 3738 2993 3741 3016
rect 3714 2916 3717 2976
rect 3658 2913 3669 2916
rect 3650 2866 3653 2886
rect 3578 2793 3581 2806
rect 3602 2803 3621 2806
rect 3646 2863 3653 2866
rect 3646 2806 3649 2863
rect 3666 2836 3669 2913
rect 3658 2833 3669 2836
rect 3706 2913 3717 2916
rect 3658 2813 3661 2833
rect 3706 2826 3709 2913
rect 3706 2823 3717 2826
rect 3646 2803 3653 2806
rect 3554 2773 3565 2776
rect 3562 2696 3565 2773
rect 3578 2716 3581 2736
rect 3554 2693 3565 2696
rect 3574 2713 3581 2716
rect 3554 2673 3557 2693
rect 3574 2636 3577 2713
rect 3574 2633 3581 2636
rect 3546 2583 3549 2606
rect 3570 2603 3573 2616
rect 3530 2573 3549 2576
rect 3522 2533 3541 2536
rect 3490 2366 3493 2526
rect 3514 2523 3533 2526
rect 3498 2423 3501 2436
rect 3506 2373 3509 2406
rect 3490 2363 3501 2366
rect 3474 2353 3481 2356
rect 3458 2343 3469 2346
rect 3466 2316 3469 2343
rect 3458 2313 3469 2316
rect 3458 2226 3461 2313
rect 3478 2306 3481 2353
rect 3490 2313 3493 2336
rect 3498 2326 3501 2363
rect 3506 2333 3509 2346
rect 3514 2336 3517 2446
rect 3522 2413 3525 2426
rect 3530 2403 3533 2523
rect 3538 2443 3541 2533
rect 3514 2333 3525 2336
rect 3538 2326 3541 2416
rect 3498 2323 3509 2326
rect 3478 2303 3485 2306
rect 3458 2223 3469 2226
rect 3418 2083 3429 2086
rect 3410 1933 3413 2056
rect 3418 1936 3421 1986
rect 3426 1943 3429 2083
rect 3442 2033 3445 2186
rect 3450 2013 3453 2126
rect 3458 1996 3461 2206
rect 3466 2186 3469 2223
rect 3474 2203 3477 2216
rect 3482 2213 3485 2303
rect 3514 2226 3517 2326
rect 3530 2323 3541 2326
rect 3506 2223 3517 2226
rect 3490 2193 3493 2206
rect 3466 2183 3473 2186
rect 3450 1993 3461 1996
rect 3418 1933 3429 1936
rect 3426 1923 3429 1933
rect 3394 1913 3405 1916
rect 3402 1846 3405 1913
rect 3418 1893 3421 1916
rect 3450 1856 3453 1993
rect 3470 1986 3473 2183
rect 3482 2103 3485 2126
rect 3498 2123 3501 2216
rect 3506 2203 3509 2223
rect 3506 2123 3509 2166
rect 3522 2133 3525 2246
rect 3530 2213 3533 2323
rect 3538 2196 3541 2256
rect 3534 2193 3541 2196
rect 3498 2083 3501 2106
rect 3534 2066 3537 2193
rect 3534 2063 3541 2066
rect 3482 2023 3501 2026
rect 3466 1983 3473 1986
rect 3450 1853 3461 1856
rect 3394 1843 3405 1846
rect 3378 1763 3381 1806
rect 3362 1626 3365 1726
rect 3370 1713 3373 1746
rect 3378 1696 3381 1736
rect 3386 1733 3389 1816
rect 3394 1733 3397 1843
rect 3402 1806 3405 1826
rect 3434 1813 3437 1836
rect 3402 1803 3413 1806
rect 3410 1756 3413 1803
rect 3402 1753 3413 1756
rect 3346 1623 3365 1626
rect 3374 1693 3381 1696
rect 3374 1626 3377 1693
rect 3374 1623 3381 1626
rect 3346 1586 3349 1623
rect 3290 1523 3309 1526
rect 3290 1403 3293 1523
rect 3298 1403 3301 1436
rect 3290 1303 3293 1326
rect 3282 1283 3289 1286
rect 3258 1093 3269 1096
rect 3210 813 3213 826
rect 3218 803 3221 926
rect 3226 833 3229 926
rect 3250 913 3253 1016
rect 3170 733 3173 746
rect 3194 713 3197 726
rect 3218 713 3221 726
rect 3150 583 3157 586
rect 3130 543 3141 546
rect 3114 433 3117 526
rect 3106 423 3125 426
rect 3098 413 3117 416
rect 3114 403 3117 413
rect 3122 396 3125 423
rect 3114 393 3125 396
rect 3098 333 3101 346
rect 3114 276 3117 393
rect 3122 343 3125 386
rect 3130 333 3133 426
rect 3138 393 3141 543
rect 3150 526 3153 583
rect 3162 543 3165 696
rect 3170 603 3173 616
rect 3178 533 3181 606
rect 3186 593 3189 616
rect 3226 613 3229 816
rect 3242 733 3245 816
rect 3258 783 3261 1093
rect 3274 1016 3277 1256
rect 3286 1196 3289 1283
rect 3282 1193 3289 1196
rect 3282 1173 3285 1193
rect 3298 1173 3301 1336
rect 3306 1323 3309 1336
rect 3314 1333 3317 1406
rect 3322 1396 3325 1586
rect 3342 1583 3349 1586
rect 3330 1503 3333 1546
rect 3342 1516 3345 1583
rect 3354 1523 3357 1616
rect 3362 1603 3365 1616
rect 3342 1513 3349 1516
rect 3346 1403 3349 1513
rect 3362 1433 3365 1536
rect 3370 1523 3373 1606
rect 3378 1506 3381 1623
rect 3374 1503 3381 1506
rect 3322 1393 3333 1396
rect 3314 1313 3317 1326
rect 3306 1203 3309 1216
rect 3314 1213 3317 1236
rect 3322 1206 3325 1393
rect 3374 1376 3377 1503
rect 3386 1386 3389 1686
rect 3394 1633 3397 1726
rect 3402 1613 3405 1753
rect 3410 1643 3413 1736
rect 3418 1713 3421 1726
rect 3426 1696 3429 1736
rect 3418 1693 3429 1696
rect 3418 1613 3421 1693
rect 3394 1543 3397 1606
rect 3402 1583 3405 1596
rect 3394 1413 3397 1526
rect 3402 1516 3405 1536
rect 3434 1516 3437 1726
rect 3442 1683 3445 1826
rect 3458 1816 3461 1853
rect 3466 1823 3469 1983
rect 3474 1923 3477 1946
rect 3482 1866 3485 1936
rect 3490 1933 3493 2016
rect 3498 2006 3501 2023
rect 3498 2003 3509 2006
rect 3506 1946 3509 2003
rect 3538 1966 3541 2063
rect 3498 1943 3509 1946
rect 3530 1963 3541 1966
rect 3498 1923 3501 1943
rect 3482 1863 3501 1866
rect 3450 1813 3461 1816
rect 3466 1813 3477 1816
rect 3450 1673 3453 1813
rect 3458 1803 3477 1806
rect 3482 1783 3485 1856
rect 3458 1733 3461 1746
rect 3458 1713 3461 1726
rect 3402 1513 3413 1516
rect 3410 1436 3413 1513
rect 3402 1433 3413 1436
rect 3426 1513 3437 1516
rect 3402 1413 3405 1433
rect 3386 1383 3393 1386
rect 3374 1373 3381 1376
rect 3314 1203 3325 1206
rect 3282 1103 3285 1136
rect 3290 1096 3293 1156
rect 3330 1153 3333 1246
rect 3338 1206 3341 1256
rect 3362 1243 3365 1346
rect 3370 1333 3373 1356
rect 3378 1253 3381 1373
rect 3390 1296 3393 1383
rect 3402 1323 3405 1406
rect 3426 1343 3429 1513
rect 3442 1486 3445 1656
rect 3450 1613 3453 1626
rect 3458 1556 3461 1646
rect 3474 1633 3477 1726
rect 3490 1663 3493 1806
rect 3498 1803 3501 1863
rect 3506 1806 3509 1826
rect 3514 1813 3517 1926
rect 3530 1846 3533 1963
rect 3530 1843 3541 1846
rect 3530 1813 3533 1826
rect 3506 1803 3517 1806
rect 3506 1653 3509 1796
rect 3514 1643 3517 1803
rect 3538 1793 3541 1843
rect 3546 1833 3549 2573
rect 3570 2536 3573 2586
rect 3578 2566 3581 2633
rect 3586 2583 3589 2716
rect 3602 2706 3605 2803
rect 3650 2736 3653 2803
rect 3666 2773 3669 2816
rect 3618 2713 3621 2736
rect 3650 2733 3661 2736
rect 3602 2703 3621 2706
rect 3578 2563 3597 2566
rect 3570 2533 3581 2536
rect 3554 2403 3557 2516
rect 3554 1933 3557 2366
rect 3562 2296 3565 2526
rect 3578 2466 3581 2533
rect 3570 2463 3581 2466
rect 3570 2406 3573 2463
rect 3594 2446 3597 2563
rect 3578 2443 3597 2446
rect 3578 2413 3581 2443
rect 3570 2403 3581 2406
rect 3594 2403 3597 2416
rect 3602 2403 3605 2426
rect 3578 2333 3581 2403
rect 3610 2373 3613 2416
rect 3562 2293 3569 2296
rect 3566 2196 3569 2293
rect 3578 2243 3581 2326
rect 3602 2323 3605 2346
rect 3562 2193 3569 2196
rect 3562 2173 3565 2193
rect 3578 2123 3581 2196
rect 3594 2193 3597 2216
rect 3586 2133 3589 2146
rect 3602 2133 3605 2316
rect 3618 2226 3621 2703
rect 3642 2683 3645 2726
rect 3642 2656 3645 2676
rect 3638 2653 3645 2656
rect 3626 2533 3629 2616
rect 3638 2556 3641 2653
rect 3658 2636 3661 2733
rect 3698 2723 3701 2806
rect 3714 2803 3717 2823
rect 3722 2786 3725 2993
rect 3746 2873 3749 2926
rect 3754 2856 3757 3056
rect 3778 3053 3781 3326
rect 3818 3323 3829 3326
rect 3818 3266 3821 3323
rect 3818 3263 3829 3266
rect 3826 3243 3829 3263
rect 3842 3246 3845 3443
rect 3858 3363 3861 3576
rect 3866 3553 3869 3603
rect 3882 3563 3885 3616
rect 3890 3613 3893 3626
rect 3874 3353 3877 3536
rect 3906 3533 3909 3663
rect 3890 3523 3909 3526
rect 3890 3403 3893 3523
rect 3922 3516 3925 3673
rect 3946 3603 3949 3726
rect 3970 3636 3973 3766
rect 3970 3633 3989 3636
rect 3954 3533 3957 3556
rect 3914 3513 3925 3516
rect 3978 3513 3981 3526
rect 3914 3463 3917 3513
rect 3906 3403 3909 3416
rect 3930 3393 3933 3416
rect 3986 3413 3989 3633
rect 4010 3606 4013 3826
rect 4018 3803 4021 3926
rect 4026 3923 4029 3936
rect 4034 3903 4037 3986
rect 4042 3953 4045 4006
rect 4058 3933 4061 3966
rect 4034 3833 4037 3876
rect 4058 3813 4061 3836
rect 4066 3813 4069 4006
rect 4090 4003 4093 4016
rect 4114 3976 4117 4053
rect 4146 4046 4149 4156
rect 4142 4043 4149 4046
rect 4106 3973 4117 3976
rect 4074 3923 4077 3936
rect 4090 3906 4093 3926
rect 4106 3923 4109 3973
rect 4114 3913 4117 3956
rect 4130 3933 4133 4006
rect 4142 3956 4145 4043
rect 4170 4036 4173 4163
rect 4202 4106 4205 4126
rect 4154 4033 4173 4036
rect 4194 4103 4205 4106
rect 4142 3953 4149 3956
rect 4146 3933 4149 3953
rect 4154 3933 4157 4033
rect 4194 4026 4197 4103
rect 4194 4023 4205 4026
rect 4138 3923 4157 3926
rect 4074 3823 4077 3836
rect 4018 3723 4021 3746
rect 4042 3723 4045 3806
rect 4082 3803 4085 3906
rect 4090 3903 4097 3906
rect 4094 3836 4097 3903
rect 4090 3833 4097 3836
rect 4090 3733 4093 3833
rect 4106 3813 4109 3826
rect 4098 3793 4101 3806
rect 4106 3803 4117 3806
rect 4122 3803 4125 3816
rect 4114 3733 4117 3756
rect 4114 3713 4117 3726
rect 4034 3613 4037 3626
rect 4106 3606 4109 3656
rect 4114 3613 4117 3646
rect 4122 3613 4125 3736
rect 4130 3733 4133 3746
rect 4138 3713 4141 3726
rect 4010 3603 4037 3606
rect 4106 3603 4117 3606
rect 4130 3603 4133 3626
rect 4018 3413 4021 3426
rect 3874 3333 3877 3346
rect 3834 3243 3845 3246
rect 3786 3203 3789 3216
rect 3810 3213 3813 3226
rect 3794 3036 3797 3136
rect 3818 3113 3821 3126
rect 3826 3076 3829 3236
rect 3786 3033 3797 3036
rect 3818 3073 3829 3076
rect 3786 3003 3789 3033
rect 3786 2926 3789 2996
rect 3818 2946 3821 3073
rect 3834 2993 3837 3243
rect 3842 3203 3845 3226
rect 3898 3216 3901 3356
rect 4034 3336 4037 3603
rect 4114 3583 4117 3603
rect 4138 3543 4141 3646
rect 4146 3603 4149 3806
rect 4154 3706 4157 3816
rect 4162 3803 4165 3936
rect 4170 3933 4173 4016
rect 4202 4003 4205 4023
rect 4210 3906 4213 4213
rect 4218 4196 4221 4276
rect 4242 4213 4245 4226
rect 4258 4196 4261 4216
rect 4218 4193 4229 4196
rect 4226 4126 4229 4193
rect 4218 4123 4229 4126
rect 4250 4193 4261 4196
rect 4218 4006 4221 4123
rect 4226 4013 4229 4106
rect 4250 4056 4253 4193
rect 4266 4173 4269 4336
rect 4290 4316 4293 4336
rect 4298 4333 4301 4436
rect 4306 4333 4309 4356
rect 4314 4333 4317 4366
rect 4326 4356 4329 4443
rect 4322 4353 4329 4356
rect 4282 4313 4293 4316
rect 4282 4266 4285 4313
rect 4282 4263 4293 4266
rect 4274 4203 4277 4246
rect 4290 4233 4293 4263
rect 4298 4243 4301 4326
rect 4322 4323 4325 4353
rect 4306 4233 4309 4256
rect 4242 4053 4253 4056
rect 4218 4003 4229 4006
rect 4202 3903 4213 3906
rect 4170 3813 4173 3836
rect 4202 3826 4205 3903
rect 4178 3803 4181 3826
rect 4186 3823 4205 3826
rect 4154 3703 4165 3706
rect 4162 3646 4165 3703
rect 4154 3643 4165 3646
rect 4154 3596 4157 3643
rect 4146 3593 4157 3596
rect 4074 3493 4077 3526
rect 4130 3523 4141 3526
rect 4066 3433 4069 3476
rect 4030 3333 4037 3336
rect 3922 3286 3925 3326
rect 3978 3306 3981 3326
rect 3970 3303 3981 3306
rect 3922 3283 3933 3286
rect 3818 2943 3829 2946
rect 3746 2853 3757 2856
rect 3714 2783 3725 2786
rect 3714 2726 3717 2783
rect 3714 2723 3725 2726
rect 3650 2633 3661 2636
rect 3638 2553 3645 2556
rect 3634 2523 3637 2536
rect 3626 2373 3629 2416
rect 3642 2323 3645 2553
rect 3650 2503 3653 2633
rect 3666 2523 3669 2616
rect 3690 2613 3693 2676
rect 3698 2603 3701 2626
rect 3706 2613 3717 2616
rect 3722 2613 3725 2723
rect 3674 2523 3677 2546
rect 3658 2356 3661 2406
rect 3654 2353 3661 2356
rect 3614 2223 3621 2226
rect 3562 2093 3565 2116
rect 3562 1993 3565 2016
rect 3586 1983 3589 2006
rect 3602 2003 3605 2126
rect 3614 2116 3617 2223
rect 3626 2123 3629 2216
rect 3634 2123 3637 2206
rect 3642 2203 3645 2246
rect 3654 2236 3657 2353
rect 3654 2233 3661 2236
rect 3658 2203 3661 2233
rect 3666 2186 3669 2346
rect 3682 2293 3685 2326
rect 3658 2183 3669 2186
rect 3614 2113 3621 2116
rect 3618 2033 3621 2113
rect 3562 1916 3565 1936
rect 3578 1933 3581 1946
rect 3602 1923 3621 1926
rect 3562 1913 3573 1916
rect 3570 1846 3573 1913
rect 3562 1843 3573 1846
rect 3562 1823 3565 1843
rect 3586 1813 3589 1826
rect 3626 1823 3629 1936
rect 3642 1933 3645 2136
rect 3658 2036 3661 2183
rect 3674 2166 3677 2206
rect 3690 2203 3693 2316
rect 3714 2233 3717 2536
rect 3722 2523 3725 2546
rect 3730 2536 3733 2796
rect 3746 2736 3749 2853
rect 3762 2746 3765 2926
rect 3786 2923 3797 2926
rect 3826 2923 3829 2943
rect 3770 2896 3773 2916
rect 3770 2893 3781 2896
rect 3778 2836 3781 2893
rect 3770 2833 3781 2836
rect 3770 2813 3773 2833
rect 3762 2743 3769 2746
rect 3746 2733 3757 2736
rect 3738 2676 3741 2716
rect 3746 2693 3749 2706
rect 3738 2673 3745 2676
rect 3742 2546 3745 2673
rect 3754 2576 3757 2733
rect 3766 2696 3769 2743
rect 3762 2693 3769 2696
rect 3762 2673 3765 2693
rect 3762 2593 3765 2606
rect 3770 2603 3773 2666
rect 3778 2613 3781 2816
rect 3794 2796 3797 2923
rect 3834 2906 3837 2926
rect 3830 2903 3837 2906
rect 3830 2836 3833 2903
rect 3818 2813 3821 2836
rect 3830 2833 3837 2836
rect 3786 2793 3797 2796
rect 3786 2713 3789 2793
rect 3786 2693 3789 2706
rect 3754 2573 3765 2576
rect 3742 2543 3749 2546
rect 3730 2533 3741 2536
rect 3730 2413 3733 2426
rect 3738 2343 3741 2533
rect 3738 2313 3741 2326
rect 3746 2253 3749 2543
rect 3762 2466 3765 2573
rect 3786 2563 3789 2606
rect 3794 2583 3797 2626
rect 3802 2573 3805 2776
rect 3826 2723 3829 2806
rect 3834 2753 3837 2833
rect 3834 2686 3837 2726
rect 3826 2683 3837 2686
rect 3810 2593 3813 2616
rect 3826 2586 3829 2683
rect 3842 2666 3845 3166
rect 3858 3163 3861 3216
rect 3866 3203 3877 3206
rect 3874 3113 3877 3203
rect 3874 3066 3877 3086
rect 3850 3046 3853 3066
rect 3870 3063 3877 3066
rect 3850 3043 3861 3046
rect 3858 2996 3861 3043
rect 3850 2993 3861 2996
rect 3850 2903 3853 2993
rect 3858 2923 3861 2976
rect 3870 2926 3873 3063
rect 3870 2923 3877 2926
rect 3850 2813 3853 2836
rect 3838 2663 3845 2666
rect 3838 2606 3841 2663
rect 3838 2603 3845 2606
rect 3826 2583 3837 2586
rect 3754 2463 3765 2466
rect 3754 2386 3757 2463
rect 3794 2426 3797 2556
rect 3818 2523 3821 2566
rect 3826 2516 3829 2556
rect 3818 2513 3829 2516
rect 3794 2423 3813 2426
rect 3778 2403 3781 2416
rect 3754 2383 3761 2386
rect 3758 2266 3761 2383
rect 3794 2336 3797 2416
rect 3786 2333 3797 2336
rect 3754 2263 3761 2266
rect 3754 2236 3757 2263
rect 3698 2213 3701 2226
rect 3714 2213 3717 2226
rect 3706 2173 3709 2206
rect 3670 2163 3677 2166
rect 3670 2086 3673 2163
rect 3690 2123 3693 2146
rect 3738 2133 3741 2236
rect 3750 2233 3757 2236
rect 3750 2166 3753 2233
rect 3750 2163 3757 2166
rect 3670 2083 3677 2086
rect 3658 2033 3669 2036
rect 3650 2003 3653 2016
rect 3658 1993 3661 2006
rect 3666 1983 3669 2033
rect 3674 2016 3677 2083
rect 3674 2013 3685 2016
rect 3698 2013 3701 2106
rect 3674 1973 3677 2006
rect 3682 1933 3685 2013
rect 3714 1983 3717 2006
rect 3610 1793 3613 1806
rect 3642 1793 3645 1926
rect 3690 1913 3693 1926
rect 3698 1856 3701 1936
rect 3714 1933 3717 1976
rect 3722 1926 3725 1936
rect 3706 1923 3725 1926
rect 3730 1903 3733 1926
rect 3690 1853 3701 1856
rect 3690 1813 3693 1853
rect 3738 1813 3741 1936
rect 3754 1853 3757 2163
rect 3762 2133 3765 2246
rect 3770 2203 3773 2286
rect 3786 2273 3789 2333
rect 3794 2283 3797 2326
rect 3786 2203 3789 2226
rect 3762 2103 3765 2126
rect 3786 2026 3789 2196
rect 3810 2193 3813 2423
rect 3818 2413 3821 2513
rect 3834 2496 3837 2583
rect 3830 2493 3837 2496
rect 3830 2426 3833 2493
rect 3830 2423 3837 2426
rect 3834 2333 3837 2423
rect 3842 2363 3845 2603
rect 3850 2573 3853 2806
rect 3858 2603 3861 2616
rect 3874 2593 3877 2923
rect 3882 2876 3885 3216
rect 3898 3213 3905 3216
rect 3890 3183 3893 3206
rect 3890 3123 3893 3136
rect 3902 3106 3905 3213
rect 3914 3133 3917 3206
rect 3922 3203 3925 3216
rect 3930 3203 3933 3283
rect 3970 3246 3973 3303
rect 3970 3243 3981 3246
rect 3938 3193 3941 3216
rect 3954 3213 3957 3226
rect 3978 3193 3981 3243
rect 3986 3183 3989 3206
rect 3994 3203 3997 3326
rect 4030 3276 4033 3333
rect 4042 3303 4045 3326
rect 4026 3273 4033 3276
rect 4026 3146 4029 3273
rect 4026 3143 4037 3146
rect 3890 2923 3893 3106
rect 3898 3103 3905 3106
rect 3898 3083 3901 3103
rect 3906 3003 3909 3036
rect 3946 3033 3949 3136
rect 3898 2893 3901 2936
rect 3882 2873 3893 2876
rect 3890 2646 3893 2873
rect 3914 2796 3917 2926
rect 3930 2916 3933 3016
rect 3938 2933 3941 3006
rect 3970 2976 3973 3126
rect 3986 3026 3989 3116
rect 4026 3106 4029 3126
rect 4018 3103 4029 3106
rect 4018 3036 4021 3103
rect 4034 3046 4037 3143
rect 4042 3133 4045 3186
rect 4050 3063 4053 3426
rect 4082 3423 4085 3516
rect 4122 3483 4125 3506
rect 4146 3456 4149 3593
rect 4170 3536 4173 3626
rect 4186 3616 4189 3823
rect 4210 3786 4213 3816
rect 4226 3803 4229 4003
rect 4242 3996 4245 4053
rect 4250 4003 4253 4026
rect 4242 3993 4253 3996
rect 4234 3903 4237 3926
rect 4250 3833 4253 3993
rect 4250 3793 4253 3816
rect 4210 3783 4221 3786
rect 4194 3733 4205 3736
rect 4194 3633 4197 3666
rect 4202 3623 4205 3726
rect 4210 3713 4213 3736
rect 4210 3616 4213 3626
rect 4186 3613 4197 3616
rect 4202 3613 4213 3616
rect 4166 3533 4173 3536
rect 4186 3533 4189 3546
rect 4154 3503 4157 3516
rect 4166 3456 4169 3533
rect 4138 3453 4149 3456
rect 4138 3446 4141 3453
rect 4122 3443 4141 3446
rect 4122 3376 4125 3443
rect 4138 3386 4141 3436
rect 4146 3413 4149 3446
rect 4154 3433 4157 3456
rect 4166 3453 4173 3456
rect 4162 3413 4165 3436
rect 4138 3383 4145 3386
rect 4122 3373 4133 3376
rect 4074 3216 4077 3346
rect 4106 3333 4109 3346
rect 4070 3213 4077 3216
rect 4058 3143 4061 3186
rect 4070 3146 4073 3213
rect 4066 3143 4073 3146
rect 4066 3046 4069 3143
rect 4074 3106 4077 3136
rect 4082 3123 4085 3206
rect 4090 3133 4093 3306
rect 4130 3276 4133 3373
rect 4122 3273 4133 3276
rect 4142 3276 4145 3383
rect 4154 3303 4157 3326
rect 4142 3273 4149 3276
rect 4098 3113 4101 3206
rect 4122 3186 4125 3273
rect 4122 3183 4133 3186
rect 4106 3133 4109 3146
rect 4114 3123 4117 3166
rect 4122 3123 4125 3136
rect 4074 3103 4085 3106
rect 4034 3043 4045 3046
rect 4018 3033 4029 3036
rect 3986 3023 3993 3026
rect 3954 2973 3973 2976
rect 3954 2933 3957 2973
rect 3962 2923 3965 2936
rect 3922 2903 3925 2916
rect 3930 2913 3949 2916
rect 3930 2806 3933 2846
rect 3922 2803 3933 2806
rect 3946 2803 3949 2913
rect 3954 2813 3973 2816
rect 3906 2793 3917 2796
rect 3962 2796 3965 2806
rect 3970 2803 3973 2813
rect 3978 2796 3981 3016
rect 3990 2836 3993 3023
rect 3986 2833 3993 2836
rect 3986 2813 3989 2833
rect 3962 2793 3981 2796
rect 3906 2716 3909 2793
rect 3922 2723 3925 2756
rect 3962 2746 3965 2793
rect 3954 2743 3965 2746
rect 3906 2713 3917 2716
rect 3882 2643 3893 2646
rect 3882 2533 3885 2643
rect 3890 2476 3893 2616
rect 3898 2603 3901 2626
rect 3906 2603 3909 2616
rect 3914 2613 3917 2713
rect 3930 2693 3933 2716
rect 3954 2696 3957 2743
rect 3978 2703 3981 2736
rect 3986 2703 3989 2726
rect 3954 2693 3965 2696
rect 3962 2636 3965 2693
rect 3954 2633 3965 2636
rect 3898 2523 3901 2586
rect 3906 2496 3909 2596
rect 3922 2593 3925 2606
rect 3930 2603 3933 2616
rect 3946 2613 3949 2626
rect 3954 2536 3957 2633
rect 3994 2593 3997 2616
rect 4002 2583 4005 2986
rect 4010 2933 4013 3016
rect 4018 2933 4021 3016
rect 4026 3003 4029 3033
rect 4042 2996 4045 3043
rect 4062 3043 4069 3046
rect 4062 2996 4065 3043
rect 4082 3036 4085 3103
rect 4034 2993 4045 2996
rect 4058 2993 4065 2996
rect 4074 3033 4085 3036
rect 4018 2803 4021 2926
rect 4026 2786 4029 2816
rect 4034 2796 4037 2993
rect 4058 2946 4061 2993
rect 4050 2943 4061 2946
rect 4050 2846 4053 2943
rect 4050 2843 4061 2846
rect 4042 2813 4045 2826
rect 4034 2793 4045 2796
rect 4018 2783 4029 2786
rect 4018 2736 4021 2783
rect 4018 2733 4029 2736
rect 4026 2713 4029 2733
rect 4042 2716 4045 2793
rect 4058 2773 4061 2843
rect 4066 2716 4069 2936
rect 4074 2933 4077 3033
rect 4098 2936 4101 3096
rect 4106 3003 4109 3026
rect 4090 2933 4101 2936
rect 4090 2916 4093 2933
rect 4086 2913 4093 2916
rect 4074 2803 4077 2856
rect 4086 2846 4089 2913
rect 4098 2853 4101 2926
rect 4106 2856 4109 2936
rect 4114 2933 4117 3016
rect 4130 3013 4133 3183
rect 4146 3146 4149 3273
rect 4170 3213 4173 3453
rect 4138 3143 4149 3146
rect 4138 3093 4141 3143
rect 4178 3133 4181 3526
rect 4194 3436 4197 3613
rect 4186 3433 4197 3436
rect 4218 3433 4221 3783
rect 4226 3733 4229 3756
rect 4226 3583 4229 3606
rect 4234 3503 4237 3526
rect 4186 3406 4189 3433
rect 4194 3423 4221 3426
rect 4218 3413 4221 3423
rect 4234 3413 4237 3426
rect 4242 3416 4245 3746
rect 4258 3613 4261 4016
rect 4266 4003 4269 4126
rect 4282 4016 4285 4226
rect 4298 4223 4309 4226
rect 4306 4203 4309 4216
rect 4298 4096 4301 4116
rect 4298 4093 4309 4096
rect 4306 4046 4309 4093
rect 4274 4013 4285 4016
rect 4298 4043 4309 4046
rect 4266 3743 4269 3836
rect 4266 3713 4269 3736
rect 4274 3616 4277 4013
rect 4298 4003 4301 4043
rect 4306 4013 4309 4026
rect 4282 3913 4285 3936
rect 4290 3933 4293 3956
rect 4306 3933 4309 4006
rect 4314 3913 4317 3926
rect 4322 3836 4325 4006
rect 4330 3986 4333 4336
rect 4338 4333 4341 4416
rect 4346 4363 4349 4466
rect 4346 4323 4349 4346
rect 4362 4333 4365 4546
rect 4378 4513 4381 4536
rect 4394 4533 4397 4566
rect 4418 4533 4421 4606
rect 4434 4533 4437 4546
rect 4442 4526 4445 4616
rect 4450 4563 4453 4606
rect 4482 4603 4485 4616
rect 4490 4566 4493 4606
rect 4498 4573 4501 4616
rect 4522 4583 4525 4606
rect 4490 4563 4509 4566
rect 4394 4496 4397 4526
rect 4410 4523 4421 4526
rect 4426 4523 4445 4526
rect 4386 4493 4397 4496
rect 4386 4446 4389 4493
rect 4386 4443 4397 4446
rect 4394 4423 4397 4443
rect 4378 4413 4397 4416
rect 4378 4333 4381 4413
rect 4410 4396 4413 4506
rect 4426 4456 4429 4523
rect 4418 4453 4429 4456
rect 4418 4403 4421 4453
rect 4426 4413 4429 4446
rect 4402 4393 4413 4396
rect 4402 4336 4405 4393
rect 4402 4333 4413 4336
rect 4418 4333 4421 4356
rect 4442 4333 4445 4426
rect 4458 4413 4461 4526
rect 4482 4426 4485 4546
rect 4506 4523 4509 4563
rect 4570 4543 4573 4606
rect 4466 4423 4485 4426
rect 4450 4333 4453 4346
rect 4362 4313 4365 4326
rect 4330 3983 4349 3986
rect 4346 3933 4349 3983
rect 4354 3966 4357 4296
rect 4386 4263 4389 4326
rect 4410 4313 4413 4333
rect 4378 4213 4381 4236
rect 4426 4196 4429 4326
rect 4458 4323 4461 4386
rect 4466 4373 4469 4423
rect 4474 4403 4477 4416
rect 4482 4393 4485 4406
rect 4474 4313 4477 4326
rect 4450 4213 4453 4246
rect 4426 4193 4437 4196
rect 4378 4113 4381 4126
rect 4434 4086 4437 4193
rect 4458 4136 4461 4236
rect 4426 4083 4437 4086
rect 4450 4133 4461 4136
rect 4426 4056 4429 4083
rect 4426 4053 4437 4056
rect 4378 4003 4381 4016
rect 4434 3976 4437 4053
rect 4426 3973 4437 3976
rect 4354 3963 4373 3966
rect 4370 3946 4373 3963
rect 4370 3943 4377 3946
rect 4374 3896 4377 3943
rect 4370 3893 4377 3896
rect 4306 3833 4325 3836
rect 4306 3756 4309 3833
rect 4322 3813 4325 3826
rect 4306 3753 4317 3756
rect 4282 3733 4285 3746
rect 4290 3726 4293 3736
rect 4290 3723 4309 3726
rect 4314 3706 4317 3753
rect 4330 3726 4333 3846
rect 4354 3796 4357 3816
rect 4370 3806 4373 3893
rect 4386 3813 4389 3896
rect 4346 3793 4357 3796
rect 4362 3793 4365 3806
rect 4370 3803 4381 3806
rect 4394 3803 4397 3926
rect 4402 3813 4405 3826
rect 4346 3746 4349 3793
rect 4346 3743 4357 3746
rect 4330 3723 4341 3726
rect 4310 3703 4317 3706
rect 4266 3613 4277 3616
rect 4266 3596 4269 3613
rect 4262 3593 4269 3596
rect 4262 3526 4265 3593
rect 4274 3533 4277 3606
rect 4250 3423 4253 3526
rect 4262 3523 4269 3526
rect 4242 3413 4253 3416
rect 4186 3403 4197 3406
rect 4194 3326 4197 3403
rect 4190 3323 4197 3326
rect 4190 3156 4193 3323
rect 4190 3153 4197 3156
rect 4186 3133 4189 3146
rect 4122 2993 4125 3006
rect 4106 2853 4117 2856
rect 4086 2843 4093 2846
rect 4090 2813 4093 2843
rect 4114 2813 4117 2853
rect 4074 2723 4077 2796
rect 4090 2773 4093 2806
rect 4122 2753 4125 2926
rect 4130 2803 4133 2936
rect 4146 2856 4149 3126
rect 4162 2993 4165 3126
rect 4170 3096 4173 3126
rect 4170 3093 4181 3096
rect 4178 3036 4181 3093
rect 4170 3033 4181 3036
rect 4194 3033 4197 3153
rect 4202 3133 4205 3306
rect 4210 3123 4213 3406
rect 4250 3396 4253 3413
rect 4242 3393 4253 3396
rect 4242 3266 4245 3393
rect 4242 3263 4253 3266
rect 4250 3246 4253 3263
rect 4250 3243 4257 3246
rect 4226 3136 4229 3206
rect 4254 3196 4257 3243
rect 4250 3193 4257 3196
rect 4218 3046 4221 3136
rect 4226 3133 4237 3136
rect 4210 3043 4221 3046
rect 4162 2923 4165 2936
rect 4170 2923 4173 3033
rect 4202 3013 4205 3026
rect 4194 2993 4197 3006
rect 4210 2946 4213 3043
rect 4194 2943 4213 2946
rect 4146 2853 4165 2856
rect 4034 2713 4045 2716
rect 4034 2693 4037 2713
rect 4058 2633 4061 2716
rect 4066 2713 4077 2716
rect 4066 2623 4069 2696
rect 4074 2653 4077 2706
rect 4082 2633 4093 2636
rect 3922 2523 3925 2536
rect 3954 2533 3965 2536
rect 3906 2493 3913 2496
rect 3890 2473 3901 2476
rect 3874 2413 3877 2436
rect 3890 2406 3893 2416
rect 3898 2413 3901 2473
rect 3910 2406 3913 2493
rect 3858 2393 3861 2406
rect 3866 2403 3893 2406
rect 3906 2403 3913 2406
rect 3922 2403 3925 2426
rect 3930 2403 3933 2456
rect 3946 2403 3949 2526
rect 3962 2456 3965 2533
rect 3954 2453 3965 2456
rect 3954 2433 3957 2453
rect 3954 2413 3973 2416
rect 3954 2403 3957 2413
rect 3826 2233 3829 2326
rect 3850 2323 3853 2336
rect 3858 2306 3861 2326
rect 3854 2303 3861 2306
rect 3834 2193 3837 2216
rect 3854 2176 3857 2303
rect 3866 2196 3869 2403
rect 3906 2346 3909 2403
rect 3890 2326 3893 2346
rect 3906 2343 3925 2346
rect 3874 2303 3877 2326
rect 3882 2213 3885 2326
rect 3890 2323 3897 2326
rect 3894 2206 3897 2323
rect 3890 2203 3897 2206
rect 3866 2193 3877 2196
rect 3854 2173 3861 2176
rect 3858 2153 3861 2173
rect 3762 2013 3765 2026
rect 3786 2023 3797 2026
rect 3810 2023 3813 2136
rect 3818 2123 3837 2126
rect 3842 2123 3845 2136
rect 3818 2106 3821 2123
rect 3858 2106 3861 2136
rect 3874 2106 3877 2193
rect 3890 2133 3893 2203
rect 3818 2103 3829 2106
rect 3778 1923 3781 2016
rect 3794 1946 3797 2023
rect 3826 2016 3829 2103
rect 3850 2103 3861 2106
rect 3866 2103 3877 2106
rect 3890 2103 3893 2126
rect 3850 2036 3853 2103
rect 3866 2086 3869 2103
rect 3866 2083 3877 2086
rect 3850 2033 3861 2036
rect 3786 1943 3797 1946
rect 3818 2013 3829 2016
rect 3858 2013 3861 2033
rect 3786 1923 3789 1943
rect 3818 1933 3821 2013
rect 3874 2006 3877 2083
rect 3866 2003 3877 2006
rect 3794 1853 3797 1926
rect 3834 1923 3837 1986
rect 3842 1933 3845 1946
rect 3850 1893 3853 1926
rect 3866 1903 3869 2003
rect 3906 1956 3909 2343
rect 3914 2313 3917 2336
rect 3922 2333 3925 2343
rect 3922 2263 3925 2326
rect 3930 2323 3933 2366
rect 3938 2333 3941 2396
rect 3954 2333 3957 2356
rect 3978 2343 3981 2436
rect 3986 2406 3989 2526
rect 4002 2486 4005 2526
rect 4010 2506 4013 2526
rect 4042 2523 4045 2616
rect 4106 2603 4109 2646
rect 4130 2636 4133 2776
rect 4114 2633 4133 2636
rect 4114 2596 4117 2633
rect 4122 2603 4125 2626
rect 4138 2616 4141 2636
rect 4138 2613 4149 2616
rect 4106 2593 4117 2596
rect 4082 2523 4085 2536
rect 4010 2503 4021 2506
rect 3994 2483 4005 2486
rect 3994 2413 3997 2483
rect 4018 2436 4021 2503
rect 4106 2463 4109 2593
rect 4122 2533 4125 2576
rect 4130 2496 4133 2606
rect 4146 2556 4149 2613
rect 4122 2493 4133 2496
rect 4138 2553 4149 2556
rect 4010 2433 4021 2436
rect 4002 2413 4005 2426
rect 3986 2403 3997 2406
rect 4010 2403 4013 2433
rect 3946 2313 3949 2326
rect 3962 2313 3965 2326
rect 3938 2203 3941 2216
rect 3954 2213 3957 2226
rect 3970 2213 3973 2236
rect 3946 2193 3949 2206
rect 3938 2133 3941 2146
rect 3946 2133 3957 2136
rect 3994 2133 3997 2403
rect 4018 2333 4021 2416
rect 4050 2393 4053 2416
rect 4098 2386 4101 2446
rect 4122 2416 4125 2493
rect 4138 2443 4141 2553
rect 4146 2533 4157 2536
rect 4162 2533 4165 2853
rect 4178 2833 4181 2936
rect 4194 2933 4197 2943
rect 4202 2926 4205 2936
rect 4186 2923 4205 2926
rect 4194 2856 4197 2876
rect 4190 2853 4197 2856
rect 4190 2786 4193 2853
rect 4202 2813 4205 2856
rect 4190 2783 4197 2786
rect 4194 2766 4197 2783
rect 4194 2763 4205 2766
rect 4178 2713 4181 2726
rect 4178 2536 4181 2696
rect 4170 2533 4181 2536
rect 4146 2506 4149 2526
rect 4146 2503 4157 2506
rect 4154 2446 4157 2503
rect 4170 2453 4173 2533
rect 4146 2443 4157 2446
rect 4146 2423 4149 2443
rect 4122 2413 4133 2416
rect 4098 2383 4109 2386
rect 4098 2346 4101 2366
rect 4090 2343 4101 2346
rect 4106 2343 4109 2383
rect 4090 2286 4093 2343
rect 4090 2283 4101 2286
rect 4010 2173 4013 2206
rect 4050 2203 4053 2226
rect 4058 2163 4061 2216
rect 4074 2213 4077 2266
rect 4082 2203 4085 2216
rect 3930 2123 3941 2126
rect 3898 1953 3909 1956
rect 3874 1913 3877 1926
rect 3898 1913 3901 1936
rect 3906 1933 3909 1953
rect 3914 1923 3917 1956
rect 3922 1933 3925 2006
rect 3938 1933 3941 2066
rect 3946 1943 3949 2126
rect 4018 2123 4021 2146
rect 4090 2103 4093 2126
rect 3962 1933 3965 2016
rect 4002 2003 4005 2016
rect 4082 2013 4085 2096
rect 4050 1976 4053 2006
rect 3930 1913 3933 1926
rect 3946 1913 3949 1926
rect 3970 1826 3973 1976
rect 4042 1973 4053 1976
rect 4042 1923 4045 1973
rect 4066 1933 4069 2006
rect 4074 1993 4077 2006
rect 4098 1983 4101 2283
rect 4114 2246 4117 2396
rect 4130 2363 4133 2413
rect 4138 2366 4141 2406
rect 4146 2373 4149 2416
rect 4138 2363 4149 2366
rect 4130 2333 4133 2346
rect 4146 2343 4149 2363
rect 4110 2243 4117 2246
rect 4110 2196 4113 2243
rect 4122 2203 4125 2236
rect 4110 2193 4117 2196
rect 4106 2063 4109 2136
rect 4114 2133 4117 2193
rect 4130 2163 4133 2326
rect 4154 2323 4157 2406
rect 4162 2233 4165 2416
rect 4170 2353 4173 2406
rect 4146 2193 4149 2206
rect 4154 2146 4157 2226
rect 4162 2173 4165 2206
rect 4154 2143 4165 2146
rect 4106 1993 4109 2016
rect 4114 2003 4117 2106
rect 4130 2013 4133 2126
rect 4138 2076 4141 2136
rect 4146 2096 4149 2136
rect 4162 2123 4165 2143
rect 4170 2113 4173 2166
rect 4178 2133 4181 2526
rect 4194 2523 4197 2756
rect 4202 2633 4205 2763
rect 4202 2603 4205 2626
rect 4210 2576 4213 2943
rect 4218 2823 4221 3036
rect 4226 3023 4229 3126
rect 4234 3116 4237 3133
rect 4234 3113 4241 3116
rect 4218 2603 4221 2746
rect 4226 2596 4229 3016
rect 4238 2896 4241 3113
rect 4250 2983 4253 3193
rect 4266 3013 4269 3523
rect 4282 3413 4285 3616
rect 4298 3613 4301 3636
rect 4310 3626 4313 3703
rect 4310 3623 4317 3626
rect 4314 3603 4317 3623
rect 4322 3603 4325 3716
rect 4338 3626 4341 3723
rect 4330 3623 4341 3626
rect 4330 3566 4333 3623
rect 4322 3563 4333 3566
rect 4322 3546 4325 3563
rect 4318 3543 4325 3546
rect 4274 3323 4277 3336
rect 4282 3256 4285 3366
rect 4290 3283 4293 3406
rect 4306 3403 4309 3526
rect 4318 3486 4321 3543
rect 4338 3523 4341 3536
rect 4318 3483 4325 3486
rect 4322 3416 4325 3483
rect 4322 3413 4333 3416
rect 4314 3333 4317 3406
rect 4330 3356 4333 3413
rect 4346 3363 4349 3606
rect 4354 3553 4357 3743
rect 4362 3733 4365 3756
rect 4378 3666 4381 3803
rect 4402 3723 4405 3746
rect 4370 3663 4381 3666
rect 4362 3486 4365 3576
rect 4370 3543 4373 3663
rect 4378 3603 4381 3656
rect 4386 3613 4397 3616
rect 4402 3556 4405 3606
rect 4410 3603 4413 3926
rect 4426 3766 4429 3973
rect 4450 3946 4453 4133
rect 4466 4023 4469 4126
rect 4450 3943 4461 3946
rect 4434 3813 4437 3826
rect 4450 3803 4453 3926
rect 4458 3923 4461 3943
rect 4466 3913 4469 4016
rect 4474 3893 4477 4216
rect 4490 4213 4493 4416
rect 4498 4393 4501 4406
rect 4506 4333 4509 4426
rect 4482 4173 4485 4206
rect 4498 4203 4501 4216
rect 4506 4196 4509 4226
rect 4514 4203 4517 4406
rect 4538 4383 4541 4406
rect 4562 4393 4565 4416
rect 4578 4413 4581 4576
rect 4586 4533 4589 4556
rect 4594 4523 4597 4606
rect 4602 4533 4605 4616
rect 4618 4533 4621 4586
rect 4610 4513 4613 4526
rect 4626 4513 4629 4526
rect 4634 4413 4637 4426
rect 4642 4416 4645 4536
rect 4650 4533 4653 4616
rect 4666 4463 4669 4536
rect 4674 4523 4677 4536
rect 4682 4533 4685 4606
rect 4698 4556 4701 4606
rect 4722 4603 4725 4616
rect 4698 4553 4717 4556
rect 4690 4513 4693 4526
rect 4698 4456 4701 4546
rect 4714 4466 4717 4553
rect 4778 4526 4781 4616
rect 4674 4453 4701 4456
rect 4706 4463 4717 4466
rect 4770 4523 4781 4526
rect 4642 4413 4653 4416
rect 4530 4296 4533 4316
rect 4530 4293 4541 4296
rect 4538 4236 4541 4293
rect 4530 4233 4541 4236
rect 4522 4196 4525 4206
rect 4506 4193 4525 4196
rect 4482 3986 4485 4116
rect 4498 4103 4501 4166
rect 4506 4113 4509 4126
rect 4514 4103 4517 4116
rect 4530 4093 4533 4233
rect 4570 4216 4573 4386
rect 4618 4366 4621 4406
rect 4634 4403 4645 4406
rect 4610 4363 4621 4366
rect 4546 4203 4549 4216
rect 4562 4213 4573 4216
rect 4578 4213 4581 4226
rect 4594 4213 4597 4326
rect 4610 4286 4613 4363
rect 4650 4336 4653 4413
rect 4658 4393 4661 4406
rect 4666 4343 4669 4416
rect 4674 4383 4677 4453
rect 4690 4366 4693 4446
rect 4706 4443 4709 4463
rect 4770 4436 4773 4523
rect 4770 4433 4781 4436
rect 4714 4393 4717 4416
rect 4682 4363 4693 4366
rect 4650 4333 4669 4336
rect 4610 4283 4621 4286
rect 4618 4226 4621 4283
rect 4618 4223 4629 4226
rect 4554 4193 4557 4206
rect 4490 4003 4493 4016
rect 4514 4013 4517 4056
rect 4554 4053 4557 4136
rect 4506 3993 4509 4006
rect 4482 3983 4489 3986
rect 4486 3896 4489 3983
rect 4522 3976 4525 4006
rect 4522 3973 4533 3976
rect 4482 3893 4489 3896
rect 4482 3876 4485 3893
rect 4474 3873 4485 3876
rect 4474 3776 4477 3873
rect 4474 3773 4485 3776
rect 4422 3763 4429 3766
rect 4422 3686 4425 3763
rect 4482 3756 4485 3773
rect 4458 3723 4461 3756
rect 4482 3753 4489 3756
rect 4474 3706 4477 3726
rect 4470 3703 4477 3706
rect 4422 3683 4429 3686
rect 4418 3603 4421 3616
rect 4426 3593 4429 3683
rect 4442 3613 4445 3646
rect 4470 3636 4473 3703
rect 4486 3696 4489 3753
rect 4482 3693 4489 3696
rect 4470 3633 4477 3636
rect 4482 3633 4485 3693
rect 4434 3583 4437 3606
rect 4450 3603 4453 3616
rect 4458 3613 4461 3626
rect 4402 3553 4409 3556
rect 4386 3533 4389 3546
rect 4406 3506 4409 3553
rect 4426 3533 4429 3546
rect 4402 3503 4409 3506
rect 4362 3483 4381 3486
rect 4322 3353 4333 3356
rect 4322 3326 4325 3353
rect 4306 3323 4325 3326
rect 4330 3323 4333 3336
rect 4354 3333 4357 3386
rect 4306 3306 4309 3323
rect 4306 3303 4317 3306
rect 4282 3253 4293 3256
rect 4290 3236 4293 3253
rect 4290 3233 4297 3236
rect 4274 3193 4277 3216
rect 4294 3176 4297 3233
rect 4314 3226 4317 3303
rect 4290 3173 4297 3176
rect 4306 3223 4317 3226
rect 4274 3103 4277 3126
rect 4290 3106 4293 3173
rect 4306 3123 4309 3223
rect 4322 3203 4333 3206
rect 4314 3113 4317 3136
rect 4322 3133 4325 3203
rect 4290 3103 4309 3106
rect 4306 3036 4309 3103
rect 4306 3033 4317 3036
rect 4250 2923 4253 2936
rect 4258 2903 4261 2926
rect 4234 2893 4241 2896
rect 4234 2873 4237 2893
rect 4242 2773 4245 2826
rect 4266 2823 4269 3006
rect 4290 2993 4293 3016
rect 4234 2603 4237 2716
rect 4250 2616 4253 2726
rect 4242 2613 4261 2616
rect 4266 2613 4269 2816
rect 4274 2813 4277 2836
rect 4282 2796 4285 2986
rect 4314 2976 4317 3033
rect 4330 2993 4333 3126
rect 4338 3023 4341 3136
rect 4346 3126 4349 3286
rect 4362 3203 4365 3246
rect 4370 3213 4373 3406
rect 4378 3243 4381 3483
rect 4386 3323 4389 3426
rect 4402 3343 4405 3503
rect 4418 3396 4421 3526
rect 4434 3513 4437 3526
rect 4442 3503 4445 3536
rect 4450 3533 4453 3576
rect 4426 3413 4429 3446
rect 4434 3403 4437 3426
rect 4418 3393 4437 3396
rect 4394 3333 4405 3336
rect 4418 3333 4421 3376
rect 4394 3293 4397 3326
rect 4402 3323 4413 3326
rect 4378 3213 4381 3236
rect 4394 3213 4397 3226
rect 4386 3193 4389 3206
rect 4346 3123 4365 3126
rect 4370 3116 4373 3136
rect 4346 3013 4349 3116
rect 4362 3113 4373 3116
rect 4362 3066 4365 3113
rect 4394 3106 4397 3206
rect 4402 3113 4405 3136
rect 4394 3103 4405 3106
rect 4354 3063 4365 3066
rect 4306 2973 4317 2976
rect 4306 2886 4309 2973
rect 4306 2883 4313 2886
rect 4278 2793 4285 2796
rect 4278 2646 4281 2793
rect 4278 2643 4285 2646
rect 4282 2623 4285 2643
rect 4226 2593 4245 2596
rect 4210 2573 4221 2576
rect 4186 2366 4189 2516
rect 4194 2486 4197 2506
rect 4218 2496 4221 2573
rect 4242 2513 4245 2593
rect 4250 2573 4253 2606
rect 4258 2603 4261 2613
rect 4274 2556 4277 2616
rect 4290 2606 4293 2866
rect 4310 2756 4313 2883
rect 4310 2753 4317 2756
rect 4298 2733 4309 2736
rect 4266 2553 4277 2556
rect 4286 2603 4293 2606
rect 4226 2503 4237 2506
rect 4218 2493 4229 2496
rect 4194 2483 4205 2486
rect 4202 2426 4205 2483
rect 4194 2423 4205 2426
rect 4194 2403 4197 2423
rect 4218 2413 4221 2426
rect 4210 2403 4221 2406
rect 4226 2393 4229 2493
rect 4234 2483 4237 2503
rect 4266 2486 4269 2553
rect 4286 2546 4289 2603
rect 4282 2543 4289 2546
rect 4282 2503 4285 2543
rect 4290 2493 4293 2526
rect 4298 2513 4301 2616
rect 4306 2603 4309 2726
rect 4314 2693 4317 2753
rect 4322 2733 4325 2946
rect 4330 2793 4333 2986
rect 4338 2813 4341 2926
rect 4346 2906 4349 2936
rect 4354 2933 4357 3063
rect 4370 2933 4373 3016
rect 4394 3013 4397 3026
rect 4354 2923 4373 2926
rect 4378 2906 4381 2936
rect 4346 2903 4357 2906
rect 4354 2836 4357 2903
rect 4370 2903 4381 2906
rect 4370 2856 4373 2903
rect 4370 2853 4381 2856
rect 4346 2833 4357 2836
rect 4378 2833 4381 2853
rect 4346 2813 4349 2833
rect 4386 2816 4389 2996
rect 4402 2933 4405 3103
rect 4418 3056 4421 3326
rect 4434 3223 4437 3393
rect 4450 3326 4453 3526
rect 4458 3523 4461 3556
rect 4466 3353 4469 3596
rect 4474 3506 4477 3633
rect 4498 3626 4501 3916
rect 4506 3903 4509 3946
rect 4514 3913 4517 3926
rect 4530 3923 4533 3973
rect 4538 3966 4541 4046
rect 4562 4043 4565 4213
rect 4570 4203 4589 4206
rect 4570 4113 4573 4126
rect 4586 4056 4589 4203
rect 4602 4183 4605 4216
rect 4578 4053 4589 4056
rect 4602 4056 4605 4096
rect 4610 4083 4613 4196
rect 4626 4156 4629 4223
rect 4650 4203 4653 4326
rect 4618 4153 4629 4156
rect 4618 4096 4621 4153
rect 4626 4123 4629 4136
rect 4650 4133 4653 4186
rect 4658 4173 4661 4206
rect 4634 4113 4637 4126
rect 4618 4093 4629 4096
rect 4602 4053 4613 4056
rect 4562 3993 4565 4016
rect 4578 3986 4581 4053
rect 4578 3983 4589 3986
rect 4538 3963 4549 3966
rect 4586 3963 4589 3983
rect 4610 3976 4613 4053
rect 4602 3973 4613 3976
rect 4530 3903 4533 3916
rect 4546 3896 4549 3963
rect 4562 3903 4565 3926
rect 4538 3893 4549 3896
rect 4538 3876 4541 3893
rect 4538 3873 4557 3876
rect 4506 3733 4517 3736
rect 4530 3733 4533 3816
rect 4554 3766 4557 3873
rect 4570 3846 4573 3936
rect 4586 3933 4589 3956
rect 4602 3926 4605 3973
rect 4626 3956 4629 4093
rect 4650 4083 4653 4126
rect 4658 4013 4661 4136
rect 4618 3953 4629 3956
rect 4578 3893 4581 3926
rect 4594 3923 4605 3926
rect 4570 3843 4581 3846
rect 4578 3813 4581 3843
rect 4594 3766 4597 3923
rect 4610 3893 4613 3936
rect 4546 3763 4557 3766
rect 4586 3763 4597 3766
rect 4506 3723 4517 3726
rect 4530 3643 4533 3726
rect 4546 3636 4549 3763
rect 4570 3653 4573 3726
rect 4586 3686 4589 3763
rect 4618 3746 4621 3953
rect 4626 3903 4629 3936
rect 4634 3923 4645 3926
rect 4634 3913 4637 3923
rect 4650 3913 4653 3936
rect 4658 3933 4661 3966
rect 4614 3743 4621 3746
rect 4614 3686 4617 3743
rect 4586 3683 4597 3686
rect 4594 3636 4597 3683
rect 4482 3603 4485 3626
rect 4498 3623 4505 3626
rect 4482 3513 4485 3536
rect 4490 3523 4493 3616
rect 4502 3576 4505 3623
rect 4498 3573 4505 3576
rect 4498 3553 4501 3573
rect 4514 3536 4517 3586
rect 4498 3533 4517 3536
rect 4474 3503 4485 3506
rect 4482 3386 4485 3503
rect 4490 3413 4493 3446
rect 4474 3383 4485 3386
rect 4458 3333 4469 3336
rect 4450 3323 4461 3326
rect 4426 3193 4429 3206
rect 4414 3053 4421 3056
rect 4434 3056 4437 3216
rect 4458 3203 4461 3323
rect 4466 3313 4469 3326
rect 4450 3133 4453 3146
rect 4434 3053 4441 3056
rect 4414 2976 4417 3053
rect 4438 2976 4441 3053
rect 4450 3013 4453 3116
rect 4458 2983 4461 3126
rect 4466 3106 4469 3216
rect 4474 3123 4477 3383
rect 4482 3313 4485 3356
rect 4482 3213 4485 3236
rect 4490 3206 4493 3406
rect 4498 3213 4501 3526
rect 4506 3493 4509 3526
rect 4506 3403 4509 3426
rect 4514 3343 4517 3436
rect 4506 3213 4509 3336
rect 4514 3293 4517 3326
rect 4482 3203 4493 3206
rect 4498 3203 4509 3206
rect 4482 3133 4485 3203
rect 4514 3193 4517 3206
rect 4514 3113 4517 3126
rect 4466 3103 4473 3106
rect 4470 3016 4473 3103
rect 4522 3046 4525 3636
rect 4546 3633 4557 3636
rect 4530 3603 4533 3616
rect 4538 3533 4541 3606
rect 4554 3566 4557 3633
rect 4586 3633 4597 3636
rect 4610 3683 4617 3686
rect 4586 3576 4589 3633
rect 4610 3623 4613 3683
rect 4626 3636 4629 3876
rect 4642 3806 4645 3896
rect 4650 3813 4653 3906
rect 4658 3873 4661 3926
rect 4642 3803 4661 3806
rect 4634 3733 4637 3796
rect 4634 3706 4637 3726
rect 4634 3703 4641 3706
rect 4638 3636 4641 3703
rect 4618 3633 4629 3636
rect 4634 3633 4641 3636
rect 4586 3573 4597 3576
rect 4546 3563 4557 3566
rect 4546 3543 4549 3563
rect 4594 3553 4597 3573
rect 4538 3513 4541 3526
rect 4554 3493 4557 3536
rect 4586 3533 4589 3546
rect 4602 3533 4605 3576
rect 4530 3416 4533 3446
rect 4530 3413 4541 3416
rect 4586 3413 4589 3426
rect 4538 3406 4541 3413
rect 4530 3293 4533 3406
rect 4538 3403 4549 3406
rect 4538 3333 4541 3346
rect 4538 3276 4541 3316
rect 4534 3273 4541 3276
rect 4534 3156 4537 3273
rect 4546 3173 4549 3403
rect 4562 3363 4565 3406
rect 4554 3333 4565 3336
rect 4570 3333 4573 3376
rect 4562 3323 4573 3326
rect 4578 3313 4581 3326
rect 4602 3316 4605 3526
rect 4610 3523 4613 3616
rect 4618 3546 4621 3633
rect 4626 3556 4629 3626
rect 4634 3613 4637 3633
rect 4650 3616 4653 3726
rect 4658 3643 4661 3803
rect 4666 3723 4669 4333
rect 4682 4243 4685 4363
rect 4706 4236 4709 4326
rect 4722 4276 4725 4386
rect 4770 4333 4773 4416
rect 4778 4403 4781 4433
rect 4786 4353 4789 4516
rect 4722 4273 4733 4276
rect 4682 4233 4709 4236
rect 4682 4203 4685 4233
rect 4690 4193 4693 4216
rect 4706 4213 4709 4226
rect 4698 4186 4701 4206
rect 4690 4183 4701 4186
rect 4690 4136 4693 4183
rect 4674 4023 4677 4136
rect 4682 4133 4693 4136
rect 4682 4113 4685 4126
rect 4682 4013 4685 4056
rect 4690 3973 4693 4133
rect 4714 4106 4717 4246
rect 4730 4226 4733 4273
rect 4722 4223 4733 4226
rect 4722 4203 4725 4223
rect 4762 4183 4765 4326
rect 4778 4323 4781 4346
rect 4706 4103 4717 4106
rect 4706 3966 4709 4103
rect 4730 4013 4733 4026
rect 4786 4013 4789 4126
rect 4690 3963 4709 3966
rect 4674 3933 4677 3946
rect 4674 3886 4677 3926
rect 4674 3883 4685 3886
rect 4674 3803 4677 3876
rect 4682 3813 4685 3883
rect 4690 3866 4693 3963
rect 4722 3936 4725 3976
rect 4722 3933 4733 3936
rect 4714 3873 4717 3926
rect 4730 3876 4733 3933
rect 4770 3923 4773 3946
rect 4722 3873 4733 3876
rect 4690 3863 4709 3866
rect 4674 3626 4677 3746
rect 4682 3733 4685 3806
rect 4690 3786 4693 3856
rect 4690 3783 4701 3786
rect 4690 3726 4693 3736
rect 4698 3733 4701 3783
rect 4706 3736 4709 3863
rect 4722 3853 4725 3873
rect 4730 3803 4733 3816
rect 4706 3733 4717 3736
rect 4754 3733 4757 3786
rect 4786 3783 4789 3816
rect 4690 3723 4709 3726
rect 4714 3716 4717 3733
rect 4642 3613 4653 3616
rect 4658 3613 4661 3626
rect 4666 3623 4677 3626
rect 4698 3713 4717 3716
rect 4634 3563 4637 3606
rect 4650 3593 4653 3606
rect 4626 3553 4645 3556
rect 4618 3543 4629 3546
rect 4618 3513 4621 3536
rect 4626 3533 4629 3543
rect 4626 3503 4629 3526
rect 4634 3393 4637 3546
rect 4642 3516 4645 3553
rect 4666 3533 4669 3623
rect 4698 3576 4701 3713
rect 4738 3623 4741 3726
rect 4722 3593 4725 3616
rect 4778 3613 4781 3736
rect 4682 3573 4701 3576
rect 4682 3533 4685 3573
rect 4642 3513 4653 3516
rect 4706 3513 4709 3526
rect 4650 3446 4653 3513
rect 4778 3503 4781 3526
rect 4794 3486 4797 3646
rect 4646 3443 4653 3446
rect 4786 3483 4797 3486
rect 4646 3386 4649 3443
rect 4658 3413 4661 3426
rect 4642 3383 4649 3386
rect 4618 3323 4621 3376
rect 4602 3313 4613 3316
rect 4534 3153 4541 3156
rect 4530 3103 4533 3136
rect 4466 3013 4473 3016
rect 4466 2993 4469 3013
rect 4414 2973 4421 2976
rect 4394 2913 4397 2926
rect 4402 2843 4405 2926
rect 4382 2813 4389 2816
rect 4402 2813 4405 2836
rect 4314 2513 4317 2626
rect 4330 2573 4333 2766
rect 4382 2746 4385 2813
rect 4418 2766 4421 2973
rect 4434 2973 4441 2976
rect 4434 2923 4437 2973
rect 4450 2933 4453 2946
rect 4442 2863 4445 2926
rect 4458 2923 4461 2976
rect 4450 2773 4453 2846
rect 4466 2766 4469 2926
rect 4482 2786 4485 3046
rect 4522 3043 4529 3046
rect 4498 3003 4501 3016
rect 4526 2996 4529 3043
rect 4482 2783 4493 2786
rect 4370 2743 4385 2746
rect 4402 2763 4421 2766
rect 4442 2763 4469 2766
rect 4338 2723 4357 2726
rect 4362 2713 4365 2736
rect 4322 2496 4325 2546
rect 4338 2523 4341 2626
rect 4370 2623 4373 2743
rect 4378 2653 4381 2736
rect 4386 2723 4389 2736
rect 4402 2686 4405 2763
rect 4426 2713 4429 2726
rect 4442 2716 4445 2763
rect 4442 2713 4453 2716
rect 4450 2696 4453 2713
rect 4402 2683 4413 2686
rect 4370 2603 4373 2616
rect 4394 2576 4397 2616
rect 4378 2573 4397 2576
rect 4314 2493 4325 2496
rect 4266 2483 4277 2486
rect 4186 2363 4197 2366
rect 4194 2343 4197 2363
rect 4242 2353 4245 2466
rect 4266 2403 4269 2416
rect 4274 2413 4277 2483
rect 4242 2313 4245 2326
rect 4250 2246 4253 2346
rect 4258 2333 4261 2396
rect 4314 2376 4317 2493
rect 4314 2373 4325 2376
rect 4242 2243 4253 2246
rect 4194 2133 4197 2216
rect 4226 2193 4229 2216
rect 4242 2196 4245 2243
rect 4282 2236 4285 2326
rect 4290 2243 4293 2336
rect 4298 2323 4301 2336
rect 4282 2233 4293 2236
rect 4290 2213 4293 2233
rect 4242 2193 4253 2196
rect 4234 2126 4237 2176
rect 4250 2146 4253 2193
rect 4250 2143 4261 2146
rect 4186 2103 4189 2126
rect 4226 2123 4237 2126
rect 4242 2106 4245 2136
rect 4250 2113 4253 2136
rect 4234 2103 4245 2106
rect 4146 2093 4165 2096
rect 4138 2073 4149 2076
rect 4146 2006 4149 2073
rect 4090 1923 4093 1936
rect 4122 1923 4125 2006
rect 4138 2003 4149 2006
rect 4138 1933 4141 2003
rect 4162 1976 4165 2093
rect 4234 2036 4237 2103
rect 4258 2096 4261 2143
rect 4254 2093 4261 2096
rect 4254 2046 4257 2093
rect 4266 2056 4269 2136
rect 4274 2133 4277 2206
rect 4290 2133 4293 2146
rect 4306 2133 4309 2356
rect 4322 2256 4325 2373
rect 4330 2353 4333 2506
rect 4346 2503 4349 2536
rect 4338 2413 4341 2426
rect 4318 2253 4325 2256
rect 4318 2176 4321 2253
rect 4318 2173 4325 2176
rect 4322 2143 4325 2173
rect 4274 2103 4277 2126
rect 4330 2123 4333 2246
rect 4338 2213 4341 2336
rect 4354 2286 4357 2536
rect 4378 2533 4381 2573
rect 4394 2533 4397 2546
rect 4410 2533 4413 2683
rect 4434 2613 4437 2696
rect 4450 2693 4461 2696
rect 4474 2693 4477 2776
rect 4490 2706 4493 2783
rect 4482 2703 4493 2706
rect 4442 2613 4453 2616
rect 4370 2426 4373 2526
rect 4386 2523 4405 2526
rect 4370 2423 4389 2426
rect 4362 2413 4373 2416
rect 4362 2313 4365 2336
rect 4370 2323 4373 2413
rect 4386 2396 4389 2423
rect 4394 2413 4397 2506
rect 4378 2393 4389 2396
rect 4378 2306 4381 2393
rect 4386 2316 4389 2326
rect 4410 2323 4413 2516
rect 4418 2403 4421 2526
rect 4426 2486 4429 2576
rect 4442 2533 4445 2613
rect 4434 2503 4437 2516
rect 4450 2503 4453 2586
rect 4458 2553 4461 2693
rect 4426 2483 4437 2486
rect 4434 2396 4437 2483
rect 4458 2443 4461 2526
rect 4474 2486 4477 2516
rect 4466 2483 4477 2486
rect 4426 2393 4437 2396
rect 4386 2313 4413 2316
rect 4378 2303 4389 2306
rect 4346 2196 4349 2286
rect 4354 2283 4365 2286
rect 4362 2226 4365 2283
rect 4342 2193 4349 2196
rect 4354 2223 4365 2226
rect 4266 2053 4285 2056
rect 4254 2043 4261 2046
rect 4234 2033 4245 2036
rect 4242 2013 4245 2033
rect 4258 1996 4261 2043
rect 4282 2013 4285 2053
rect 4342 2046 4345 2193
rect 4354 2056 4357 2223
rect 4370 2126 4373 2206
rect 4378 2183 4381 2206
rect 4386 2173 4389 2303
rect 4418 2216 4421 2336
rect 4426 2303 4429 2393
rect 4450 2243 4453 2426
rect 4458 2383 4461 2436
rect 4466 2413 4469 2483
rect 4458 2303 4461 2326
rect 4474 2266 4477 2316
rect 4482 2306 4485 2703
rect 4498 2686 4501 2996
rect 4522 2993 4529 2996
rect 4506 2733 4509 2806
rect 4522 2726 4525 2993
rect 4538 2803 4541 3153
rect 4554 3136 4557 3296
rect 4570 3183 4573 3206
rect 4594 3203 4597 3216
rect 4610 3176 4613 3313
rect 4626 3273 4629 3326
rect 4634 3283 4637 3336
rect 4546 3133 4557 3136
rect 4546 3093 4549 3133
rect 4554 3113 4557 3126
rect 4562 3056 4565 3136
rect 4570 3113 4573 3176
rect 4610 3173 4621 3176
rect 4578 3123 4581 3156
rect 4586 3123 4589 3146
rect 4546 3053 4565 3056
rect 4546 3013 4549 3053
rect 4570 2946 4573 3096
rect 4578 3013 4581 3106
rect 4602 3016 4605 3116
rect 4618 3043 4621 3173
rect 4634 3166 4637 3246
rect 4630 3163 4637 3166
rect 4630 3036 4633 3163
rect 4630 3033 4637 3036
rect 4594 3013 4605 3016
rect 4594 2956 4597 3013
rect 4594 2953 4605 2956
rect 4554 2943 4573 2946
rect 4554 2883 4557 2943
rect 4562 2876 4565 2936
rect 4570 2933 4573 2943
rect 4570 2923 4589 2926
rect 4562 2873 4573 2876
rect 4494 2683 4501 2686
rect 4506 2723 4525 2726
rect 4494 2386 4497 2683
rect 4506 2423 4509 2723
rect 4506 2393 4509 2406
rect 4494 2383 4501 2386
rect 4498 2306 4501 2383
rect 4514 2373 4517 2696
rect 4522 2603 4525 2636
rect 4530 2616 4533 2736
rect 4538 2703 4541 2726
rect 4554 2723 4557 2866
rect 4570 2813 4573 2873
rect 4570 2693 4573 2726
rect 4578 2713 4581 2736
rect 4546 2616 4549 2626
rect 4530 2613 4549 2616
rect 4538 2573 4541 2606
rect 4522 2436 4525 2536
rect 4530 2493 4533 2526
rect 4546 2446 4549 2536
rect 4554 2533 4557 2596
rect 4562 2533 4565 2606
rect 4586 2603 4589 2886
rect 4594 2856 4597 2936
rect 4602 2923 4605 2953
rect 4610 2913 4613 3006
rect 4626 2936 4629 3016
rect 4634 2986 4637 3033
rect 4642 3003 4645 3383
rect 4650 3316 4653 3346
rect 4658 3333 4661 3396
rect 4674 3373 4677 3416
rect 4650 3313 4657 3316
rect 4654 3246 4657 3313
rect 4650 3243 4657 3246
rect 4650 3206 4653 3243
rect 4658 3213 4661 3226
rect 4650 3203 4661 3206
rect 4658 3163 4661 3203
rect 4650 3083 4653 3136
rect 4658 3133 4661 3156
rect 4658 3113 4661 3126
rect 4666 3036 4669 3256
rect 4674 3243 4677 3366
rect 4698 3323 4701 3336
rect 4754 3323 4757 3406
rect 4786 3356 4789 3483
rect 4786 3353 4797 3356
rect 4794 3336 4797 3353
rect 4682 3213 4685 3286
rect 4762 3283 4765 3326
rect 4786 3266 4789 3336
rect 4794 3333 4801 3336
rect 4778 3263 4789 3266
rect 4674 3143 4677 3206
rect 4650 3033 4669 3036
rect 4650 3013 4653 3033
rect 4674 3023 4677 3136
rect 4682 3113 4685 3126
rect 4658 2986 4661 3006
rect 4634 2983 4645 2986
rect 4626 2933 4633 2936
rect 4594 2853 4613 2856
rect 4610 2813 4613 2853
rect 4610 2633 4613 2806
rect 4618 2723 4621 2926
rect 4630 2886 4633 2933
rect 4626 2883 4633 2886
rect 4626 2723 4629 2883
rect 4642 2866 4645 2983
rect 4654 2983 4661 2986
rect 4654 2916 4657 2983
rect 4666 2923 4669 3016
rect 4654 2913 4661 2916
rect 4634 2863 4645 2866
rect 4634 2813 4637 2863
rect 4658 2823 4661 2913
rect 4658 2756 4661 2816
rect 4682 2793 4685 2996
rect 4690 2966 4693 3206
rect 4698 3203 4701 3226
rect 4706 3213 4709 3236
rect 4706 2993 4709 3186
rect 4778 3176 4781 3263
rect 4798 3256 4801 3333
rect 4794 3253 4801 3256
rect 4794 3186 4797 3253
rect 4794 3183 4801 3186
rect 4778 3173 4789 3176
rect 4730 3123 4733 3146
rect 4786 3123 4789 3173
rect 4730 3013 4733 3026
rect 4786 3013 4789 3086
rect 4798 3016 4801 3183
rect 4794 3013 4801 3016
rect 4794 2996 4797 3013
rect 4786 2993 4797 2996
rect 4690 2963 4717 2966
rect 4706 2813 4709 2826
rect 4658 2753 4677 2756
rect 4658 2733 4661 2746
rect 4650 2706 4653 2726
rect 4666 2713 4669 2726
rect 4674 2706 4677 2753
rect 4642 2703 4653 2706
rect 4666 2703 4677 2706
rect 4602 2603 4605 2616
rect 4562 2513 4565 2526
rect 4546 2443 4557 2446
rect 4522 2433 4541 2436
rect 4514 2323 4517 2336
rect 4522 2323 4525 2416
rect 4530 2403 4533 2426
rect 4538 2413 4541 2433
rect 4554 2396 4557 2443
rect 4570 2413 4573 2536
rect 4578 2476 4581 2506
rect 4586 2493 4589 2536
rect 4610 2523 4613 2576
rect 4578 2473 4589 2476
rect 4586 2426 4589 2473
rect 4618 2456 4621 2656
rect 4642 2636 4645 2703
rect 4642 2633 4653 2636
rect 4578 2423 4589 2426
rect 4602 2453 4621 2456
rect 4546 2393 4557 2396
rect 4546 2366 4549 2393
rect 4530 2363 4549 2366
rect 4530 2326 4533 2363
rect 4538 2333 4541 2346
rect 4546 2333 4549 2356
rect 4530 2323 4549 2326
rect 4482 2303 4489 2306
rect 4498 2303 4509 2306
rect 4466 2263 4477 2266
rect 4402 2213 4421 2216
rect 4394 2133 4397 2206
rect 4410 2143 4413 2206
rect 4442 2136 4445 2206
rect 4434 2133 4445 2136
rect 4370 2123 4389 2126
rect 4434 2123 4437 2133
rect 4354 2053 4361 2056
rect 4342 2043 4349 2046
rect 4330 2003 4333 2026
rect 4346 2023 4349 2043
rect 4258 1993 4269 1996
rect 4146 1973 4165 1976
rect 4146 1953 4149 1973
rect 4210 1933 4213 1946
rect 3962 1823 3973 1826
rect 3530 1643 3533 1726
rect 3546 1713 3549 1736
rect 3594 1723 3597 1746
rect 3666 1716 3669 1736
rect 3698 1733 3701 1746
rect 3466 1593 3469 1606
rect 3450 1553 3461 1556
rect 3450 1503 3453 1553
rect 3458 1533 3461 1546
rect 3466 1523 3469 1546
rect 3554 1543 3557 1616
rect 3562 1573 3565 1626
rect 3570 1613 3573 1636
rect 3578 1613 3581 1646
rect 3570 1543 3573 1606
rect 3578 1533 3581 1556
rect 3442 1483 3453 1486
rect 3450 1366 3453 1483
rect 3442 1363 3453 1366
rect 3442 1343 3445 1363
rect 3498 1333 3501 1346
rect 3514 1333 3517 1356
rect 3386 1293 3393 1296
rect 3386 1273 3389 1293
rect 3346 1213 3349 1226
rect 3338 1203 3349 1206
rect 3354 1203 3357 1236
rect 3410 1233 3413 1326
rect 3506 1323 3517 1326
rect 3522 1316 3525 1506
rect 3538 1413 3541 1426
rect 3514 1313 3525 1316
rect 3514 1256 3517 1313
rect 3514 1253 3521 1256
rect 3306 1113 3309 1126
rect 3330 1096 3333 1146
rect 3290 1093 3301 1096
rect 3298 1026 3301 1093
rect 3266 1013 3277 1016
rect 3282 1013 3285 1026
rect 3290 1023 3301 1026
rect 3322 1093 3333 1096
rect 3266 916 3269 1013
rect 3290 966 3293 1023
rect 3298 993 3301 1006
rect 3290 963 3301 966
rect 3274 923 3277 946
rect 3298 933 3301 963
rect 3322 956 3325 1093
rect 3338 1026 3341 1186
rect 3346 1143 3349 1203
rect 3362 1193 3365 1206
rect 3362 1136 3365 1176
rect 3362 1133 3373 1136
rect 3394 1133 3397 1146
rect 3354 1043 3357 1126
rect 3370 1106 3373 1133
rect 3402 1126 3405 1146
rect 3450 1143 3453 1216
rect 3458 1213 3461 1226
rect 3466 1193 3469 1206
rect 3482 1203 3485 1216
rect 3518 1176 3521 1253
rect 3514 1173 3521 1176
rect 3498 1133 3509 1136
rect 3386 1123 3405 1126
rect 3370 1103 3381 1106
rect 3378 1036 3381 1103
rect 3370 1033 3381 1036
rect 3490 1036 3493 1126
rect 3498 1113 3501 1126
rect 3514 1116 3517 1173
rect 3510 1113 3517 1116
rect 3510 1056 3513 1113
rect 3510 1053 3517 1056
rect 3490 1033 3509 1036
rect 3338 1023 3349 1026
rect 3346 956 3349 1023
rect 3322 953 3333 956
rect 3266 913 3277 916
rect 3250 666 3253 756
rect 3258 733 3261 776
rect 3274 736 3277 913
rect 3290 793 3293 926
rect 3274 733 3281 736
rect 3250 663 3261 666
rect 3226 583 3229 606
rect 3250 593 3253 616
rect 3258 586 3261 663
rect 3266 633 3269 726
rect 3278 666 3281 733
rect 3290 706 3293 786
rect 3298 723 3301 816
rect 3306 803 3309 936
rect 3314 883 3317 926
rect 3314 733 3317 826
rect 3322 813 3325 926
rect 3330 893 3333 953
rect 3338 953 3349 956
rect 3338 933 3341 953
rect 3346 906 3349 926
rect 3354 913 3357 936
rect 3342 903 3349 906
rect 3362 903 3365 926
rect 3370 923 3373 1033
rect 3394 963 3397 1006
rect 3402 1003 3405 1016
rect 3342 836 3345 903
rect 3342 833 3349 836
rect 3330 793 3333 806
rect 3338 763 3341 816
rect 3346 773 3349 833
rect 3354 786 3357 896
rect 3362 796 3365 816
rect 3370 803 3373 896
rect 3410 893 3413 1016
rect 3506 1003 3509 1033
rect 3458 923 3461 936
rect 3474 933 3477 996
rect 3482 933 3485 946
rect 3466 913 3469 926
rect 3362 793 3381 796
rect 3354 783 3373 786
rect 3370 736 3373 783
rect 3290 703 3301 706
rect 3274 663 3281 666
rect 3242 583 3261 586
rect 3242 556 3245 583
rect 3266 566 3269 626
rect 3226 553 3245 556
rect 3226 543 3229 553
rect 3186 526 3189 536
rect 3150 523 3157 526
rect 3170 523 3189 526
rect 3154 506 3157 523
rect 3154 503 3165 506
rect 3162 436 3165 503
rect 3154 433 3165 436
rect 3114 273 3133 276
rect 3130 213 3133 273
rect 3154 233 3157 433
rect 3234 413 3237 546
rect 3242 533 3245 553
rect 3262 563 3269 566
rect 3242 503 3245 526
rect 3250 513 3253 536
rect 3262 476 3265 563
rect 3274 503 3277 663
rect 3298 646 3301 703
rect 3330 686 3333 734
rect 3362 733 3373 736
rect 3418 733 3421 766
rect 3330 683 3349 686
rect 3290 643 3301 646
rect 3290 623 3293 643
rect 3330 593 3333 616
rect 3262 473 3269 476
rect 3266 456 3269 473
rect 3266 453 3277 456
rect 3106 193 3109 206
rect 3170 193 3173 366
rect 3202 363 3205 406
rect 3274 396 3277 453
rect 3266 393 3277 396
rect 3266 376 3269 393
rect 3250 373 3269 376
rect 3194 323 3197 356
rect 3250 306 3253 373
rect 3282 333 3285 366
rect 3298 363 3301 586
rect 3346 583 3349 683
rect 3362 666 3365 733
rect 3378 676 3381 726
rect 3378 673 3389 676
rect 3410 673 3413 726
rect 3426 723 3429 736
rect 3466 733 3469 816
rect 3474 813 3477 886
rect 3482 783 3485 836
rect 3490 793 3493 956
rect 3498 933 3501 996
rect 3514 936 3517 1053
rect 3522 1013 3525 1136
rect 3530 993 3533 1346
rect 3546 1323 3549 1506
rect 3554 1353 3557 1526
rect 3562 1423 3565 1526
rect 3594 1506 3597 1716
rect 3658 1713 3669 1716
rect 3602 1613 3613 1616
rect 3618 1613 3621 1646
rect 3658 1626 3661 1713
rect 3658 1623 3669 1626
rect 3610 1593 3613 1606
rect 3626 1523 3629 1606
rect 3634 1566 3637 1616
rect 3642 1583 3645 1606
rect 3666 1583 3669 1623
rect 3634 1563 3641 1566
rect 3638 1516 3641 1563
rect 3674 1523 3677 1606
rect 3682 1523 3685 1726
rect 3690 1713 3693 1726
rect 3706 1703 3709 1726
rect 3714 1723 3717 1736
rect 3762 1733 3765 1816
rect 3802 1776 3805 1816
rect 3794 1773 3805 1776
rect 3714 1616 3717 1626
rect 3706 1613 3717 1616
rect 3722 1613 3733 1616
rect 3738 1606 3741 1726
rect 3746 1613 3749 1626
rect 3706 1593 3709 1606
rect 3578 1503 3597 1506
rect 3634 1513 3641 1516
rect 3562 1403 3565 1416
rect 3578 1403 3581 1503
rect 3634 1456 3637 1513
rect 3618 1453 3637 1456
rect 3602 1376 3605 1416
rect 3586 1373 3605 1376
rect 3586 1333 3589 1373
rect 3594 1333 3605 1336
rect 3538 1213 3541 1226
rect 3538 1133 3541 1206
rect 3562 1203 3565 1326
rect 3570 1243 3573 1326
rect 3538 1093 3541 1126
rect 3554 1026 3557 1156
rect 3578 1133 3581 1326
rect 3594 1303 3597 1326
rect 3610 1313 3613 1326
rect 3618 1296 3621 1453
rect 3690 1436 3693 1586
rect 3722 1533 3725 1606
rect 3738 1603 3749 1606
rect 3754 1603 3757 1716
rect 3778 1696 3781 1756
rect 3794 1733 3797 1773
rect 3810 1766 3813 1806
rect 3850 1793 3853 1806
rect 3882 1793 3885 1806
rect 3802 1763 3813 1766
rect 3770 1693 3781 1696
rect 3770 1596 3773 1693
rect 3786 1626 3789 1706
rect 3802 1643 3805 1763
rect 3826 1733 3829 1746
rect 3834 1733 3837 1756
rect 3842 1706 3845 1726
rect 3850 1713 3853 1736
rect 3834 1703 3845 1706
rect 3762 1593 3773 1596
rect 3782 1623 3789 1626
rect 3674 1433 3693 1436
rect 3658 1333 3661 1416
rect 3674 1333 3677 1433
rect 3690 1403 3693 1416
rect 3714 1333 3717 1526
rect 3722 1503 3725 1526
rect 3746 1513 3749 1536
rect 3722 1333 3725 1416
rect 3730 1333 3741 1336
rect 3594 1293 3621 1296
rect 3586 1153 3589 1246
rect 3586 1113 3589 1126
rect 3594 1096 3597 1293
rect 3602 1183 3605 1206
rect 3610 1196 3613 1216
rect 3618 1203 3621 1226
rect 3626 1196 3629 1306
rect 3706 1293 3709 1326
rect 3714 1246 3717 1326
rect 3730 1303 3733 1326
rect 3746 1313 3749 1326
rect 3714 1243 3725 1246
rect 3674 1203 3677 1216
rect 3690 1203 3693 1226
rect 3722 1196 3725 1243
rect 3738 1203 3741 1216
rect 3610 1193 3621 1196
rect 3626 1193 3645 1196
rect 3586 1093 3597 1096
rect 3586 1036 3589 1093
rect 3586 1033 3597 1036
rect 3554 1023 3565 1026
rect 3538 953 3541 1016
rect 3546 993 3549 1006
rect 3562 956 3565 1023
rect 3594 1013 3597 1033
rect 3602 1006 3605 1136
rect 3610 1093 3613 1126
rect 3618 1113 3621 1193
rect 3626 1166 3629 1186
rect 3626 1163 3633 1166
rect 3630 1106 3633 1163
rect 3626 1103 3633 1106
rect 3554 953 3565 956
rect 3594 1003 3605 1006
rect 3554 936 3557 953
rect 3506 933 3525 936
rect 3546 933 3557 936
rect 3578 933 3589 936
rect 3522 923 3533 926
rect 3522 886 3525 923
rect 3522 883 3533 886
rect 3482 733 3485 746
rect 3506 733 3509 876
rect 3530 836 3533 883
rect 3522 833 3533 836
rect 3522 816 3525 833
rect 3546 816 3549 933
rect 3562 823 3565 916
rect 3570 903 3573 926
rect 3594 923 3597 1003
rect 3602 913 3605 936
rect 3610 913 3613 936
rect 3618 923 3621 1006
rect 3626 916 3629 1103
rect 3642 1026 3645 1193
rect 3714 1193 3725 1196
rect 3666 1133 3669 1146
rect 3682 1093 3685 1126
rect 3634 1023 3645 1026
rect 3634 926 3637 1023
rect 3666 1013 3669 1026
rect 3682 1013 3685 1086
rect 3658 993 3661 1006
rect 3642 933 3645 986
rect 3674 946 3677 1006
rect 3690 953 3693 1136
rect 3698 1123 3701 1146
rect 3706 1113 3709 1136
rect 3666 943 3677 946
rect 3650 933 3661 936
rect 3634 923 3645 926
rect 3666 923 3669 943
rect 3622 913 3629 916
rect 3522 813 3533 816
rect 3546 813 3557 816
rect 3514 733 3517 746
rect 3554 733 3557 813
rect 3562 733 3565 746
rect 3586 733 3589 866
rect 3602 813 3605 846
rect 3610 803 3613 906
rect 3622 826 3625 913
rect 3634 853 3637 916
rect 3642 846 3645 923
rect 3618 823 3625 826
rect 3634 843 3645 846
rect 3474 686 3477 726
rect 3474 683 3485 686
rect 3362 663 3373 666
rect 3322 523 3325 536
rect 3314 413 3317 426
rect 3362 413 3365 506
rect 3338 363 3341 406
rect 3370 386 3373 663
rect 3386 466 3389 673
rect 3466 613 3469 676
rect 3482 636 3485 683
rect 3474 633 3485 636
rect 3474 613 3477 633
rect 3450 603 3469 606
rect 3474 603 3493 606
rect 3458 533 3461 596
rect 3498 533 3501 616
rect 3506 613 3509 636
rect 3514 613 3517 726
rect 3522 703 3525 716
rect 3554 703 3557 716
rect 3458 493 3461 526
rect 3466 513 3485 516
rect 3506 513 3509 526
rect 3362 383 3373 386
rect 3378 463 3389 466
rect 3266 313 3269 326
rect 3306 323 3309 346
rect 3250 303 3261 306
rect 3258 256 3261 303
rect 3362 276 3365 383
rect 3250 253 3261 256
rect 3354 273 3365 276
rect 3194 213 3197 226
rect 3234 213 3237 236
rect 3210 193 3213 206
rect 2986 113 2989 126
rect 3002 123 3005 146
rect 3082 123 3085 136
rect 3130 133 3133 176
rect 3250 146 3253 253
rect 3250 143 3261 146
rect 3146 103 3149 126
rect 3258 113 3261 143
rect 3282 133 3285 196
rect 3306 193 3309 216
rect 3314 183 3317 216
rect 3354 206 3357 273
rect 3378 266 3381 463
rect 3426 403 3429 426
rect 3434 393 3437 416
rect 3458 413 3461 456
rect 3466 426 3469 513
rect 3466 423 3493 426
rect 3466 393 3469 406
rect 3474 386 3477 423
rect 3506 403 3509 416
rect 3514 403 3517 536
rect 3522 413 3525 626
rect 3530 593 3533 606
rect 3546 596 3549 636
rect 3554 603 3557 616
rect 3562 613 3565 626
rect 3546 593 3557 596
rect 3466 383 3477 386
rect 3418 336 3421 356
rect 3410 333 3421 336
rect 3410 323 3421 326
rect 3418 303 3421 316
rect 3442 313 3445 336
rect 3370 263 3381 266
rect 3370 213 3373 263
rect 3354 203 3365 206
rect 3298 123 3301 166
rect 3362 123 3365 203
rect 3394 176 3397 206
rect 3410 203 3413 226
rect 3466 223 3469 383
rect 3506 343 3509 356
rect 3482 313 3485 326
rect 3498 323 3501 336
rect 3506 326 3509 336
rect 3530 333 3533 426
rect 3538 413 3541 526
rect 3554 423 3557 593
rect 3570 436 3573 726
rect 3578 623 3581 636
rect 3586 613 3589 626
rect 3594 603 3597 736
rect 3618 733 3621 823
rect 3610 713 3621 716
rect 3610 703 3613 713
rect 3626 706 3629 806
rect 3634 713 3637 843
rect 3642 723 3645 826
rect 3658 766 3661 846
rect 3666 803 3669 916
rect 3682 913 3685 936
rect 3674 813 3677 826
rect 3650 763 3661 766
rect 3650 723 3653 763
rect 3658 733 3661 746
rect 3674 733 3677 806
rect 3690 803 3693 936
rect 3698 923 3701 1106
rect 3706 1013 3709 1096
rect 3714 993 3717 1193
rect 3722 916 3725 1166
rect 3730 1106 3733 1126
rect 3730 1103 3741 1106
rect 3738 1036 3741 1103
rect 3730 1033 3741 1036
rect 3730 1003 3733 1033
rect 3738 993 3741 1006
rect 3754 956 3757 1536
rect 3762 1183 3765 1593
rect 3782 1536 3785 1623
rect 3794 1613 3805 1616
rect 3774 1533 3785 1536
rect 3774 1436 3777 1533
rect 3770 1433 3777 1436
rect 3770 1316 3773 1433
rect 3778 1333 3781 1416
rect 3786 1413 3789 1526
rect 3794 1523 3797 1606
rect 3810 1603 3813 1656
rect 3834 1626 3837 1703
rect 3858 1646 3861 1726
rect 3850 1643 3861 1646
rect 3834 1623 3845 1626
rect 3818 1593 3821 1606
rect 3810 1423 3813 1526
rect 3834 1516 3837 1536
rect 3826 1513 3837 1516
rect 3826 1446 3829 1513
rect 3826 1443 3837 1446
rect 3818 1413 3821 1426
rect 3834 1423 3837 1443
rect 3770 1313 3777 1316
rect 3774 1236 3777 1313
rect 3770 1233 3777 1236
rect 3714 913 3725 916
rect 3746 953 3757 956
rect 3714 816 3717 913
rect 3746 893 3749 953
rect 3754 933 3757 946
rect 3762 916 3765 956
rect 3758 913 3765 916
rect 3758 836 3761 913
rect 3758 833 3765 836
rect 3714 813 3721 816
rect 3682 733 3693 736
rect 3618 703 3629 706
rect 3578 533 3581 556
rect 3586 533 3589 546
rect 3594 503 3597 516
rect 3570 433 3581 436
rect 3554 333 3557 416
rect 3506 323 3525 326
rect 3562 323 3565 416
rect 3570 413 3573 426
rect 3474 213 3477 236
rect 3482 223 3501 226
rect 3466 193 3469 206
rect 3490 203 3493 216
rect 3386 173 3397 176
rect 3386 133 3389 173
rect 3418 133 3421 146
rect 3442 113 3445 126
rect 3498 123 3501 216
rect 3506 213 3509 246
rect 3522 213 3525 323
rect 3530 213 3533 246
rect 3570 236 3573 406
rect 3578 346 3581 433
rect 3602 413 3605 526
rect 3594 393 3597 406
rect 3578 343 3589 346
rect 3594 343 3597 376
rect 3586 323 3589 343
rect 3586 293 3589 316
rect 3570 233 3581 236
rect 3522 133 3525 206
rect 3570 203 3573 216
rect 3578 203 3581 233
rect 3594 213 3597 336
rect 3610 333 3613 606
rect 3618 466 3621 703
rect 3642 616 3645 716
rect 3650 696 3653 716
rect 3666 703 3669 726
rect 3674 723 3685 726
rect 3698 706 3701 746
rect 3690 703 3701 706
rect 3650 693 3657 696
rect 3634 613 3645 616
rect 3634 536 3637 613
rect 3654 606 3657 693
rect 3690 636 3693 703
rect 3690 633 3701 636
rect 3650 603 3657 606
rect 3650 536 3653 603
rect 3626 533 3637 536
rect 3646 533 3653 536
rect 3626 486 3629 533
rect 3626 483 3637 486
rect 3618 463 3625 466
rect 3622 376 3625 463
rect 3618 373 3625 376
rect 3618 316 3621 373
rect 3634 356 3637 483
rect 3646 436 3649 533
rect 3646 433 3653 436
rect 3650 413 3653 433
rect 3658 393 3661 526
rect 3666 523 3669 616
rect 3698 613 3701 633
rect 3706 606 3709 806
rect 3718 756 3721 813
rect 3698 603 3709 606
rect 3714 753 3721 756
rect 3714 603 3717 753
rect 3674 533 3677 546
rect 3682 443 3685 536
rect 3666 413 3669 426
rect 3674 413 3685 416
rect 3698 413 3701 603
rect 3610 313 3621 316
rect 3626 353 3637 356
rect 3626 313 3629 353
rect 3674 346 3677 406
rect 3682 356 3685 413
rect 3682 353 3693 356
rect 3610 236 3613 313
rect 3634 306 3637 336
rect 3626 303 3637 306
rect 3610 233 3621 236
rect 3618 213 3621 233
rect 3570 123 3573 146
rect 3602 93 3605 206
rect 3626 193 3629 303
rect 3642 293 3645 316
rect 3626 123 3629 176
rect 3642 143 3645 206
rect 3650 163 3653 226
rect 3658 213 3661 346
rect 3674 343 3685 346
rect 3682 323 3685 343
rect 3674 203 3677 216
rect 3682 213 3685 316
rect 3690 296 3693 353
rect 3706 313 3709 446
rect 3714 403 3717 536
rect 3722 366 3725 736
rect 3730 683 3733 816
rect 3738 793 3741 806
rect 3746 803 3749 816
rect 3762 813 3765 833
rect 3738 733 3741 786
rect 3754 773 3757 806
rect 3746 733 3757 736
rect 3746 673 3749 726
rect 3730 523 3733 606
rect 3746 566 3749 666
rect 3754 616 3757 726
rect 3762 703 3765 726
rect 3770 663 3773 1233
rect 3778 1133 3781 1216
rect 3778 783 3781 936
rect 3786 903 3789 1406
rect 3794 1233 3797 1326
rect 3818 1313 3821 1406
rect 3842 1316 3845 1623
rect 3850 1613 3853 1643
rect 3866 1613 3869 1636
rect 3874 1616 3877 1736
rect 3890 1726 3893 1736
rect 3898 1733 3901 1786
rect 3914 1733 3917 1816
rect 3930 1733 3933 1746
rect 3882 1633 3885 1726
rect 3890 1723 3901 1726
rect 3898 1653 3901 1723
rect 3922 1703 3925 1726
rect 3938 1713 3941 1726
rect 3922 1633 3941 1636
rect 3874 1613 3885 1616
rect 3858 1413 3861 1606
rect 3866 1603 3877 1606
rect 3874 1403 3877 1536
rect 3882 1523 3885 1613
rect 3898 1553 3901 1616
rect 3906 1576 3909 1626
rect 3922 1613 3925 1633
rect 3906 1573 3917 1576
rect 3882 1386 3885 1406
rect 3866 1383 3885 1386
rect 3842 1313 3853 1316
rect 3794 1133 3797 1206
rect 3802 1123 3805 1216
rect 3818 1203 3829 1206
rect 3834 1166 3837 1306
rect 3850 1236 3853 1313
rect 3842 1233 3853 1236
rect 3866 1236 3869 1383
rect 3890 1246 3893 1536
rect 3914 1533 3917 1573
rect 3930 1563 3933 1606
rect 3938 1603 3941 1626
rect 3922 1516 3925 1536
rect 3906 1386 3909 1406
rect 3902 1383 3909 1386
rect 3902 1266 3905 1383
rect 3902 1263 3909 1266
rect 3890 1243 3897 1246
rect 3866 1233 3885 1236
rect 3842 1183 3845 1233
rect 3850 1193 3853 1216
rect 3866 1203 3869 1216
rect 3882 1186 3885 1233
rect 3874 1183 3885 1186
rect 3834 1163 3853 1166
rect 3794 1013 3797 1036
rect 3810 1013 3813 1146
rect 3802 936 3805 1006
rect 3818 1003 3821 1016
rect 3826 1013 3829 1136
rect 3850 1056 3853 1163
rect 3834 1053 3853 1056
rect 3834 1036 3837 1053
rect 3834 1033 3845 1036
rect 3794 933 3805 936
rect 3794 923 3797 933
rect 3810 923 3813 966
rect 3834 933 3837 1026
rect 3842 1016 3845 1033
rect 3842 1013 3849 1016
rect 3846 936 3849 1013
rect 3874 996 3877 1183
rect 3894 1176 3897 1243
rect 3906 1223 3909 1263
rect 3914 1206 3917 1516
rect 3922 1513 3933 1516
rect 3930 1446 3933 1513
rect 3922 1443 3933 1446
rect 3922 1376 3925 1443
rect 3946 1403 3949 1796
rect 3962 1726 3965 1823
rect 3978 1733 3981 1816
rect 3962 1723 3973 1726
rect 3954 1613 3965 1616
rect 3954 1523 3957 1606
rect 3970 1493 3973 1723
rect 3978 1613 3981 1626
rect 3994 1593 3997 1816
rect 4018 1803 4021 1816
rect 4026 1783 4029 1806
rect 4042 1803 4045 1906
rect 4002 1733 4005 1756
rect 4018 1733 4021 1756
rect 4002 1583 4005 1606
rect 4018 1603 4021 1716
rect 4042 1713 4045 1726
rect 4050 1636 4053 1816
rect 4130 1813 4133 1926
rect 4058 1743 4061 1806
rect 4154 1756 4157 1816
rect 4162 1803 4165 1916
rect 4170 1903 4173 1926
rect 4226 1826 4229 1926
rect 4242 1836 4245 1926
rect 4258 1913 4261 1926
rect 4266 1836 4269 1993
rect 4242 1833 4249 1836
rect 4226 1823 4237 1826
rect 4178 1783 4181 1806
rect 4210 1766 4213 1816
rect 4234 1803 4237 1823
rect 4246 1776 4249 1833
rect 4258 1833 4269 1836
rect 4258 1786 4261 1833
rect 4258 1783 4277 1786
rect 4282 1783 4285 1946
rect 4306 1933 4309 1946
rect 4346 1933 4349 2016
rect 4358 1976 4361 2053
rect 4354 1973 4361 1976
rect 4338 1913 4341 1926
rect 4354 1916 4357 1973
rect 4362 1933 4365 1956
rect 4378 1933 4381 2016
rect 4426 1973 4429 2006
rect 4394 1933 4397 1966
rect 4442 1956 4445 2016
rect 4450 2006 4453 2226
rect 4458 2213 4461 2236
rect 4466 2213 4469 2263
rect 4466 2123 4469 2136
rect 4474 2016 4477 2246
rect 4486 2236 4489 2303
rect 4506 2246 4509 2303
rect 4482 2233 4489 2236
rect 4498 2243 4509 2246
rect 4482 2213 4485 2233
rect 4498 2223 4501 2243
rect 4530 2213 4533 2306
rect 4522 2193 4525 2206
rect 4538 2203 4541 2226
rect 4546 2213 4549 2323
rect 4554 2306 4557 2376
rect 4578 2336 4581 2423
rect 4602 2393 4605 2453
rect 4618 2413 4621 2426
rect 4562 2333 4573 2336
rect 4578 2333 4597 2336
rect 4562 2323 4589 2326
rect 4554 2303 4565 2306
rect 4562 2236 4565 2303
rect 4554 2233 4565 2236
rect 4546 2183 4549 2206
rect 4554 2203 4557 2233
rect 4570 2143 4573 2206
rect 4578 2193 4581 2216
rect 4594 2163 4597 2333
rect 4602 2323 4605 2386
rect 4626 2363 4629 2616
rect 4634 2383 4637 2616
rect 4650 2613 4653 2633
rect 4666 2596 4669 2703
rect 4658 2593 4669 2596
rect 4658 2526 4661 2593
rect 4674 2533 4677 2606
rect 4682 2593 4685 2616
rect 4690 2603 4693 2776
rect 4698 2613 4701 2626
rect 4706 2606 4709 2796
rect 4714 2773 4717 2963
rect 4762 2813 4765 2936
rect 4786 2836 4789 2993
rect 4786 2833 4797 2836
rect 4794 2816 4797 2833
rect 4730 2723 4733 2746
rect 4770 2713 4773 2816
rect 4794 2813 4801 2816
rect 4786 2723 4789 2806
rect 4798 2716 4801 2813
rect 4794 2713 4801 2716
rect 4794 2696 4797 2713
rect 4786 2693 4797 2696
rect 4786 2626 4789 2693
rect 4786 2623 4793 2626
rect 4698 2603 4709 2606
rect 4658 2523 4669 2526
rect 4682 2523 4685 2546
rect 4618 2323 4621 2336
rect 4626 2333 4629 2356
rect 4642 2333 4645 2406
rect 4666 2393 4669 2523
rect 4698 2376 4701 2603
rect 4714 2543 4717 2606
rect 4722 2593 4725 2616
rect 4722 2523 4725 2536
rect 4778 2523 4781 2606
rect 4790 2506 4793 2623
rect 4786 2503 4793 2506
rect 4786 2436 4789 2503
rect 4786 2433 4793 2436
rect 4722 2403 4725 2416
rect 4698 2373 4717 2376
rect 4650 2326 4653 2346
rect 4658 2333 4661 2366
rect 4514 2023 4517 2136
rect 4570 2123 4573 2136
rect 4594 2123 4597 2146
rect 4602 2123 4605 2216
rect 4618 2183 4621 2316
rect 4634 2213 4637 2326
rect 4650 2323 4669 2326
rect 4674 2316 4677 2336
rect 4658 2313 4677 2316
rect 4650 2213 4653 2226
rect 4642 2133 4645 2206
rect 4658 2203 4661 2313
rect 4674 2203 4677 2216
rect 4698 2213 4701 2336
rect 4714 2266 4717 2373
rect 4706 2263 4717 2266
rect 4706 2206 4709 2263
rect 4738 2213 4741 2396
rect 4778 2333 4781 2416
rect 4790 2336 4793 2433
rect 4790 2333 4797 2336
rect 4754 2306 4757 2326
rect 4794 2313 4797 2333
rect 4754 2303 4765 2306
rect 4762 2246 4765 2303
rect 4802 2296 4805 2606
rect 4754 2243 4765 2246
rect 4794 2293 4805 2296
rect 4754 2213 4757 2243
rect 4762 2213 4765 2226
rect 4698 2203 4709 2206
rect 4674 2123 4677 2196
rect 4698 2133 4701 2203
rect 4722 2123 4725 2136
rect 4778 2123 4781 2206
rect 4794 2036 4797 2293
rect 4794 2033 4801 2036
rect 4458 2013 4477 2016
rect 4450 2003 4469 2006
rect 4442 1953 4449 1956
rect 4434 1933 4437 1946
rect 4350 1913 4357 1916
rect 4350 1846 4353 1913
rect 4350 1843 4357 1846
rect 4354 1823 4357 1843
rect 4202 1763 4213 1766
rect 4242 1773 4249 1776
rect 4146 1753 4157 1756
rect 4098 1733 4117 1736
rect 4098 1723 4101 1733
rect 4026 1633 4053 1636
rect 4026 1596 4029 1633
rect 4010 1593 4029 1596
rect 4010 1536 4013 1593
rect 4034 1586 4037 1616
rect 4058 1613 4061 1666
rect 4074 1613 4077 1646
rect 4042 1593 4045 1606
rect 4002 1533 4013 1536
rect 4026 1536 4029 1586
rect 4034 1583 4049 1586
rect 4026 1533 4037 1536
rect 3986 1493 3989 1526
rect 4002 1466 4005 1533
rect 4002 1463 4013 1466
rect 3922 1373 3933 1376
rect 3930 1266 3933 1373
rect 3954 1333 3957 1356
rect 3962 1333 3973 1336
rect 3978 1333 3981 1416
rect 4010 1366 4013 1463
rect 4018 1403 4021 1526
rect 4034 1436 4037 1533
rect 4046 1506 4049 1583
rect 4058 1513 4061 1536
rect 4066 1523 4069 1606
rect 4082 1603 4085 1626
rect 4090 1603 4093 1616
rect 4098 1613 4101 1656
rect 4106 1603 4109 1716
rect 4114 1623 4117 1726
rect 4130 1636 4133 1656
rect 4146 1653 4149 1753
rect 4130 1633 4137 1636
rect 4122 1583 4125 1606
rect 4046 1503 4053 1506
rect 4026 1433 4037 1436
rect 4002 1363 4013 1366
rect 3890 1173 3897 1176
rect 3906 1203 3917 1206
rect 3922 1263 3933 1266
rect 3874 993 3885 996
rect 3842 933 3849 936
rect 3858 933 3861 976
rect 3882 946 3885 993
rect 3874 943 3885 946
rect 3842 916 3845 933
rect 3874 926 3877 943
rect 3834 913 3845 916
rect 3786 876 3789 896
rect 3786 873 3797 876
rect 3794 826 3797 873
rect 3786 823 3797 826
rect 3786 776 3789 823
rect 3810 816 3813 906
rect 3834 836 3837 913
rect 3850 903 3853 916
rect 3834 833 3841 836
rect 3810 813 3821 816
rect 3778 773 3789 776
rect 3754 613 3773 616
rect 3762 583 3765 606
rect 3778 603 3781 773
rect 3794 733 3797 746
rect 3786 706 3789 726
rect 3786 703 3793 706
rect 3790 636 3793 703
rect 3802 673 3805 806
rect 3818 756 3821 813
rect 3838 786 3841 833
rect 3850 793 3853 806
rect 3838 783 3845 786
rect 3810 753 3821 756
rect 3810 733 3813 753
rect 3810 723 3821 726
rect 3842 706 3845 783
rect 3858 746 3861 926
rect 3870 923 3877 926
rect 3890 923 3893 1173
rect 3898 1133 3901 1156
rect 3906 1133 3909 1203
rect 3914 1133 3917 1196
rect 3922 1173 3925 1263
rect 3938 1203 3941 1226
rect 3962 1193 3965 1216
rect 3930 1133 3933 1186
rect 3954 1156 3957 1176
rect 3954 1153 3961 1156
rect 3898 1003 3901 1016
rect 3906 1003 3909 1126
rect 3922 1123 3933 1126
rect 3938 1113 3941 1126
rect 3946 1096 3949 1136
rect 3942 1093 3949 1096
rect 3914 1013 3917 1056
rect 3930 1013 3933 1036
rect 3914 1003 3925 1006
rect 3914 923 3917 1003
rect 3942 976 3945 1093
rect 3958 1086 3961 1153
rect 3970 1133 3973 1326
rect 4002 1266 4005 1363
rect 4026 1333 4029 1433
rect 4050 1426 4053 1503
rect 4050 1423 4061 1426
rect 4026 1306 4029 1326
rect 4034 1313 4037 1416
rect 4042 1363 4045 1416
rect 4058 1366 4061 1423
rect 4050 1363 4061 1366
rect 4050 1336 4053 1363
rect 4074 1346 4077 1536
rect 4098 1526 4101 1536
rect 4090 1523 4101 1526
rect 4090 1506 4093 1523
rect 4086 1503 4093 1506
rect 4086 1446 4089 1503
rect 4098 1456 4101 1516
rect 4106 1493 4109 1526
rect 4114 1483 4117 1526
rect 4098 1453 4109 1456
rect 4086 1443 4093 1446
rect 4090 1423 4093 1443
rect 4106 1423 4109 1453
rect 4122 1406 4125 1536
rect 4134 1506 4137 1633
rect 4154 1613 4157 1636
rect 4162 1613 4165 1756
rect 4186 1713 4189 1726
rect 4202 1686 4205 1763
rect 4242 1753 4245 1773
rect 4274 1766 4277 1783
rect 4274 1763 4285 1766
rect 4250 1733 4269 1736
rect 4250 1723 4253 1733
rect 4202 1683 4213 1686
rect 4146 1593 4149 1606
rect 4162 1526 4165 1606
rect 4146 1523 4165 1526
rect 4134 1503 4141 1506
rect 4138 1436 4141 1503
rect 4162 1436 4165 1516
rect 4170 1506 4173 1616
rect 4178 1523 4181 1576
rect 4186 1523 4189 1546
rect 4170 1503 4177 1506
rect 4106 1403 4125 1406
rect 4130 1433 4141 1436
rect 4154 1433 4165 1436
rect 4066 1336 4069 1346
rect 4074 1343 4085 1346
rect 4042 1333 4053 1336
rect 4042 1323 4053 1326
rect 4058 1323 4061 1336
rect 4066 1333 4077 1336
rect 4022 1303 4029 1306
rect 4002 1263 4009 1266
rect 4006 1166 4009 1263
rect 4022 1236 4025 1303
rect 4022 1233 4029 1236
rect 3994 1163 4009 1166
rect 3954 1083 3961 1086
rect 3954 986 3957 1083
rect 3962 993 3965 1006
rect 3970 1003 3973 1126
rect 3994 1056 3997 1163
rect 4018 1133 4021 1216
rect 4026 1126 4029 1233
rect 3986 1053 3997 1056
rect 4018 1123 4029 1126
rect 3954 983 3965 986
rect 3942 973 3949 976
rect 3870 836 3873 923
rect 3870 833 3877 836
rect 3874 816 3877 833
rect 3882 823 3885 906
rect 3890 896 3893 916
rect 3922 906 3925 936
rect 3946 916 3949 973
rect 3954 916 3957 926
rect 3914 903 3925 906
rect 3890 893 3901 896
rect 3898 836 3901 893
rect 3890 833 3901 836
rect 3874 813 3885 816
rect 3834 703 3845 706
rect 3854 743 3861 746
rect 3786 633 3793 636
rect 3786 613 3789 633
rect 3834 626 3837 703
rect 3854 696 3857 743
rect 3854 693 3861 696
rect 3834 623 3845 626
rect 3742 563 3749 566
rect 3742 486 3745 563
rect 3786 546 3789 586
rect 3818 556 3821 606
rect 3826 583 3829 606
rect 3818 553 3829 556
rect 3762 523 3765 546
rect 3778 543 3789 546
rect 3778 496 3781 543
rect 3810 513 3813 536
rect 3778 493 3789 496
rect 3742 483 3749 486
rect 3730 413 3733 426
rect 3746 413 3749 483
rect 3786 426 3789 493
rect 3786 423 3805 426
rect 3722 363 3729 366
rect 3690 293 3701 296
rect 3698 246 3701 293
rect 3726 286 3729 363
rect 3738 323 3741 406
rect 3746 393 3749 406
rect 3762 333 3765 346
rect 3690 243 3701 246
rect 3722 283 3729 286
rect 3690 223 3693 243
rect 3722 213 3725 283
rect 3690 166 3693 206
rect 3706 193 3709 206
rect 3674 163 3693 166
rect 3674 123 3677 163
rect 3730 156 3733 206
rect 3738 203 3741 216
rect 3754 213 3757 226
rect 3786 223 3789 416
rect 3794 323 3797 406
rect 3802 376 3805 423
rect 3810 393 3813 406
rect 3802 373 3809 376
rect 3806 316 3809 373
rect 3826 333 3829 553
rect 3842 533 3845 623
rect 3850 613 3853 676
rect 3858 603 3861 693
rect 3866 546 3869 736
rect 3882 733 3885 813
rect 3890 803 3893 833
rect 3898 763 3901 816
rect 3914 756 3917 903
rect 3930 803 3933 916
rect 3938 913 3957 916
rect 3938 903 3941 913
rect 3962 906 3965 983
rect 3954 903 3965 906
rect 3914 753 3933 756
rect 3890 733 3901 736
rect 3874 673 3877 726
rect 3890 613 3893 726
rect 3898 716 3901 733
rect 3898 713 3909 716
rect 3906 626 3909 713
rect 3898 623 3909 626
rect 3930 626 3933 753
rect 3938 733 3941 746
rect 3954 733 3957 903
rect 3970 863 3973 926
rect 3962 733 3973 736
rect 3978 733 3981 746
rect 3946 703 3949 726
rect 3954 723 3965 726
rect 3986 706 3989 1053
rect 3994 1013 3997 1046
rect 4010 1013 4013 1026
rect 4002 916 4005 1006
rect 4018 993 4021 1123
rect 4034 1106 4037 1306
rect 4042 1206 4045 1323
rect 4050 1213 4053 1316
rect 4042 1203 4053 1206
rect 4042 1133 4045 1146
rect 4050 1126 4053 1203
rect 4058 1133 4061 1196
rect 4050 1123 4061 1126
rect 4034 1103 4045 1106
rect 4026 1013 4029 1036
rect 4042 1016 4045 1103
rect 4034 1013 4045 1016
rect 4002 913 4021 916
rect 4026 913 4029 926
rect 4034 916 4037 1013
rect 4066 1006 4069 1326
rect 4082 1303 4085 1343
rect 4106 1266 4109 1403
rect 4106 1263 4121 1266
rect 4074 1133 4077 1156
rect 4082 1053 4085 1226
rect 4106 1193 4109 1216
rect 4118 1166 4121 1263
rect 4106 1163 4121 1166
rect 4090 1013 4093 1066
rect 4066 1003 4077 1006
rect 4058 933 4061 996
rect 4066 926 4069 936
rect 4066 923 4077 926
rect 4082 923 4085 1006
rect 4106 936 4109 1163
rect 4130 1136 4133 1433
rect 4138 1363 4141 1406
rect 4146 1403 4149 1416
rect 4154 1396 4157 1433
rect 4174 1426 4177 1503
rect 4146 1393 4157 1396
rect 4170 1423 4177 1426
rect 4146 1256 4149 1393
rect 4170 1376 4173 1423
rect 4186 1413 4189 1516
rect 4162 1373 4173 1376
rect 4146 1253 4153 1256
rect 4150 1176 4153 1253
rect 4162 1236 4165 1373
rect 4162 1233 4173 1236
rect 4122 1133 4133 1136
rect 4146 1173 4153 1176
rect 4146 1136 4149 1173
rect 4146 1133 4153 1136
rect 4162 1133 4165 1216
rect 4122 1116 4125 1133
rect 4118 1113 4125 1116
rect 4118 956 4121 1113
rect 4130 1003 4133 1126
rect 4118 953 4125 956
rect 4034 913 4045 916
rect 4002 823 4005 856
rect 4018 813 4021 913
rect 4026 813 4029 836
rect 4002 716 4005 736
rect 3978 703 3989 706
rect 3998 713 4005 716
rect 3930 623 3941 626
rect 3874 593 3877 606
rect 3866 543 3885 546
rect 3858 533 3869 536
rect 3858 523 3861 533
rect 3842 343 3845 516
rect 3866 356 3869 526
rect 3874 413 3877 536
rect 3882 366 3885 543
rect 3890 393 3893 536
rect 3898 523 3901 623
rect 3922 603 3933 606
rect 3938 603 3941 623
rect 3946 613 3949 676
rect 3978 626 3981 703
rect 3978 623 3989 626
rect 3938 533 3949 536
rect 3938 413 3941 526
rect 3970 443 3973 606
rect 3978 533 3981 546
rect 3986 453 3989 623
rect 3998 606 4001 713
rect 4010 613 4013 726
rect 4018 683 4021 726
rect 4026 716 4029 806
rect 4042 756 4045 913
rect 4066 886 4069 906
rect 4058 883 4069 886
rect 4058 816 4061 883
rect 4074 823 4077 923
rect 4090 826 4093 936
rect 4106 933 4113 936
rect 4098 883 4101 926
rect 4110 886 4113 933
rect 4122 903 4125 953
rect 4130 933 4133 956
rect 4138 886 4141 1126
rect 4150 1066 4153 1133
rect 4146 1063 4153 1066
rect 4146 1006 4149 1063
rect 4154 1013 4157 1046
rect 4170 1043 4173 1233
rect 4178 1176 4181 1406
rect 4194 1203 4197 1616
rect 4210 1603 4213 1683
rect 4258 1666 4261 1726
rect 4226 1613 4229 1666
rect 4250 1663 4261 1666
rect 4242 1613 4245 1646
rect 4202 1536 4205 1556
rect 4234 1553 4237 1606
rect 4250 1593 4253 1663
rect 4258 1613 4261 1636
rect 4282 1626 4285 1763
rect 4306 1733 4309 1756
rect 4322 1733 4325 1816
rect 4274 1623 4285 1626
rect 4202 1533 4209 1536
rect 4206 1446 4209 1533
rect 4218 1523 4221 1536
rect 4234 1533 4237 1546
rect 4274 1533 4277 1623
rect 4282 1593 4285 1606
rect 4234 1503 4237 1526
rect 4250 1503 4253 1526
rect 4290 1456 4293 1536
rect 4298 1523 4301 1606
rect 4306 1603 4309 1626
rect 4314 1603 4317 1726
rect 4330 1703 4333 1726
rect 4346 1713 4349 1726
rect 4354 1696 4357 1736
rect 4346 1693 4357 1696
rect 4322 1613 4325 1646
rect 4330 1593 4333 1606
rect 4346 1596 4349 1693
rect 4362 1603 4365 1916
rect 4370 1896 4373 1926
rect 4386 1913 4389 1926
rect 4370 1893 4381 1896
rect 4378 1766 4381 1893
rect 4394 1793 4397 1926
rect 4418 1923 4437 1926
rect 4434 1913 4437 1923
rect 4446 1906 4449 1953
rect 4466 1936 4469 2003
rect 4474 1943 4477 2013
rect 4482 2013 4501 2016
rect 4482 1996 4485 2013
rect 4490 2003 4501 2006
rect 4482 1993 4493 1996
rect 4458 1933 4469 1936
rect 4490 1933 4493 1993
rect 4514 1933 4517 2016
rect 4538 1993 4541 2006
rect 4522 1933 4525 1956
rect 4562 1933 4565 2016
rect 4442 1903 4449 1906
rect 4370 1763 4381 1766
rect 4370 1703 4373 1763
rect 4386 1733 4389 1746
rect 4386 1613 4389 1666
rect 4346 1593 4357 1596
rect 4306 1533 4317 1536
rect 4322 1533 4325 1566
rect 4354 1546 4357 1593
rect 4346 1543 4357 1546
rect 4314 1483 4317 1516
rect 4322 1503 4325 1516
rect 4290 1453 4301 1456
rect 4202 1443 4209 1446
rect 4202 1413 4205 1443
rect 4218 1403 4221 1426
rect 4266 1403 4269 1416
rect 4298 1396 4301 1453
rect 4346 1426 4349 1543
rect 4378 1536 4381 1606
rect 4394 1603 4397 1726
rect 4402 1596 4405 1816
rect 4410 1806 4413 1816
rect 4410 1803 4421 1806
rect 4346 1423 4357 1426
rect 4290 1393 4301 1396
rect 4226 1313 4229 1326
rect 4178 1173 4185 1176
rect 4170 1013 4173 1026
rect 4182 1016 4185 1173
rect 4194 1026 4197 1176
rect 4234 1133 4237 1216
rect 4242 1126 4245 1246
rect 4266 1223 4269 1334
rect 4282 1246 4285 1336
rect 4290 1316 4293 1393
rect 4314 1333 4317 1376
rect 4290 1313 4301 1316
rect 4278 1243 4285 1246
rect 4278 1186 4281 1243
rect 4298 1236 4301 1313
rect 4290 1233 4301 1236
rect 4278 1183 4285 1186
rect 4282 1163 4285 1183
rect 4282 1133 4285 1156
rect 4194 1023 4201 1026
rect 4182 1013 4189 1016
rect 4146 1003 4157 1006
rect 4110 883 4117 886
rect 4082 823 4093 826
rect 4058 813 4069 816
rect 4034 753 4045 756
rect 4034 733 4037 753
rect 4042 733 4053 736
rect 4026 713 4037 716
rect 3998 603 4005 606
rect 4018 603 4021 666
rect 4026 613 4029 706
rect 4034 663 4037 713
rect 4042 673 4045 726
rect 4050 716 4053 733
rect 4050 713 4057 716
rect 4054 666 4057 713
rect 4050 663 4057 666
rect 4026 603 4037 606
rect 3954 403 3957 416
rect 3882 363 3893 366
rect 3858 353 3869 356
rect 3802 313 3809 316
rect 3802 213 3805 313
rect 3842 213 3845 226
rect 3858 213 3861 353
rect 3874 323 3877 336
rect 3890 316 3893 363
rect 3874 313 3893 316
rect 3714 153 3733 156
rect 2722 0 2725 16
rect 3642 0 3645 96
rect 3714 63 3717 153
rect 3730 123 3733 136
rect 3762 123 3765 206
rect 3778 193 3781 206
rect 3818 113 3821 206
rect 3826 193 3829 206
rect 3850 146 3853 206
rect 3866 203 3869 216
rect 3874 213 3877 313
rect 3850 143 3861 146
rect 3834 123 3837 136
rect 3858 123 3861 143
rect 3746 0 3749 66
rect 3866 0 3869 116
rect 3890 0 3893 16
rect 3914 13 3917 206
rect 3930 193 3933 336
rect 3970 326 3973 346
rect 3986 336 3989 446
rect 3994 413 3997 536
rect 4002 523 4005 603
rect 4010 523 4013 536
rect 4026 513 4029 603
rect 3986 333 3993 336
rect 3962 323 3973 326
rect 3962 256 3965 323
rect 3962 253 3973 256
rect 3954 213 3957 226
rect 3970 213 3973 253
rect 3962 146 3965 206
rect 3978 203 3981 326
rect 3990 246 3993 333
rect 4002 293 4005 456
rect 4034 413 4037 536
rect 4042 533 4045 546
rect 4050 406 4053 663
rect 4066 576 4069 813
rect 4074 703 4077 726
rect 4082 716 4085 823
rect 4114 816 4117 883
rect 4106 813 4117 816
rect 4130 883 4141 886
rect 4090 733 4093 746
rect 4106 733 4109 813
rect 4130 756 4133 883
rect 4146 803 4149 926
rect 4154 853 4157 1003
rect 4162 936 4165 1006
rect 4170 1003 4181 1006
rect 4186 996 4189 1013
rect 4178 993 4189 996
rect 4162 933 4173 936
rect 4170 923 4173 933
rect 4130 753 4149 756
rect 4106 723 4117 726
rect 4082 713 4101 716
rect 4090 613 4093 676
rect 4082 583 4085 606
rect 4098 603 4101 713
rect 4106 613 4109 686
rect 4122 596 4125 736
rect 4130 703 4133 726
rect 4138 686 4141 746
rect 4146 726 4149 753
rect 4154 743 4157 806
rect 4146 723 4153 726
rect 4134 683 4141 686
rect 4134 606 4137 683
rect 4150 676 4153 723
rect 4162 683 4165 816
rect 4178 803 4181 993
rect 4186 933 4189 956
rect 4198 946 4201 1023
rect 4194 943 4201 946
rect 4194 873 4197 943
rect 4146 673 4153 676
rect 4134 603 4141 606
rect 4118 593 4125 596
rect 4066 573 4085 576
rect 4034 403 4053 406
rect 3986 243 3993 246
rect 4010 243 4013 336
rect 4026 323 4029 356
rect 4034 323 4037 403
rect 4042 323 4045 336
rect 4058 333 4061 416
rect 4066 393 4069 536
rect 4082 493 4085 573
rect 4090 533 4093 546
rect 4074 343 4077 436
rect 4090 413 4093 516
rect 4106 506 4109 536
rect 4118 526 4121 593
rect 4118 523 4125 526
rect 4106 503 4113 506
rect 4082 323 4085 406
rect 4098 396 4101 496
rect 4110 436 4113 503
rect 4106 433 4113 436
rect 4106 403 4109 433
rect 4098 393 4109 396
rect 3986 213 3989 243
rect 4042 213 4045 246
rect 4002 173 4005 206
rect 3962 143 3973 146
rect 3946 123 3949 136
rect 3970 123 3973 143
rect 4018 123 4021 206
rect 3962 0 3965 16
rect 4026 13 4029 176
rect 4058 123 4061 136
rect 4090 123 4093 226
rect 4098 186 4101 326
rect 4106 203 4109 393
rect 4122 243 4125 523
rect 4130 506 4133 586
rect 4138 523 4141 603
rect 4146 563 4149 673
rect 4170 613 4173 726
rect 4154 593 4157 606
rect 4162 583 4165 606
rect 4178 603 4181 796
rect 4186 783 4189 816
rect 4194 733 4197 806
rect 4202 793 4205 926
rect 4210 796 4213 1056
rect 4226 1013 4229 1126
rect 4234 1123 4245 1126
rect 4234 1013 4237 1076
rect 4250 1013 4253 1046
rect 4258 1033 4261 1126
rect 4242 946 4245 1006
rect 4258 1003 4261 1026
rect 4266 993 4269 1006
rect 4290 976 4293 1233
rect 4322 1226 4325 1416
rect 4330 1333 4333 1406
rect 4354 1333 4357 1423
rect 4338 1243 4341 1326
rect 4354 1266 4357 1326
rect 4346 1263 4357 1266
rect 4322 1223 4341 1226
rect 4298 1206 4301 1216
rect 4298 1203 4317 1206
rect 4298 1113 4301 1146
rect 4322 1143 4325 1216
rect 4330 1153 4333 1206
rect 4314 1113 4317 1126
rect 4234 943 4245 946
rect 4282 973 4293 976
rect 4234 923 4237 943
rect 4218 813 4221 916
rect 4242 826 4245 936
rect 4250 923 4253 936
rect 4282 906 4285 973
rect 4306 913 4309 1026
rect 4322 923 4325 1136
rect 4330 1063 4333 1126
rect 4338 1023 4341 1223
rect 4346 1096 4349 1263
rect 4362 1216 4365 1536
rect 4370 1533 4381 1536
rect 4386 1593 4405 1596
rect 4386 1533 4389 1593
rect 4394 1533 4397 1546
rect 4370 1523 4373 1533
rect 4378 1486 4381 1526
rect 4394 1503 4397 1516
rect 4378 1483 4389 1486
rect 4386 1426 4389 1483
rect 4370 1423 4389 1426
rect 4370 1223 4373 1423
rect 4378 1326 4381 1416
rect 4386 1403 4397 1406
rect 4410 1396 4413 1796
rect 4418 1733 4421 1803
rect 4426 1726 4429 1826
rect 4442 1803 4445 1903
rect 4458 1813 4461 1926
rect 4482 1913 4485 1926
rect 4458 1783 4461 1806
rect 4482 1776 4485 1816
rect 4466 1773 4485 1776
rect 4434 1733 4437 1756
rect 4466 1733 4469 1773
rect 4418 1723 4429 1726
rect 4418 1613 4421 1723
rect 4458 1676 4461 1726
rect 4474 1693 4477 1736
rect 4482 1733 4485 1746
rect 4458 1673 4469 1676
rect 4450 1613 4453 1666
rect 4466 1626 4469 1673
rect 4498 1663 4501 1926
rect 4554 1906 4557 1926
rect 4546 1903 4557 1906
rect 4546 1846 4549 1903
rect 4570 1866 4573 2026
rect 4618 2006 4621 2016
rect 4626 2013 4629 2026
rect 4618 2003 4637 2006
rect 4578 1933 4581 1966
rect 4586 1923 4589 1956
rect 4566 1863 4573 1866
rect 4546 1843 4557 1846
rect 4538 1733 4541 1816
rect 4546 1813 4549 1826
rect 4554 1733 4557 1843
rect 4566 1816 4569 1863
rect 4562 1813 4569 1816
rect 4514 1713 4517 1726
rect 4458 1623 4469 1626
rect 4426 1603 4437 1606
rect 4442 1523 4445 1606
rect 4458 1603 4461 1623
rect 4514 1613 4517 1626
rect 4530 1613 4533 1726
rect 4458 1523 4461 1536
rect 4394 1393 4413 1396
rect 4394 1333 4397 1393
rect 4418 1373 4421 1406
rect 4426 1383 4429 1516
rect 4458 1483 4461 1516
rect 4474 1426 4477 1526
rect 4482 1513 4485 1526
rect 4498 1456 4501 1526
rect 4494 1453 4501 1456
rect 4434 1336 4437 1426
rect 4474 1423 4485 1426
rect 4450 1403 4453 1416
rect 4474 1403 4477 1416
rect 4482 1336 4485 1423
rect 4494 1386 4497 1453
rect 4494 1383 4501 1386
rect 4498 1366 4501 1383
rect 4498 1363 4509 1366
rect 4378 1323 4397 1326
rect 4354 1213 4365 1216
rect 4354 1196 4357 1213
rect 4370 1203 4373 1216
rect 4378 1203 4381 1316
rect 4394 1216 4397 1323
rect 4410 1263 4413 1334
rect 4434 1333 4453 1336
rect 4434 1313 4437 1326
rect 4450 1256 4453 1333
rect 4478 1333 4485 1336
rect 4498 1333 4501 1356
rect 4450 1253 4457 1256
rect 4354 1193 4365 1196
rect 4354 1113 4357 1126
rect 4346 1093 4353 1096
rect 4350 1016 4353 1093
rect 4346 1013 4353 1016
rect 4282 903 4293 906
rect 4242 823 4253 826
rect 4210 793 4217 796
rect 4186 706 4189 726
rect 4186 703 4193 706
rect 4190 636 4193 703
rect 4202 673 4205 786
rect 4214 706 4217 793
rect 4226 733 4229 746
rect 4234 713 4237 816
rect 4250 766 4253 823
rect 4274 783 4277 806
rect 4290 803 4293 903
rect 4298 803 4301 816
rect 4242 763 4253 766
rect 4242 733 4245 763
rect 4250 733 4261 736
rect 4266 733 4269 746
rect 4274 736 4277 756
rect 4274 733 4281 736
rect 4290 733 4293 796
rect 4306 753 4309 816
rect 4298 733 4309 736
rect 4242 723 4253 726
rect 4214 703 4237 706
rect 4186 633 4193 636
rect 4186 613 4189 633
rect 4170 526 4173 566
rect 4162 523 4173 526
rect 4130 503 4141 506
rect 4138 436 4141 503
rect 4162 446 4165 523
rect 4194 516 4197 606
rect 4234 576 4237 703
rect 4266 683 4269 726
rect 4278 676 4281 733
rect 4274 673 4281 676
rect 4298 673 4301 726
rect 4234 573 4261 576
rect 4210 523 4213 546
rect 4186 513 4197 516
rect 4162 443 4173 446
rect 4130 433 4141 436
rect 4130 316 4133 433
rect 4138 323 4141 406
rect 4146 403 4149 416
rect 4154 413 4157 426
rect 4146 333 4149 356
rect 4162 353 4165 406
rect 4146 316 4149 326
rect 4130 313 4149 316
rect 4146 226 4149 313
rect 4138 223 4149 226
rect 4138 213 4141 223
rect 4154 216 4157 246
rect 4162 223 4165 336
rect 4170 283 4173 443
rect 4186 413 4189 513
rect 4178 393 4181 406
rect 4178 266 4181 336
rect 4170 263 4181 266
rect 4146 213 4157 216
rect 4130 196 4133 206
rect 4138 203 4149 206
rect 4130 193 4141 196
rect 4146 193 4149 203
rect 4098 183 4105 186
rect 4102 106 4105 183
rect 4098 103 4105 106
rect 4098 86 4101 103
rect 4090 83 4101 86
rect 4090 36 4093 83
rect 4090 33 4101 36
rect 4066 0 4069 16
rect 4098 13 4101 33
rect 4114 0 4117 76
rect 4138 73 4141 193
rect 4154 153 4157 206
rect 4162 203 4165 216
rect 4170 203 4173 263
rect 4178 213 4181 246
rect 4186 193 4189 206
rect 4202 203 4205 366
rect 4210 323 4213 406
rect 4234 393 4237 406
rect 4258 393 4261 573
rect 4274 566 4277 673
rect 4282 593 4285 616
rect 4306 603 4309 733
rect 4274 563 4285 566
rect 4282 466 4285 563
rect 4314 546 4317 806
rect 4322 733 4325 806
rect 4330 793 4333 936
rect 4338 913 4341 936
rect 4322 613 4325 726
rect 4330 613 4333 746
rect 4338 733 4341 756
rect 4338 683 4341 726
rect 4346 723 4349 1013
rect 4362 996 4365 1193
rect 4386 1133 4389 1216
rect 4394 1213 4405 1216
rect 4394 1173 4397 1206
rect 4402 1203 4405 1213
rect 4394 1123 4397 1156
rect 4402 1106 4405 1136
rect 4394 1103 4405 1106
rect 4410 1103 4413 1166
rect 4394 1036 4397 1103
rect 4370 1023 4373 1036
rect 4394 1033 4405 1036
rect 4402 1013 4405 1033
rect 4410 1023 4413 1036
rect 4358 993 4365 996
rect 4358 936 4361 993
rect 4358 933 4365 936
rect 4354 903 4357 916
rect 4354 733 4357 806
rect 4362 803 4365 933
rect 4370 926 4373 1006
rect 4370 923 4381 926
rect 4378 836 4381 923
rect 4394 906 4397 926
rect 4370 833 4381 836
rect 4390 903 4397 906
rect 4370 796 4373 833
rect 4378 803 4381 816
rect 4362 793 4373 796
rect 4390 796 4393 903
rect 4402 803 4405 1006
rect 4410 1003 4413 1016
rect 4418 1003 4421 1226
rect 4426 1073 4429 1126
rect 4434 1056 4437 1206
rect 4442 1116 4445 1246
rect 4454 1166 4457 1253
rect 4478 1246 4481 1333
rect 4478 1243 4485 1246
rect 4450 1163 4457 1166
rect 4450 1133 4453 1163
rect 4442 1113 4449 1116
rect 4430 1053 4437 1056
rect 4430 996 4433 1053
rect 4446 1046 4449 1113
rect 4442 1043 4449 1046
rect 4442 1023 4445 1043
rect 4458 1016 4461 1136
rect 4466 1133 4469 1216
rect 4474 1126 4477 1226
rect 4482 1133 4485 1243
rect 4490 1203 4493 1326
rect 4506 1316 4509 1363
rect 4498 1313 4509 1316
rect 4498 1243 4501 1313
rect 4498 1183 4501 1206
rect 4506 1153 4509 1306
rect 4514 1223 4517 1536
rect 4522 1533 4525 1606
rect 4530 1603 4541 1606
rect 4562 1603 4565 1813
rect 4570 1733 4573 1806
rect 4578 1723 4581 1856
rect 4602 1843 4605 1966
rect 4626 1933 4629 1996
rect 4642 1933 4645 1956
rect 4594 1813 4597 1836
rect 4586 1743 4589 1806
rect 4586 1626 4589 1736
rect 4602 1733 4605 1826
rect 4610 1793 4613 1816
rect 4594 1676 4597 1726
rect 4594 1673 4605 1676
rect 4570 1623 4589 1626
rect 4522 1513 4525 1526
rect 4530 1513 4533 1536
rect 4570 1523 4573 1623
rect 4578 1556 4581 1616
rect 4602 1613 4605 1673
rect 4594 1586 4597 1606
rect 4594 1583 4601 1586
rect 4578 1553 4589 1556
rect 4586 1533 4589 1553
rect 4598 1526 4601 1583
rect 4522 1303 4525 1506
rect 4578 1456 4581 1526
rect 4554 1453 4581 1456
rect 4594 1523 4601 1526
rect 4530 1406 4533 1416
rect 4538 1413 4541 1426
rect 4530 1403 4549 1406
rect 4466 1113 4469 1126
rect 4474 1123 4481 1126
rect 4478 1046 4481 1123
rect 4478 1043 4485 1046
rect 4458 1013 4465 1016
rect 4418 993 4433 996
rect 4410 903 4413 916
rect 4390 793 4397 796
rect 4362 673 4365 793
rect 4370 733 4373 746
rect 4378 716 4381 756
rect 4394 733 4397 793
rect 4374 713 4381 716
rect 4386 713 4389 726
rect 4394 723 4405 726
rect 4374 626 4377 713
rect 4374 623 4381 626
rect 4314 543 4325 546
rect 4314 516 4317 536
rect 4322 523 4325 543
rect 4274 463 4285 466
rect 4306 513 4317 516
rect 4306 466 4309 513
rect 4306 463 4317 466
rect 4274 403 4277 463
rect 4282 413 4285 446
rect 4314 413 4317 463
rect 4242 323 4245 356
rect 4290 333 4293 366
rect 4306 286 4309 336
rect 4314 323 4317 406
rect 4322 333 4325 376
rect 4330 366 4333 606
rect 4338 533 4341 606
rect 4354 593 4357 606
rect 4362 563 4365 616
rect 4378 603 4381 623
rect 4386 613 4389 686
rect 4362 443 4365 536
rect 4386 533 4389 606
rect 4370 506 4373 526
rect 4370 503 4381 506
rect 4346 393 4349 406
rect 4378 396 4381 503
rect 4410 456 4413 746
rect 4418 676 4421 993
rect 4434 923 4437 936
rect 4442 866 4445 1006
rect 4450 983 4453 1006
rect 4462 956 4465 1013
rect 4458 953 4465 956
rect 4450 933 4453 946
rect 4450 903 4453 916
rect 4434 863 4445 866
rect 4434 816 4437 863
rect 4430 813 4437 816
rect 4430 746 4433 813
rect 4430 743 4437 746
rect 4426 683 4429 726
rect 4418 673 4429 676
rect 4418 593 4421 606
rect 4410 453 4417 456
rect 4394 413 4397 426
rect 4370 393 4381 396
rect 4330 363 4341 366
rect 4290 283 4309 286
rect 4250 213 4253 226
rect 4290 213 4293 283
rect 4298 213 4301 236
rect 4314 213 4317 286
rect 4338 256 4341 363
rect 4330 253 4341 256
rect 4330 213 4333 253
rect 4362 223 4365 336
rect 4370 303 4373 393
rect 4394 286 4397 376
rect 4414 366 4417 453
rect 4410 363 4417 366
rect 4410 346 4413 363
rect 4402 343 4413 346
rect 4402 326 4405 343
rect 4402 323 4413 326
rect 4386 283 4397 286
rect 4386 236 4389 283
rect 4386 233 4397 236
rect 4394 213 4397 233
rect 4410 213 4413 323
rect 4426 213 4429 673
rect 4434 603 4437 743
rect 4442 713 4445 806
rect 4458 733 4461 953
rect 4466 923 4469 936
rect 4474 913 4477 1026
rect 4482 926 4485 1043
rect 4490 1026 4493 1136
rect 4506 1133 4509 1146
rect 4498 1043 4501 1126
rect 4490 1023 4501 1026
rect 4498 956 4501 1023
rect 4514 1013 4517 1206
rect 4522 1163 4525 1216
rect 4530 1026 4533 1334
rect 4538 1333 4541 1366
rect 4554 1356 4557 1453
rect 4570 1403 4573 1416
rect 4546 1353 4557 1356
rect 4538 1133 4541 1316
rect 4546 1306 4549 1353
rect 4554 1323 4557 1346
rect 4546 1303 4553 1306
rect 4550 1226 4553 1303
rect 4550 1223 4557 1226
rect 4546 1203 4549 1216
rect 4554 1046 4557 1223
rect 4562 1213 4565 1386
rect 4594 1343 4597 1523
rect 4578 1333 4589 1336
rect 4602 1326 4605 1426
rect 4610 1333 4613 1746
rect 4618 1613 4621 1926
rect 4626 1776 4629 1846
rect 4634 1786 4637 1926
rect 4642 1803 4645 1916
rect 4650 1813 4653 1856
rect 4634 1783 4645 1786
rect 4626 1773 4637 1776
rect 4642 1773 4645 1783
rect 4626 1733 4629 1766
rect 4634 1656 4637 1773
rect 4642 1706 4645 1736
rect 4650 1733 4653 1806
rect 4658 1733 4661 1936
rect 4674 1923 4677 1946
rect 4706 1943 4709 2006
rect 4730 1993 4733 2016
rect 4786 1933 4789 2016
rect 4698 1913 4701 1926
rect 4666 1793 4669 1816
rect 4674 1803 4677 1816
rect 4666 1733 4669 1756
rect 4650 1723 4661 1726
rect 4642 1703 4653 1706
rect 4634 1653 4641 1656
rect 4626 1503 4629 1646
rect 4638 1576 4641 1653
rect 4634 1573 4641 1576
rect 4618 1376 4621 1416
rect 4634 1383 4637 1573
rect 4650 1556 4653 1703
rect 4646 1553 4653 1556
rect 4646 1436 4649 1553
rect 4642 1433 4649 1436
rect 4642 1396 4645 1433
rect 4658 1423 4661 1536
rect 4666 1506 4669 1666
rect 4674 1533 4677 1626
rect 4666 1503 4677 1506
rect 4674 1426 4677 1503
rect 4674 1423 4685 1426
rect 4650 1406 4653 1416
rect 4650 1403 4669 1406
rect 4642 1393 4653 1396
rect 4618 1373 4637 1376
rect 4618 1333 4621 1366
rect 4586 1323 4605 1326
rect 4586 1213 4589 1323
rect 4610 1313 4613 1326
rect 4594 1196 4597 1216
rect 4586 1193 4597 1196
rect 4562 1103 4565 1126
rect 4522 1023 4533 1026
rect 4538 1043 4557 1046
rect 4490 953 4501 956
rect 4490 933 4493 953
rect 4482 923 4493 926
rect 4482 816 4485 826
rect 4474 813 4485 816
rect 4442 613 4445 676
rect 4466 673 4469 726
rect 4474 703 4477 813
rect 4482 656 4485 806
rect 4490 803 4493 923
rect 4514 916 4517 936
rect 4506 913 4517 916
rect 4506 856 4509 913
rect 4506 853 4517 856
rect 4498 813 4501 836
rect 4498 803 4509 806
rect 4506 733 4509 746
rect 4514 726 4517 853
rect 4522 733 4525 1023
rect 4538 993 4541 1043
rect 4570 1036 4573 1136
rect 4586 1133 4589 1193
rect 4554 1033 4573 1036
rect 4546 1013 4549 1026
rect 4546 976 4549 1006
rect 4538 973 4549 976
rect 4538 916 4541 973
rect 4554 923 4557 1033
rect 4578 1026 4581 1126
rect 4594 1123 4597 1156
rect 4602 1106 4605 1206
rect 4610 1156 4613 1216
rect 4618 1173 4621 1206
rect 4626 1196 4629 1336
rect 4634 1333 4637 1373
rect 4634 1203 4637 1226
rect 4642 1213 4645 1326
rect 4626 1193 4645 1196
rect 4650 1193 4653 1393
rect 4610 1153 4617 1156
rect 4570 1023 4581 1026
rect 4570 1013 4573 1023
rect 4562 1003 4573 1006
rect 4578 1003 4581 1016
rect 4586 1013 4589 1106
rect 4598 1103 4605 1106
rect 4598 1006 4601 1103
rect 4614 1096 4617 1153
rect 4642 1146 4645 1193
rect 4658 1173 4661 1386
rect 4638 1143 4645 1146
rect 4610 1093 4617 1096
rect 4610 1023 4613 1093
rect 4594 1003 4601 1006
rect 4618 1003 4621 1016
rect 4626 1003 4629 1136
rect 4638 1026 4641 1143
rect 4638 1023 4645 1026
rect 4562 976 4565 996
rect 4562 973 4573 976
rect 4538 913 4549 916
rect 4530 813 4533 826
rect 4546 813 4549 913
rect 4570 856 4573 973
rect 4562 853 4573 856
rect 4546 793 4549 806
rect 4562 803 4565 853
rect 4538 733 4541 756
rect 4546 733 4549 746
rect 4474 653 4485 656
rect 4474 606 4477 653
rect 4490 613 4493 726
rect 4506 723 4517 726
rect 4522 723 4533 726
rect 4506 676 4509 723
rect 4502 673 4509 676
rect 4502 626 4505 673
rect 4522 666 4525 723
rect 4530 696 4533 716
rect 4530 693 4541 696
rect 4514 663 4525 666
rect 4502 623 4509 626
rect 4434 423 4437 536
rect 4442 506 4445 606
rect 4450 583 4453 606
rect 4458 593 4461 606
rect 4474 603 4485 606
rect 4506 603 4509 623
rect 4514 613 4517 663
rect 4538 646 4541 693
rect 4562 683 4565 726
rect 4570 723 4573 836
rect 4578 796 4581 816
rect 4578 793 4585 796
rect 4582 716 4585 793
rect 4594 733 4597 1003
rect 4634 973 4637 1006
rect 4578 713 4585 716
rect 4530 643 4541 646
rect 4450 533 4453 556
rect 4458 533 4461 546
rect 4442 503 4449 506
rect 4446 436 4449 503
rect 4442 433 4449 436
rect 4442 413 4445 433
rect 4434 306 4437 326
rect 4458 323 4461 466
rect 4482 456 4485 603
rect 4506 546 4509 556
rect 4522 553 4525 606
rect 4530 596 4533 643
rect 4538 613 4541 626
rect 4530 593 4541 596
rect 4562 593 4565 606
rect 4578 603 4581 713
rect 4602 673 4605 726
rect 4610 656 4613 756
rect 4602 653 4613 656
rect 4586 613 4589 636
rect 4602 606 4605 653
rect 4602 603 4613 606
rect 4538 546 4541 593
rect 4506 543 4525 546
rect 4498 463 4501 526
rect 4506 516 4509 536
rect 4522 533 4525 543
rect 4530 543 4541 546
rect 4530 523 4533 543
rect 4562 533 4565 566
rect 4506 513 4517 516
rect 4482 453 4501 456
rect 4474 393 4477 406
rect 4498 396 4501 453
rect 4514 436 4517 513
rect 4538 456 4541 476
rect 4538 453 4545 456
rect 4506 433 4517 436
rect 4506 413 4509 433
rect 4498 393 4509 396
rect 4434 303 4445 306
rect 4442 246 4445 303
rect 4434 243 4445 246
rect 4162 123 4165 136
rect 4186 123 4189 156
rect 4210 0 4213 16
rect 4242 13 4245 196
rect 4290 183 4293 206
rect 4274 123 4277 136
rect 4306 123 4309 206
rect 4322 193 4325 206
rect 4354 123 4357 206
rect 4362 183 4365 206
rect 4386 123 4389 136
rect 4418 123 4421 206
rect 4434 193 4437 243
rect 4442 213 4445 226
rect 4466 223 4469 336
rect 4482 333 4485 376
rect 4506 346 4509 393
rect 4542 376 4545 453
rect 4554 406 4557 416
rect 4562 413 4565 526
rect 4570 523 4573 546
rect 4578 513 4581 586
rect 4610 583 4613 603
rect 4586 506 4589 556
rect 4594 533 4597 566
rect 4578 503 4589 506
rect 4554 403 4573 406
rect 4498 343 4509 346
rect 4538 373 4545 376
rect 4498 323 4501 343
rect 4538 313 4541 373
rect 4546 296 4549 336
rect 4538 293 4549 296
rect 4538 236 4541 293
rect 4538 233 4549 236
rect 4450 126 4453 206
rect 4466 183 4469 216
rect 4490 213 4493 226
rect 4546 213 4549 233
rect 4554 193 4557 336
rect 4562 213 4565 316
rect 4490 133 4493 186
rect 4450 123 4469 126
rect 4538 123 4541 146
rect 4570 143 4573 206
rect 4578 153 4581 503
rect 4610 466 4613 536
rect 4618 533 4621 806
rect 4626 683 4629 826
rect 4634 613 4637 816
rect 4642 803 4645 1023
rect 4650 1013 4653 1136
rect 4658 1123 4661 1166
rect 4666 1096 4669 1326
rect 4674 1313 4677 1416
rect 4674 1133 4677 1176
rect 4682 1163 4685 1423
rect 4690 1413 4693 1806
rect 4714 1803 4717 1816
rect 4754 1813 4757 1926
rect 4762 1903 4765 1926
rect 4798 1916 4801 2033
rect 4794 1913 4801 1916
rect 4794 1846 4797 1913
rect 4794 1843 4805 1846
rect 4770 1806 4773 1816
rect 4778 1813 4781 1826
rect 4770 1803 4789 1806
rect 4802 1786 4805 1843
rect 4786 1783 4805 1786
rect 4714 1646 4717 1766
rect 4714 1643 4721 1646
rect 4718 1596 4721 1643
rect 4714 1593 4721 1596
rect 4714 1533 4717 1593
rect 4730 1533 4733 1616
rect 4738 1506 4741 1776
rect 4734 1503 4741 1506
rect 4734 1436 4737 1503
rect 4746 1446 4749 1536
rect 4762 1533 4765 1736
rect 4786 1646 4789 1783
rect 4786 1643 4805 1646
rect 4770 1606 4773 1616
rect 4778 1613 4781 1626
rect 4770 1603 4789 1606
rect 4770 1456 4773 1546
rect 4802 1523 4805 1643
rect 4770 1453 4777 1456
rect 4746 1443 4753 1446
rect 4734 1433 4741 1436
rect 4706 1403 4709 1416
rect 4730 1376 4733 1416
rect 4714 1373 4733 1376
rect 4690 1333 4693 1346
rect 4698 1333 4701 1366
rect 4714 1333 4717 1373
rect 4730 1333 4733 1346
rect 4738 1336 4741 1433
rect 4750 1366 4753 1443
rect 4774 1386 4777 1453
rect 4746 1363 4753 1366
rect 4770 1383 4777 1386
rect 4770 1363 4773 1383
rect 4746 1343 4749 1363
rect 4738 1333 4749 1336
rect 4786 1333 4789 1416
rect 4706 1323 4717 1326
rect 4698 1186 4701 1266
rect 4722 1236 4725 1326
rect 4730 1323 4741 1326
rect 4746 1256 4749 1333
rect 4742 1253 4749 1256
rect 4722 1233 4733 1236
rect 4722 1213 4725 1226
rect 4690 1183 4701 1186
rect 4674 1113 4677 1126
rect 4690 1113 4693 1183
rect 4666 1093 4677 1096
rect 4674 1036 4677 1093
rect 4666 1033 4677 1036
rect 4698 1033 4701 1136
rect 4706 1123 4709 1156
rect 4714 1133 4717 1196
rect 4730 1153 4733 1233
rect 4722 1123 4725 1146
rect 4742 1136 4745 1253
rect 4738 1133 4745 1136
rect 4666 1013 4669 1033
rect 4666 896 4669 916
rect 4658 893 4669 896
rect 4658 846 4661 893
rect 4658 843 4669 846
rect 4650 813 4653 826
rect 4650 796 4653 806
rect 4642 793 4653 796
rect 4658 793 4661 806
rect 4626 553 4629 606
rect 4642 603 4645 793
rect 4650 733 4661 736
rect 4666 733 4669 843
rect 4674 803 4677 1006
rect 4706 1005 4709 1116
rect 4738 1056 4741 1133
rect 4738 1053 4749 1056
rect 4730 1013 4733 1036
rect 4746 966 4749 1053
rect 4754 976 4757 1156
rect 4778 1133 4781 1216
rect 4754 973 4761 976
rect 4738 963 4749 966
rect 4690 886 4693 934
rect 4714 913 4717 926
rect 4690 883 4709 886
rect 4658 706 4661 726
rect 4674 723 4677 796
rect 4690 723 4693 746
rect 4698 716 4701 736
rect 4690 713 4701 716
rect 4658 703 4669 706
rect 4650 613 4653 686
rect 4658 593 4661 606
rect 4626 533 4629 546
rect 4618 473 4621 526
rect 4626 496 4629 526
rect 4634 513 4637 526
rect 4626 493 4633 496
rect 4610 463 4621 466
rect 4618 413 4621 463
rect 4630 406 4633 493
rect 4594 393 4597 406
rect 4626 403 4633 406
rect 4594 203 4597 376
rect 4610 273 4613 336
rect 4618 333 4621 346
rect 4626 296 4629 403
rect 4634 333 4637 376
rect 4642 313 4645 586
rect 4658 536 4661 556
rect 4654 533 4661 536
rect 4654 466 4657 533
rect 4654 463 4661 466
rect 4658 376 4661 463
rect 4654 373 4661 376
rect 4654 306 4657 373
rect 4650 303 4657 306
rect 4602 213 4605 226
rect 4618 213 4621 296
rect 4626 293 4637 296
rect 4634 246 4637 293
rect 4626 243 4637 246
rect 4626 223 4629 243
rect 4650 226 4653 303
rect 4666 293 4669 703
rect 4674 413 4677 536
rect 4682 513 4685 596
rect 4690 533 4693 713
rect 4706 586 4709 883
rect 4714 876 4717 906
rect 4738 903 4741 963
rect 4758 876 4761 973
rect 4770 906 4773 926
rect 4778 923 4781 1006
rect 4786 933 4789 1016
rect 4770 903 4781 906
rect 4714 873 4733 876
rect 4730 756 4733 873
rect 4754 873 4761 876
rect 4754 806 4757 873
rect 4778 836 4781 903
rect 4770 833 4781 836
rect 4770 813 4773 833
rect 4754 803 4765 806
rect 4714 753 4733 756
rect 4714 683 4717 753
rect 4722 713 4725 726
rect 4730 613 4733 736
rect 4738 733 4749 736
rect 4702 583 4709 586
rect 4702 526 4705 583
rect 4698 523 4705 526
rect 4698 393 4701 523
rect 4714 466 4717 536
rect 4722 476 4725 596
rect 4730 533 4733 546
rect 4738 536 4741 726
rect 4746 543 4749 733
rect 4754 713 4757 726
rect 4762 706 4765 803
rect 4754 703 4765 706
rect 4754 593 4757 703
rect 4786 613 4789 726
rect 4738 533 4757 536
rect 4738 513 4741 526
rect 4722 473 4733 476
rect 4714 463 4725 466
rect 4722 413 4725 463
rect 4730 406 4733 473
rect 4754 466 4757 533
rect 4746 463 4757 466
rect 4746 446 4749 463
rect 4722 403 4733 406
rect 4742 443 4749 446
rect 4682 296 4685 336
rect 4706 323 4709 346
rect 4674 293 4685 296
rect 4646 223 4653 226
rect 4570 133 4589 136
rect 4594 133 4597 196
rect 4610 193 4613 206
rect 4570 123 4573 133
rect 4602 123 4605 156
rect 4626 133 4629 206
rect 4646 166 4649 223
rect 4634 123 4637 166
rect 4646 163 4653 166
rect 4642 133 4645 146
rect 4650 113 4653 163
rect 4658 133 4661 216
rect 4674 166 4677 293
rect 4722 256 4725 403
rect 4742 376 4745 443
rect 4778 413 4781 536
rect 4742 373 4749 376
rect 4746 333 4749 373
rect 4762 333 4781 336
rect 4762 323 4765 333
rect 4770 313 4773 326
rect 4714 253 4725 256
rect 4698 193 4701 216
rect 4714 186 4717 253
rect 4762 206 4765 216
rect 4770 213 4773 226
rect 4762 203 4781 206
rect 4714 183 4725 186
rect 4674 163 4685 166
rect 4722 163 4725 183
rect 4682 133 4685 163
rect 4706 123 4709 146
rect 4762 133 4781 136
rect 4762 123 4765 133
rect 4770 113 4773 126
rect 4809 37 4829 4703
rect 4833 13 4853 4727
rect 4866 693 4869 3066
<< metal3 >>
rect 1681 4732 3254 4737
rect 1937 4722 1966 4727
rect 1961 4717 1966 4722
rect 2617 4722 2646 4727
rect 2617 4717 2622 4722
rect 1961 4712 2622 4717
rect 2089 4692 2814 4697
rect 2089 4687 2094 4692
rect 1145 4682 2094 4687
rect 2809 4687 2814 4692
rect 2809 4682 2838 4687
rect 2857 4672 2942 4677
rect 2857 4667 2862 4672
rect 2105 4662 2862 4667
rect 2937 4667 2942 4672
rect 2937 4662 3150 4667
rect 1153 4652 1238 4657
rect 1153 4647 1158 4652
rect 1129 4642 1158 4647
rect 1233 4647 1238 4652
rect 1841 4652 2086 4657
rect 1841 4647 1846 4652
rect 1233 4642 1734 4647
rect 1793 4642 1846 4647
rect 2081 4647 2086 4652
rect 2081 4642 2926 4647
rect 2921 4637 2926 4642
rect 3009 4642 3038 4647
rect 3169 4642 3366 4647
rect 3009 4637 3014 4642
rect 1073 4632 1174 4637
rect 2921 4632 3014 4637
rect 3169 4627 3174 4642
rect 241 4622 286 4627
rect 385 4622 430 4627
rect 657 4622 702 4627
rect 809 4622 854 4627
rect 921 4622 1022 4627
rect 1041 4622 1086 4627
rect 1105 4622 1134 4627
rect 1177 4622 1222 4627
rect 1857 4622 1902 4627
rect 1921 4622 2406 4627
rect 921 4617 926 4622
rect 273 4612 406 4617
rect 713 4612 798 4617
rect 273 4597 278 4612
rect 793 4607 798 4612
rect 865 4612 926 4617
rect 1017 4617 1022 4622
rect 1105 4617 1110 4622
rect 2401 4617 2406 4622
rect 2537 4622 2902 4627
rect 3145 4622 3174 4627
rect 3361 4627 3366 4642
rect 3361 4622 4046 4627
rect 2537 4617 2542 4622
rect 1017 4612 1110 4617
rect 1121 4612 1158 4617
rect 2401 4612 2542 4617
rect 3057 4612 3350 4617
rect 865 4607 870 4612
rect 793 4602 870 4607
rect 1089 4602 1142 4607
rect 1353 4602 1406 4607
rect 1465 4602 1510 4607
rect 1649 4602 1670 4607
rect 2001 4602 2046 4607
rect 2185 4602 2230 4607
rect 2313 4602 2382 4607
rect 2561 4602 2606 4607
rect 2705 4602 2750 4607
rect 2857 4602 2934 4607
rect 3281 4602 3374 4607
rect 3769 4602 3798 4607
rect 4121 4602 4166 4607
rect 4385 4602 4422 4607
rect 4481 4602 4598 4607
rect 4681 4602 4726 4607
rect 89 4592 278 4597
rect 377 4592 406 4597
rect 505 4592 614 4597
rect 937 4592 966 4597
rect 993 4592 1078 4597
rect 1153 4592 1270 4597
rect 1305 4592 1582 4597
rect 1809 4592 1958 4597
rect 2137 4592 2174 4597
rect 2577 4592 2726 4597
rect 2801 4592 2870 4597
rect 2921 4592 2942 4597
rect 3057 4592 3086 4597
rect 3201 4592 3230 4597
rect 3329 4592 3430 4597
rect 3529 4592 3598 4597
rect 3721 4592 4078 4597
rect 4217 4592 4342 4597
rect 4569 4592 4702 4597
rect 1073 4587 1158 4592
rect 2017 4587 2118 4592
rect 841 4582 862 4587
rect 1993 4582 2022 4587
rect 2113 4582 2398 4587
rect 2657 4582 2686 4587
rect 2681 4577 2686 4582
rect 2753 4582 2814 4587
rect 3569 4582 3606 4587
rect 4521 4582 4622 4587
rect 2753 4577 2758 4582
rect 3625 4577 3862 4582
rect 233 4572 270 4577
rect 465 4572 590 4577
rect 465 4567 470 4572
rect 377 4562 470 4567
rect 585 4567 590 4572
rect 1089 4572 1174 4577
rect 1889 4572 2126 4577
rect 2681 4572 2758 4577
rect 3041 4572 3318 4577
rect 3481 4572 3550 4577
rect 3601 4572 3630 4577
rect 3857 4572 4054 4577
rect 4097 4572 4190 4577
rect 1089 4567 1094 4572
rect 585 4562 718 4567
rect 977 4562 1094 4567
rect 1169 4567 1174 4572
rect 2145 4567 2262 4572
rect 3481 4567 3486 4572
rect 1169 4562 1278 4567
rect 1297 4562 1414 4567
rect 1297 4557 1302 4562
rect 257 4552 374 4557
rect 481 4552 574 4557
rect 1105 4552 1158 4557
rect 1265 4552 1302 4557
rect 1409 4557 1414 4562
rect 1753 4562 1854 4567
rect 2033 4562 2150 4567
rect 2257 4562 2334 4567
rect 3337 4562 3438 4567
rect 3457 4562 3486 4567
rect 3545 4567 3550 4572
rect 4097 4567 4102 4572
rect 3545 4562 3846 4567
rect 4017 4562 4102 4567
rect 4185 4567 4190 4572
rect 4225 4572 4374 4577
rect 4497 4572 4582 4577
rect 4225 4567 4230 4572
rect 4185 4562 4230 4567
rect 4369 4567 4374 4572
rect 4369 4562 4454 4567
rect 1753 4557 1758 4562
rect 1409 4552 1526 4557
rect 1729 4552 1758 4557
rect 1849 4557 1854 4562
rect 1897 4557 1998 4562
rect 3233 4557 3342 4562
rect 3433 4557 3438 4562
rect 3841 4557 4022 4562
rect 4473 4557 4566 4562
rect 1849 4552 1902 4557
rect 1993 4552 2022 4557
rect 257 4547 262 4552
rect 2017 4547 2022 4552
rect 2121 4552 2246 4557
rect 2321 4552 2390 4557
rect 2409 4552 2526 4557
rect 2777 4552 2806 4557
rect 2961 4552 3070 4557
rect 3105 4552 3238 4557
rect 3433 4552 3478 4557
rect 3537 4552 3590 4557
rect 3649 4552 3822 4557
rect 4041 4552 4150 4557
rect 4241 4552 4478 4557
rect 4561 4552 4590 4557
rect 2121 4547 2126 4552
rect 2409 4547 2414 4552
rect 137 4542 174 4547
rect 193 4542 262 4547
rect 305 4542 366 4547
rect 361 4537 366 4542
rect 465 4542 550 4547
rect 561 4542 606 4547
rect 729 4542 766 4547
rect 809 4542 958 4547
rect 1161 4542 1190 4547
rect 1305 4542 1398 4547
rect 1585 4542 1686 4547
rect 1761 4542 1814 4547
rect 1865 4542 1998 4547
rect 2017 4542 2126 4547
rect 2145 4542 2174 4547
rect 2353 4542 2414 4547
rect 2521 4547 2526 4552
rect 3105 4547 3110 4552
rect 3473 4547 3478 4552
rect 2521 4542 2798 4547
rect 3041 4542 3110 4547
rect 3249 4542 3462 4547
rect 3473 4542 3550 4547
rect 3577 4542 3662 4547
rect 3897 4542 4174 4547
rect 4273 4542 4438 4547
rect 4481 4542 4574 4547
rect 4617 4542 4702 4547
rect 465 4537 470 4542
rect 113 4532 222 4537
rect 361 4532 470 4537
rect 545 4537 550 4542
rect 2169 4537 2174 4542
rect 2257 4537 2358 4542
rect 3681 4537 3878 4542
rect 545 4532 614 4537
rect 1497 4532 1566 4537
rect 1729 4532 1934 4537
rect 2169 4532 2262 4537
rect 2377 4532 2510 4537
rect 745 4527 846 4532
rect 1497 4527 1502 4532
rect 209 4522 262 4527
rect 585 4522 750 4527
rect 841 4522 870 4527
rect 1001 4522 1214 4527
rect 1225 4522 1318 4527
rect 1385 4522 1438 4527
rect 1473 4522 1502 4527
rect 1561 4527 1566 4532
rect 1561 4522 1598 4527
rect 1849 4522 2078 4527
rect 2505 4517 2510 4532
rect 2689 4532 2718 4537
rect 2833 4532 2894 4537
rect 3025 4532 3054 4537
rect 3121 4532 3318 4537
rect 3393 4532 3686 4537
rect 3873 4532 3926 4537
rect 4185 4532 4350 4537
rect 4593 4532 4678 4537
rect 2689 4517 2694 4532
rect 3049 4527 3126 4532
rect 3921 4527 4190 4532
rect 2929 4522 2974 4527
rect 3433 4522 3710 4527
rect 3761 4522 3902 4527
rect 4257 4522 4462 4527
rect 89 4512 150 4517
rect 489 4512 542 4517
rect 561 4512 622 4517
rect 761 4512 918 4517
rect 961 4512 1150 4517
rect 1249 4512 1334 4517
rect 1353 4512 1630 4517
rect 1809 4512 1918 4517
rect 2137 4512 2398 4517
rect 2505 4512 2694 4517
rect 3113 4512 3198 4517
rect 3481 4512 3622 4517
rect 3689 4512 3734 4517
rect 3769 4512 3934 4517
rect 3945 4512 4046 4517
rect 4073 4512 4174 4517
rect 4377 4512 4630 4517
rect 4689 4512 4790 4517
rect 913 4507 918 4512
rect 1937 4507 2022 4512
rect 3113 4507 3118 4512
rect 129 4502 518 4507
rect 529 4502 710 4507
rect 769 4502 902 4507
rect 913 4502 1022 4507
rect 1233 4502 1310 4507
rect 1425 4502 1798 4507
rect 897 4497 902 4502
rect 1793 4497 1798 4502
rect 1881 4502 1942 4507
rect 2017 4502 2110 4507
rect 2241 4502 2486 4507
rect 2937 4502 2982 4507
rect 3065 4502 3118 4507
rect 3193 4507 3198 4512
rect 3193 4502 3222 4507
rect 3369 4502 3422 4507
rect 3601 4502 3646 4507
rect 3785 4502 3878 4507
rect 4329 4502 4414 4507
rect 1881 4497 1886 4502
rect 3417 4497 3422 4502
rect 3521 4497 3606 4502
rect 249 4492 542 4497
rect 593 4492 646 4497
rect 897 4492 1094 4497
rect 1129 4492 1214 4497
rect 1505 4492 1622 4497
rect 1793 4492 1886 4497
rect 1905 4492 2006 4497
rect 2153 4492 2470 4497
rect 3041 4492 3294 4497
rect 3417 4492 3526 4497
rect 3625 4492 3702 4497
rect 665 4487 870 4492
rect 1129 4487 1134 4492
rect 201 4482 230 4487
rect 225 4477 230 4482
rect 361 4482 670 4487
rect 865 4482 1134 4487
rect 1209 4487 1214 4492
rect 2041 4487 2134 4492
rect 1209 4482 1686 4487
rect 1969 4482 2046 4487
rect 2129 4482 2286 4487
rect 2841 4482 3118 4487
rect 3265 4482 3398 4487
rect 3545 4482 4206 4487
rect 361 4477 366 4482
rect 3113 4477 3270 4482
rect 225 4472 366 4477
rect 385 4472 414 4477
rect 409 4467 414 4472
rect 497 4472 854 4477
rect 1497 4472 1958 4477
rect 497 4467 502 4472
rect 849 4467 1502 4472
rect 1953 4467 1958 4472
rect 2057 4472 2574 4477
rect 3585 4472 3638 4477
rect 4369 4472 4446 4477
rect 2057 4467 2062 4472
rect 3017 4467 3094 4472
rect 3289 4467 3358 4472
rect 4369 4467 4374 4472
rect 409 4462 502 4467
rect 1953 4462 2062 4467
rect 2593 4462 2806 4467
rect 2825 4462 3022 4467
rect 3089 4462 3294 4467
rect 3353 4462 3422 4467
rect 3489 4462 3566 4467
rect 609 4457 694 4462
rect 2593 4457 2598 4462
rect 537 4452 614 4457
rect 689 4452 1694 4457
rect 2137 4452 2318 4457
rect 2449 4452 2598 4457
rect 2801 4452 2806 4462
rect 3489 4457 3494 4462
rect 3033 4452 3078 4457
rect 3305 4452 3342 4457
rect 3441 4452 3494 4457
rect 3561 4457 3566 4462
rect 3657 4462 3886 4467
rect 4345 4462 4374 4467
rect 4441 4467 4446 4472
rect 4441 4462 4670 4467
rect 3657 4457 3662 4462
rect 3561 4452 3662 4457
rect 3881 4457 3886 4462
rect 3881 4452 3910 4457
rect 3929 4452 4318 4457
rect 2449 4447 2454 4452
rect 2801 4447 3006 4452
rect 3681 4447 3862 4452
rect 3929 4447 3934 4452
rect 353 4442 534 4447
rect 625 4442 678 4447
rect 1713 4442 1806 4447
rect 529 4437 630 4442
rect 729 4437 798 4442
rect 1121 4437 1206 4442
rect 1497 4437 1662 4442
rect 1713 4437 1718 4442
rect 481 4432 510 4437
rect 649 4432 734 4437
rect 793 4432 1126 4437
rect 1201 4432 1230 4437
rect 1225 4427 1230 4432
rect 1329 4432 1502 4437
rect 1657 4432 1718 4437
rect 1801 4437 1806 4442
rect 1905 4442 2158 4447
rect 2425 4442 2454 4447
rect 3001 4442 3030 4447
rect 1905 4437 1910 4442
rect 3025 4437 3030 4442
rect 3129 4442 3286 4447
rect 3353 4442 3382 4447
rect 3129 4437 3134 4442
rect 1801 4432 1910 4437
rect 2121 4432 2190 4437
rect 2281 4432 2694 4437
rect 2721 4432 2846 4437
rect 2865 4432 2982 4437
rect 3025 4432 3134 4437
rect 1329 4427 1334 4432
rect 3377 4427 3382 4442
rect 3505 4442 3686 4447
rect 3857 4442 3934 4447
rect 4313 4447 4318 4452
rect 4313 4442 4430 4447
rect 4689 4442 4710 4447
rect 3505 4427 3510 4442
rect 3953 4437 4102 4442
rect 3529 4432 3958 4437
rect 4097 4432 4302 4437
rect 4529 4432 4614 4437
rect 4529 4427 4534 4432
rect 193 4422 238 4427
rect 457 4422 502 4427
rect 529 4422 558 4427
rect 625 4422 662 4427
rect 737 4422 782 4427
rect 1041 4422 1070 4427
rect 1065 4417 1070 4422
rect 1137 4422 1206 4427
rect 1225 4422 1334 4427
rect 1353 4422 1382 4427
rect 1513 4422 1646 4427
rect 1745 4422 1790 4427
rect 1881 4422 1910 4427
rect 1929 4422 1950 4427
rect 1985 4422 2102 4427
rect 2177 4422 2222 4427
rect 2377 4422 2422 4427
rect 2505 4422 2550 4427
rect 2577 4422 2622 4427
rect 2745 4422 2790 4427
rect 2833 4422 2886 4427
rect 2969 4422 3006 4427
rect 3377 4422 3510 4427
rect 3929 4422 4086 4427
rect 4393 4422 4446 4427
rect 4505 4422 4534 4427
rect 4609 4427 4614 4432
rect 4609 4422 4638 4427
rect 1137 4417 1142 4422
rect 1377 4417 1518 4422
rect 1985 4417 1990 4422
rect 409 4412 438 4417
rect 545 4412 654 4417
rect 689 4412 718 4417
rect 801 4412 902 4417
rect 1065 4412 1142 4417
rect 1697 4412 1766 4417
rect 1961 4412 1990 4417
rect 2097 4417 2102 4422
rect 3729 4417 3910 4422
rect 2097 4412 2126 4417
rect 2305 4412 2470 4417
rect 2537 4412 2670 4417
rect 2913 4412 2950 4417
rect 3153 4412 3190 4417
rect 3633 4412 3734 4417
rect 3905 4412 4014 4417
rect 4473 4412 4582 4417
rect 433 4407 550 4412
rect 801 4407 806 4412
rect 257 4402 390 4407
rect 641 4402 806 4407
rect 897 4407 902 4412
rect 2145 4407 2286 4412
rect 2785 4407 2894 4412
rect 897 4402 926 4407
rect 1161 4402 1190 4407
rect 1417 4402 1494 4407
rect 1505 4402 1558 4407
rect 1681 4402 1894 4407
rect 257 4397 262 4402
rect 217 4392 262 4397
rect 385 4397 390 4402
rect 1889 4397 1894 4402
rect 1977 4402 2150 4407
rect 2281 4402 2518 4407
rect 2681 4402 2790 4407
rect 2889 4402 2926 4407
rect 2985 4402 3062 4407
rect 3569 4402 3598 4407
rect 3745 4402 4038 4407
rect 4169 4402 4374 4407
rect 1977 4397 1982 4402
rect 2609 4397 2686 4402
rect 3593 4397 3750 4402
rect 4169 4397 4174 4402
rect 385 4392 1118 4397
rect 1473 4392 1534 4397
rect 1545 4392 1606 4397
rect 1777 4392 1870 4397
rect 1889 4392 1982 4397
rect 2049 4392 2430 4397
rect 2457 4392 2614 4397
rect 2801 4392 2854 4397
rect 2873 4392 2910 4397
rect 3049 4392 3110 4397
rect 3185 4392 3214 4397
rect 3329 4392 3438 4397
rect 3505 4392 3550 4397
rect 3769 4392 3806 4397
rect 3993 4392 4086 4397
rect 4145 4392 4174 4397
rect 4369 4397 4374 4402
rect 4481 4402 4638 4407
rect 4481 4397 4486 4402
rect 4369 4392 4486 4397
rect 4497 4392 4566 4397
rect 4657 4392 4718 4397
rect 3825 4387 3942 4392
rect 4273 4387 4350 4392
rect 89 4382 238 4387
rect 273 4382 414 4387
rect 697 4382 982 4387
rect 1561 4382 1670 4387
rect 2089 4382 2342 4387
rect 2513 4382 2598 4387
rect 2673 4382 2886 4387
rect 2937 4382 3350 4387
rect 3425 4382 3494 4387
rect 3561 4382 3830 4387
rect 3937 4382 4278 4387
rect 4345 4382 4462 4387
rect 4537 4382 4574 4387
rect 4673 4382 4726 4387
rect 3489 4377 3566 4382
rect 377 4372 686 4377
rect 993 4372 1062 4377
rect 1153 4372 1206 4377
rect 2001 4372 2614 4377
rect 2641 4372 2934 4377
rect 3841 4372 3926 4377
rect 3993 4372 4110 4377
rect 4289 4372 4470 4377
rect 681 4367 998 4372
rect 3057 4367 3134 4372
rect 3593 4367 3766 4372
rect 4105 4367 4294 4372
rect 241 4362 358 4367
rect 1049 4362 1142 4367
rect 1217 4362 1310 4367
rect 1689 4362 1822 4367
rect 1953 4362 2022 4367
rect 2553 4362 2742 4367
rect 2833 4362 2862 4367
rect 2945 4362 3062 4367
rect 3129 4362 3598 4367
rect 3761 4362 3894 4367
rect 4057 4362 4086 4367
rect 4313 4362 4350 4367
rect 4361 4362 4518 4367
rect 4625 4362 4766 4367
rect 241 4357 246 4362
rect 217 4352 246 4357
rect 353 4357 358 4362
rect 489 4357 630 4362
rect 1137 4357 1222 4362
rect 353 4352 494 4357
rect 625 4352 1022 4357
rect 1689 4347 1694 4362
rect 257 4342 398 4347
rect 393 4337 398 4342
rect 505 4342 614 4347
rect 1121 4342 1158 4347
rect 1273 4342 1446 4347
rect 1577 4342 1630 4347
rect 1665 4342 1694 4347
rect 1817 4347 1822 4362
rect 2065 4357 2478 4362
rect 2857 4357 2950 4362
rect 3913 4357 4006 4362
rect 4625 4357 4630 4362
rect 1985 4352 2014 4357
rect 2041 4352 2070 4357
rect 2473 4352 2502 4357
rect 2521 4352 2686 4357
rect 2721 4352 2766 4357
rect 3073 4352 3118 4357
rect 3609 4352 3750 4357
rect 3857 4352 3918 4357
rect 4001 4352 4310 4357
rect 4417 4352 4630 4357
rect 4761 4357 4766 4362
rect 4761 4352 4790 4357
rect 2041 4347 2046 4352
rect 1817 4342 2046 4347
rect 2497 4347 2502 4352
rect 3425 4347 3590 4352
rect 2497 4342 3238 4347
rect 505 4337 510 4342
rect 3233 4337 3238 4342
rect 3401 4342 3430 4347
rect 3585 4342 3614 4347
rect 3401 4337 3406 4342
rect 3609 4337 3614 4342
rect 3705 4342 4318 4347
rect 4345 4342 4382 4347
rect 4449 4342 4558 4347
rect 3705 4337 3710 4342
rect 4553 4337 4558 4342
rect 4641 4342 4782 4347
rect 4641 4337 4646 4342
rect 249 4332 326 4337
rect 393 4332 510 4337
rect 745 4332 1150 4337
rect 1297 4332 1374 4337
rect 1545 4332 1678 4337
rect 1761 4332 1806 4337
rect 2033 4332 2126 4337
rect 2217 4332 2542 4337
rect 2705 4332 2750 4337
rect 3017 4332 3046 4337
rect 3129 4332 3214 4337
rect 3233 4332 3406 4337
rect 3425 4332 3502 4337
rect 3537 4332 3590 4337
rect 3609 4332 3710 4337
rect 3729 4332 3838 4337
rect 3897 4332 3926 4337
rect 4193 4332 4222 4337
rect 4297 4332 4334 4337
rect 4553 4332 4646 4337
rect 2121 4327 2222 4332
rect 3041 4327 3134 4332
rect 3921 4327 4198 4332
rect 241 4322 358 4327
rect 553 4322 814 4327
rect 1993 4322 2014 4327
rect 2041 4322 2102 4327
rect 2241 4322 2414 4327
rect 2529 4322 2582 4327
rect 2657 4322 2798 4327
rect 2905 4322 2966 4327
rect 3153 4322 3190 4327
rect 1777 4317 1886 4322
rect 225 4312 286 4317
rect 457 4312 502 4317
rect 697 4312 742 4317
rect 753 4312 918 4317
rect 993 4312 1078 4317
rect 1129 4312 1182 4317
rect 1321 4312 1414 4317
rect 1497 4312 1582 4317
rect 1673 4312 1782 4317
rect 1881 4312 2286 4317
rect 2369 4312 3038 4317
rect 3537 4312 4534 4317
rect 2281 4307 2374 4312
rect 489 4302 558 4307
rect 641 4302 854 4307
rect 1257 4302 1494 4307
rect 1793 4302 1870 4307
rect 1993 4302 2142 4307
rect 2217 4302 2262 4307
rect 2393 4302 2438 4307
rect 2593 4302 2622 4307
rect 2793 4302 2854 4307
rect 2897 4302 2982 4307
rect 3041 4302 3198 4307
rect 2617 4297 2798 4302
rect 3473 4297 3598 4302
rect 3689 4297 4054 4302
rect 617 4292 646 4297
rect 857 4292 1710 4297
rect 1809 4292 2038 4297
rect 2281 4292 2374 4297
rect 2817 4292 2894 4297
rect 3033 4292 3062 4297
rect 3209 4292 3478 4297
rect 3593 4292 3694 4297
rect 4049 4292 4078 4297
rect 4185 4292 4358 4297
rect 641 4287 646 4292
rect 745 4287 862 4292
rect 2057 4287 2286 4292
rect 2369 4287 2470 4292
rect 2817 4287 2822 4292
rect 3057 4287 3214 4292
rect 641 4282 750 4287
rect 1177 4282 2062 4287
rect 2465 4282 2822 4287
rect 3489 4282 3582 4287
rect 3705 4282 3838 4287
rect 3873 4282 3950 4287
rect 3977 4282 4014 4287
rect 4025 4282 4254 4287
rect 1057 4277 1158 4282
rect 769 4272 806 4277
rect 841 4272 870 4277
rect 865 4267 870 4272
rect 1033 4272 1062 4277
rect 1153 4272 2454 4277
rect 2977 4272 3470 4277
rect 3881 4272 4030 4277
rect 4081 4272 4222 4277
rect 1033 4267 1038 4272
rect 2977 4267 2982 4272
rect 3465 4267 3614 4272
rect 4241 4267 4326 4272
rect 625 4262 718 4267
rect 865 4262 1038 4267
rect 1057 4262 1814 4267
rect 1857 4262 1886 4267
rect 1929 4262 2398 4267
rect 2473 4262 2822 4267
rect 2473 4257 2478 4262
rect 281 4252 358 4257
rect 809 4252 846 4257
rect 1073 4252 1318 4257
rect 1689 4252 2286 4257
rect 2369 4252 2478 4257
rect 2817 4257 2822 4262
rect 2865 4262 2934 4267
rect 2953 4262 2982 4267
rect 3609 4262 3774 4267
rect 3793 4262 3886 4267
rect 3897 4262 4246 4267
rect 4321 4262 4390 4267
rect 2865 4257 2870 4262
rect 2817 4252 2870 4257
rect 2929 4257 2934 4262
rect 3001 4257 3446 4262
rect 3769 4257 3774 4262
rect 2929 4252 3006 4257
rect 3441 4252 3598 4257
rect 3769 4252 4118 4257
rect 281 4247 286 4252
rect 185 4242 286 4247
rect 353 4247 358 4252
rect 1313 4247 1558 4252
rect 2281 4247 2374 4252
rect 2665 4247 2782 4252
rect 4113 4247 4118 4252
rect 4217 4252 4310 4257
rect 4217 4247 4222 4252
rect 4329 4247 4398 4252
rect 353 4242 382 4247
rect 569 4242 598 4247
rect 1097 4242 1134 4247
rect 1233 4242 1294 4247
rect 1553 4242 1950 4247
rect 2121 4242 2262 4247
rect 2393 4242 2606 4247
rect 2641 4242 2670 4247
rect 2777 4242 2806 4247
rect 2881 4242 2910 4247
rect 3009 4242 3414 4247
rect 3465 4242 3558 4247
rect 3649 4242 3734 4247
rect 3769 4242 3998 4247
rect 4017 4242 4094 4247
rect 4113 4242 4222 4247
rect 4273 4242 4334 4247
rect 4393 4242 4454 4247
rect 4681 4242 4718 4247
rect 1945 4237 2126 4242
rect 2905 4237 3014 4242
rect 3553 4237 3654 4242
rect 297 4232 326 4237
rect 393 4232 654 4237
rect 1105 4232 1542 4237
rect 321 4227 398 4232
rect 1537 4227 1542 4232
rect 1681 4232 1926 4237
rect 2145 4232 2382 4237
rect 2681 4232 2814 4237
rect 3033 4232 3286 4237
rect 1681 4227 1686 4232
rect 2145 4227 2150 4232
rect 2377 4227 2686 4232
rect 3281 4227 3286 4232
rect 3385 4232 3534 4237
rect 3721 4232 3846 4237
rect 4289 4232 4382 4237
rect 4457 4232 4518 4237
rect 3385 4227 3390 4232
rect 609 4222 654 4227
rect 737 4222 758 4227
rect 833 4222 926 4227
rect 1089 4222 1190 4227
rect 1249 4222 1278 4227
rect 1321 4222 1406 4227
rect 1489 4222 1518 4227
rect 1537 4222 1686 4227
rect 1705 4222 1830 4227
rect 1841 4222 1902 4227
rect 1977 4222 2150 4227
rect 2241 4222 2286 4227
rect 2705 4222 2750 4227
rect 2817 4222 2862 4227
rect 2937 4222 3022 4227
rect 3089 4222 3150 4227
rect 3201 4222 3262 4227
rect 3281 4222 3390 4227
rect 3409 4222 3558 4227
rect 3593 4222 3646 4227
rect 3809 4222 3894 4227
rect 4241 4222 4302 4227
rect 4505 4222 4582 4227
rect 4665 4222 4710 4227
rect 1825 4217 1830 4222
rect 2817 4217 2822 4222
rect 81 4212 414 4217
rect 553 4212 582 4217
rect 673 4212 798 4217
rect 1825 4212 1998 4217
rect 2257 4212 2822 4217
rect 2865 4212 2958 4217
rect 3025 4212 3086 4217
rect 3201 4212 3230 4217
rect 3425 4212 3478 4217
rect 3497 4212 3638 4217
rect 3665 4212 3742 4217
rect 3825 4212 4206 4217
rect 4329 4212 4478 4217
rect 4497 4212 4598 4217
rect 577 4207 678 4212
rect 1697 4207 1806 4212
rect 3081 4207 3206 4212
rect 3665 4207 3670 4212
rect 785 4202 966 4207
rect 1417 4202 1702 4207
rect 1801 4202 1974 4207
rect 2009 4202 2246 4207
rect 2977 4202 3062 4207
rect 3441 4202 3670 4207
rect 3737 4207 3742 4212
rect 4329 4207 4334 4212
rect 3737 4202 3822 4207
rect 4305 4202 4334 4207
rect 4473 4207 4478 4212
rect 4473 4202 4550 4207
rect 2553 4197 2718 4202
rect 241 4192 390 4197
rect 497 4192 750 4197
rect 1057 4192 1198 4197
rect 1353 4192 1438 4197
rect 1617 4192 1646 4197
rect 1713 4192 1742 4197
rect 1785 4192 1870 4197
rect 2177 4192 2222 4197
rect 2369 4192 2478 4197
rect 2529 4192 2558 4197
rect 2713 4192 2742 4197
rect 2865 4192 2894 4197
rect 2921 4192 2974 4197
rect 3081 4192 3222 4197
rect 3241 4192 3318 4197
rect 3465 4192 3574 4197
rect 3585 4192 3606 4197
rect 3617 4192 3726 4197
rect 3849 4192 3934 4197
rect 3985 4192 4030 4197
rect 4049 4192 4110 4197
rect 4129 4192 4246 4197
rect 4265 4192 4486 4197
rect 4553 4192 4694 4197
rect 3585 4187 3590 4192
rect 4129 4187 4134 4192
rect 529 4182 558 4187
rect 553 4167 558 4182
rect 745 4182 1110 4187
rect 1441 4182 1510 4187
rect 1817 4182 1958 4187
rect 1969 4182 2358 4187
rect 2433 4182 2894 4187
rect 745 4167 750 4182
rect 2353 4177 2438 4182
rect 2889 4177 2894 4182
rect 2977 4182 3070 4187
rect 3161 4182 3590 4187
rect 3609 4182 4134 4187
rect 4241 4187 4246 4192
rect 4241 4182 4294 4187
rect 4457 4182 4606 4187
rect 4649 4182 4766 4187
rect 2977 4177 2982 4182
rect 3065 4177 3166 4182
rect 4289 4177 4462 4182
rect 1393 4172 1462 4177
rect 1769 4172 1830 4177
rect 2177 4172 2206 4177
rect 2457 4172 2862 4177
rect 2889 4172 2982 4177
rect 3185 4172 3222 4177
rect 3281 4172 3358 4177
rect 3849 4172 3894 4177
rect 3945 4172 4006 4177
rect 4073 4172 4270 4177
rect 4481 4172 4526 4177
rect 3481 4167 3758 4172
rect 4521 4167 4526 4172
rect 4633 4172 4662 4177
rect 4633 4167 4638 4172
rect 553 4162 750 4167
rect 1937 4162 2014 4167
rect 2105 4162 2310 4167
rect 2409 4162 2830 4167
rect 2841 4162 2870 4167
rect 3001 4162 3030 4167
rect 3025 4157 3030 4162
rect 3129 4162 3486 4167
rect 3753 4162 3838 4167
rect 3905 4162 4174 4167
rect 4281 4162 4502 4167
rect 4521 4162 4638 4167
rect 3129 4157 3134 4162
rect 3833 4157 3910 4162
rect 4169 4157 4286 4162
rect 769 4152 1942 4157
rect 2145 4152 2478 4157
rect 2593 4152 2798 4157
rect 3025 4152 3134 4157
rect 3217 4152 3270 4157
rect 2145 4147 2150 4152
rect 2473 4147 2598 4152
rect 3265 4147 3270 4152
rect 3337 4152 3366 4157
rect 3497 4152 3742 4157
rect 3929 4152 4150 4157
rect 3337 4147 3342 4152
rect 193 4142 230 4147
rect 1937 4142 1966 4147
rect 1961 4137 1966 4142
rect 2025 4142 2150 4147
rect 2185 4142 2366 4147
rect 2401 4142 2454 4147
rect 2617 4142 2726 4147
rect 2817 4142 2846 4147
rect 3153 4142 3246 4147
rect 3265 4142 3342 4147
rect 3449 4142 3510 4147
rect 3569 4142 3646 4147
rect 3761 4142 3862 4147
rect 3889 4142 3974 4147
rect 4081 4142 4134 4147
rect 4185 4142 4286 4147
rect 2025 4137 2030 4142
rect 2721 4137 2822 4142
rect 3761 4137 3766 4142
rect 1017 4132 1078 4137
rect 1609 4132 1646 4137
rect 1657 4132 1694 4137
rect 1961 4132 2030 4137
rect 2241 4132 2470 4137
rect 2489 4132 2598 4137
rect 2649 4132 2702 4137
rect 3433 4132 3486 4137
rect 3649 4132 3766 4137
rect 3857 4137 3862 4142
rect 4185 4137 4190 4142
rect 3857 4132 3878 4137
rect 2489 4127 2494 4132
rect 153 4122 174 4127
rect 209 4122 246 4127
rect 473 4122 598 4127
rect 913 4122 950 4127
rect 961 4122 1054 4127
rect 1145 4122 1334 4127
rect 1433 4122 1526 4127
rect 1769 4122 1886 4127
rect 2185 4122 2206 4127
rect 2217 4122 2342 4127
rect 2457 4122 2494 4127
rect 2593 4127 2598 4132
rect 3873 4127 3878 4132
rect 4065 4132 4190 4137
rect 4281 4137 4286 4142
rect 4521 4142 4662 4147
rect 4521 4137 4526 4142
rect 4281 4132 4526 4137
rect 4657 4137 4662 4142
rect 4657 4132 4686 4137
rect 4065 4127 4070 4132
rect 2593 4122 2622 4127
rect 2681 4122 2806 4127
rect 3017 4122 3342 4127
rect 3529 4122 3646 4127
rect 3777 4122 3854 4127
rect 3873 4122 4070 4127
rect 4089 4122 4118 4127
rect 1521 4117 1750 4122
rect 3641 4117 3782 4122
rect 4113 4117 4118 4122
rect 4201 4122 4270 4127
rect 4625 4122 4790 4127
rect 4201 4117 4206 4122
rect 161 4112 206 4117
rect 289 4112 334 4117
rect 353 4112 454 4117
rect 497 4112 622 4117
rect 633 4112 678 4117
rect 697 4112 766 4117
rect 1009 4112 1054 4117
rect 1409 4112 1502 4117
rect 1745 4112 1870 4117
rect 2057 4112 2214 4117
rect 2249 4112 2294 4117
rect 2505 4112 2550 4117
rect 2601 4112 2670 4117
rect 2713 4112 2758 4117
rect 2825 4112 2998 4117
rect 3521 4112 3622 4117
rect 4113 4112 4206 4117
rect 4297 4112 4382 4117
rect 4505 4112 4574 4117
rect 4633 4112 4686 4117
rect 353 4107 358 4112
rect 201 4102 358 4107
rect 449 4107 454 4112
rect 697 4107 702 4112
rect 449 4102 502 4107
rect 553 4102 702 4107
rect 761 4107 766 4112
rect 2337 4107 2486 4112
rect 2825 4107 2830 4112
rect 761 4102 790 4107
rect 1073 4102 1302 4107
rect 1385 4102 1414 4107
rect 1409 4097 1414 4102
rect 1529 4102 1614 4107
rect 1633 4102 1830 4107
rect 1905 4102 2038 4107
rect 2313 4102 2342 4107
rect 2481 4102 2830 4107
rect 2993 4107 2998 4112
rect 2993 4102 3022 4107
rect 3129 4102 3374 4107
rect 3393 4102 3510 4107
rect 3745 4102 3806 4107
rect 4225 4102 4286 4107
rect 1529 4097 1534 4102
rect 1905 4097 1910 4102
rect 521 4092 558 4097
rect 809 4092 990 4097
rect 1409 4092 1534 4097
rect 1553 4092 1582 4097
rect 1809 4092 1910 4097
rect 2033 4097 2038 4102
rect 3129 4097 3134 4102
rect 2033 4092 3134 4097
rect 3369 4097 3374 4102
rect 3369 4092 3446 4097
rect 3633 4092 3734 4097
rect 809 4087 814 4092
rect 281 4082 510 4087
rect 569 4082 814 4087
rect 985 4087 990 4092
rect 1577 4087 1814 4092
rect 3441 4087 3550 4092
rect 3633 4087 3638 4092
rect 985 4082 1126 4087
rect 1281 4082 1310 4087
rect 1833 4082 2126 4087
rect 2321 4082 2558 4087
rect 2833 4082 3422 4087
rect 3545 4082 3638 4087
rect 3729 4087 3734 4092
rect 3817 4092 4094 4097
rect 3817 4087 3822 4092
rect 3729 4082 3822 4087
rect 4281 4087 4286 4102
rect 4489 4102 4518 4107
rect 4489 4087 4494 4102
rect 4529 4092 4606 4097
rect 4281 4082 4494 4087
rect 4609 4082 4654 4087
rect 505 4077 574 4082
rect 2321 4077 2326 4082
rect 2577 4077 2678 4082
rect 1145 4072 1262 4077
rect 1281 4072 1318 4077
rect 1337 4072 1534 4077
rect 913 4067 1150 4072
rect 1257 4067 1262 4072
rect 1337 4067 1342 4072
rect 361 4062 918 4067
rect 1257 4062 1342 4067
rect 1529 4067 1534 4072
rect 1617 4072 1902 4077
rect 2073 4072 2326 4077
rect 2337 4072 2390 4077
rect 2481 4072 2582 4077
rect 2673 4072 3078 4077
rect 3433 4072 3526 4077
rect 1617 4067 1622 4072
rect 1897 4067 2078 4072
rect 3073 4067 3222 4072
rect 3345 4067 3438 4072
rect 1529 4062 1622 4067
rect 2121 4062 2150 4067
rect 2305 4062 2662 4067
rect 3217 4062 3350 4067
rect 2145 4057 2310 4062
rect 2681 4057 3054 4062
rect 737 4052 766 4057
rect 937 4052 1542 4057
rect 1913 4052 2110 4057
rect 2361 4052 2438 4057
rect 2593 4052 2686 4057
rect 3049 4052 3198 4057
rect 513 4047 606 4052
rect 761 4047 942 4052
rect 2457 4047 2574 4052
rect 3193 4047 3198 4052
rect 3369 4052 3454 4057
rect 3617 4052 3702 4057
rect 3369 4047 3374 4052
rect 3617 4047 3622 4052
rect 457 4042 518 4047
rect 601 4042 718 4047
rect 1121 4042 1286 4047
rect 1553 4042 1838 4047
rect 1881 4042 1910 4047
rect 2057 4042 2462 4047
rect 2569 4042 3038 4047
rect 3193 4042 3374 4047
rect 3593 4042 3622 4047
rect 3697 4047 3702 4052
rect 4233 4052 4486 4057
rect 4513 4052 4686 4057
rect 4233 4047 4238 4052
rect 3697 4042 4238 4047
rect 4481 4047 4486 4052
rect 4481 4042 4566 4047
rect 961 4037 1070 4042
rect 1121 4037 1126 4042
rect 1281 4037 1286 4042
rect 1481 4037 1558 4042
rect 1905 4037 2062 4042
rect 161 4032 270 4037
rect 465 4032 598 4037
rect 593 4027 598 4032
rect 705 4032 814 4037
rect 833 4032 966 4037
rect 1065 4032 1126 4037
rect 1153 4032 1230 4037
rect 1281 4032 1486 4037
rect 2081 4032 2110 4037
rect 2417 4032 2878 4037
rect 2961 4032 2990 4037
rect 3545 4032 3742 4037
rect 4329 4032 4446 4037
rect 705 4027 710 4032
rect 833 4027 838 4032
rect 2873 4027 2966 4032
rect 4329 4027 4334 4032
rect 129 4022 174 4027
rect 233 4022 366 4027
rect 433 4022 478 4027
rect 545 4022 574 4027
rect 593 4022 710 4027
rect 729 4022 838 4027
rect 977 4022 1030 4027
rect 1049 4022 1166 4027
rect 1217 4022 1262 4027
rect 1505 4022 1630 4027
rect 1737 4022 1782 4027
rect 1873 4022 2510 4027
rect 2769 4022 2854 4027
rect 569 4007 574 4022
rect 729 4007 734 4022
rect 1873 4017 1878 4022
rect 2505 4017 2670 4022
rect 2769 4017 2774 4022
rect 2849 4017 2854 4022
rect 3001 4022 3174 4027
rect 3393 4022 3518 4027
rect 3569 4022 3686 4027
rect 4249 4022 4334 4027
rect 4441 4027 4446 4032
rect 4441 4022 4470 4027
rect 4673 4022 4734 4027
rect 3001 4017 3006 4022
rect 857 4012 958 4017
rect 1081 4012 1190 4017
rect 1281 4012 1438 4017
rect 1457 4012 1526 4017
rect 1593 4012 1878 4017
rect 2073 4012 2142 4017
rect 2401 4012 2486 4017
rect 2665 4012 2774 4017
rect 2801 4012 2830 4017
rect 2849 4012 3006 4017
rect 3193 4012 3374 4017
rect 3409 4012 3454 4017
rect 3553 4012 3622 4017
rect 4265 4012 4662 4017
rect 857 4007 862 4012
rect 305 4002 502 4007
rect 569 4002 734 4007
rect 801 4002 862 4007
rect 953 4007 958 4012
rect 1281 4007 1286 4012
rect 953 4002 982 4007
rect 1129 4002 1286 4007
rect 1433 4007 1438 4012
rect 1433 4002 1582 4007
rect 1665 4002 2150 4007
rect 2281 4002 2398 4007
rect 2465 4002 2510 4007
rect 2601 4002 2646 4007
rect 2793 4002 2822 4007
rect 1577 3997 1670 4002
rect 3193 3997 3198 4012
rect 769 3992 862 3997
rect 913 3992 1086 3997
rect 1305 3992 1374 3997
rect 1417 3992 1502 3997
rect 1689 3992 1718 3997
rect 1993 3992 2062 3997
rect 2169 3992 2262 3997
rect 1305 3987 1310 3992
rect 801 3982 1310 3987
rect 1369 3987 1374 3992
rect 2169 3987 2174 3992
rect 1369 3982 1406 3987
rect 1401 3977 1406 3982
rect 1513 3982 2086 3987
rect 2145 3982 2174 3987
rect 2257 3987 2262 3992
rect 2353 3992 2454 3997
rect 2529 3992 2558 3997
rect 2665 3992 2774 3997
rect 2353 3987 2358 3992
rect 2449 3987 2534 3992
rect 2665 3987 2670 3992
rect 2257 3982 2358 3987
rect 2609 3982 2670 3987
rect 2769 3987 2774 3992
rect 3025 3992 3150 3997
rect 3169 3992 3198 3997
rect 3369 3997 3374 4012
rect 3705 4002 3838 4007
rect 4025 4002 4070 4007
rect 4089 4002 4134 4007
rect 4305 4002 4382 4007
rect 3609 3997 3710 4002
rect 3833 3997 3838 4002
rect 3369 3992 3614 3997
rect 3833 3992 3862 3997
rect 3881 3992 4006 3997
rect 4505 3992 4566 3997
rect 3025 3987 3030 3992
rect 2769 3982 2894 3987
rect 3001 3982 3030 3987
rect 3145 3987 3150 3992
rect 3881 3987 3886 3992
rect 3145 3982 3334 3987
rect 3345 3982 3494 3987
rect 3553 3982 3582 3987
rect 3609 3982 3886 3987
rect 4001 3987 4006 3992
rect 4001 3982 4038 3987
rect 1513 3977 1518 3982
rect 3345 3977 3350 3982
rect 3489 3977 3494 3982
rect 281 3972 574 3977
rect 609 3972 702 3977
rect 1145 3972 1174 3977
rect 1313 3972 1358 3977
rect 1401 3972 1518 3977
rect 2081 3972 2246 3977
rect 2337 3972 2622 3977
rect 2729 3972 2758 3977
rect 2841 3972 3350 3977
rect 3393 3972 3478 3977
rect 3489 3972 3638 3977
rect 3761 3972 3894 3977
rect 4137 3972 4270 3977
rect 281 3967 286 3972
rect 257 3962 286 3967
rect 569 3967 574 3972
rect 721 3967 1078 3972
rect 2241 3967 2342 3972
rect 2753 3967 2846 3972
rect 3633 3967 3766 3972
rect 569 3962 726 3967
rect 1073 3962 1102 3967
rect 2497 3962 2526 3967
rect 2633 3962 2718 3967
rect 3041 3962 3614 3967
rect 3937 3962 4062 3967
rect 2361 3957 2462 3962
rect 2521 3957 2638 3962
rect 2713 3957 2718 3962
rect 2865 3957 3046 3962
rect 4137 3957 4142 3972
rect 625 3952 654 3957
rect 649 3947 654 3952
rect 737 3952 950 3957
rect 1001 3952 1070 3957
rect 1105 3952 1302 3957
rect 737 3947 742 3952
rect 1297 3947 1302 3952
rect 1369 3952 2366 3957
rect 2457 3952 2486 3957
rect 2713 3952 2870 3957
rect 3065 3952 3158 3957
rect 3321 3952 3430 3957
rect 3569 3952 3606 3957
rect 3689 3952 3798 3957
rect 3817 3952 3918 3957
rect 3937 3952 4046 3957
rect 4113 3952 4142 3957
rect 4265 3957 4270 3972
rect 4313 3972 4486 3977
rect 4689 3972 4726 3977
rect 4313 3957 4318 3972
rect 4265 3952 4318 3957
rect 4481 3957 4486 3972
rect 4585 3962 4662 3967
rect 4481 3952 4590 3957
rect 1369 3947 1374 3952
rect 3449 3947 3518 3952
rect 3817 3947 3822 3952
rect 265 3942 558 3947
rect 649 3942 742 3947
rect 761 3942 798 3947
rect 841 3942 998 3947
rect 1033 3942 1086 3947
rect 1297 3942 1374 3947
rect 2377 3942 2454 3947
rect 2577 3942 2630 3947
rect 2889 3942 3054 3947
rect 3169 3942 3310 3947
rect 3393 3942 3454 3947
rect 3513 3942 3558 3947
rect 3617 3942 3822 3947
rect 3913 3947 3918 3952
rect 3913 3942 4510 3947
rect 4673 3942 4774 3947
rect 1801 3937 1870 3942
rect 3049 3937 3174 3942
rect 3305 3937 3398 3942
rect 3553 3937 3622 3942
rect 929 3932 1038 3937
rect 1577 3932 1614 3937
rect 1729 3932 1806 3937
rect 1865 3932 2502 3937
rect 2689 3932 2766 3937
rect 3417 3932 3502 3937
rect 3745 3932 3838 3937
rect 3881 3932 4262 3937
rect 1057 3927 1126 3932
rect 2689 3927 2694 3932
rect 537 3922 590 3927
rect 601 3922 670 3927
rect 929 3922 1062 3927
rect 1121 3922 1246 3927
rect 1553 3922 1654 3927
rect 1817 3922 1854 3927
rect 2361 3922 2398 3927
rect 2521 3922 2646 3927
rect 2665 3922 2694 3927
rect 2761 3927 2766 3932
rect 2761 3922 2814 3927
rect 2825 3922 2910 3927
rect 3129 3922 3182 3927
rect 3201 3922 3318 3927
rect 3337 3922 3406 3927
rect 3585 3922 3654 3927
rect 3825 3922 4142 3927
rect 4257 3922 4326 3927
rect 4409 3922 4534 3927
rect 2425 3917 2526 3922
rect 2641 3917 2646 3922
rect 3201 3917 3206 3922
rect 129 3912 174 3917
rect 361 3912 406 3917
rect 529 3912 814 3917
rect 1001 3912 1110 3917
rect 1409 3912 1510 3917
rect 1521 3912 1598 3917
rect 1593 3907 1598 3912
rect 1665 3912 1702 3917
rect 1865 3912 1998 3917
rect 1665 3907 1670 3912
rect 1993 3907 1998 3912
rect 2217 3912 2350 3917
rect 2409 3912 2430 3917
rect 2641 3912 2750 3917
rect 2921 3912 3206 3917
rect 3313 3917 3318 3922
rect 4137 3917 4262 3922
rect 3313 3912 4118 3917
rect 4281 3912 4470 3917
rect 4513 3912 4638 3917
rect 4649 3912 4678 3917
rect 2217 3907 2222 3912
rect 2345 3907 2414 3912
rect 2745 3907 2926 3912
rect 161 3902 262 3907
rect 281 3902 374 3907
rect 777 3902 926 3907
rect 1345 3902 1462 3907
rect 1593 3902 1670 3907
rect 1857 3902 1942 3907
rect 1993 3902 2222 3907
rect 2441 3902 2502 3907
rect 2561 3902 2678 3907
rect 3161 3902 3246 3907
rect 3273 3902 3358 3907
rect 3585 3902 3614 3907
rect 3801 3902 3838 3907
rect 3881 3902 3966 3907
rect 4033 3902 4086 3907
rect 4233 3902 4262 3907
rect 257 3897 262 3902
rect 4257 3897 4262 3902
rect 4361 3902 4534 3907
rect 4561 3902 4654 3907
rect 4361 3897 4366 3902
rect 257 3892 326 3897
rect 433 3892 470 3897
rect 561 3892 590 3897
rect 585 3887 590 3892
rect 681 3892 806 3897
rect 817 3892 878 3897
rect 993 3892 1030 3897
rect 1297 3892 1318 3897
rect 1361 3892 1390 3897
rect 681 3887 686 3892
rect 1385 3887 1390 3892
rect 1473 3892 1574 3897
rect 2265 3892 2422 3897
rect 2529 3892 2870 3897
rect 2889 3892 2982 3897
rect 3001 3892 3150 3897
rect 3473 3892 3814 3897
rect 4257 3892 4366 3897
rect 4385 3892 4582 3897
rect 4609 3892 4646 3897
rect 1473 3887 1478 3892
rect 2265 3887 2270 3892
rect 193 3882 254 3887
rect 585 3882 686 3887
rect 1081 3882 1278 3887
rect 1385 3882 1478 3887
rect 1913 3882 1974 3887
rect 2241 3882 2270 3887
rect 2417 3887 2422 3892
rect 2889 3887 2894 3892
rect 2417 3882 2518 3887
rect 2801 3882 2894 3887
rect 2977 3887 2982 3892
rect 3225 3887 3438 3892
rect 2977 3882 3230 3887
rect 3433 3882 3462 3887
rect 1081 3877 1086 3882
rect 1057 3872 1086 3877
rect 1273 3877 1278 3882
rect 2513 3877 2806 3882
rect 1273 3872 1318 3877
rect 1537 3872 1630 3877
rect 1729 3872 1766 3877
rect 1793 3872 1918 3877
rect 2209 3872 2430 3877
rect 2825 3872 2862 3877
rect 2897 3872 2966 3877
rect 3105 3872 3158 3877
rect 3241 3872 3486 3877
rect 2961 3867 3110 3872
rect 3153 3867 3246 3872
rect 3481 3867 3486 3872
rect 3825 3872 4038 3877
rect 4625 3872 4662 3877
rect 4673 3872 4718 3877
rect 3825 3867 3830 3872
rect 201 3862 246 3867
rect 705 3862 806 3867
rect 873 3862 1150 3867
rect 1337 3862 1518 3867
rect 705 3857 710 3862
rect 625 3852 710 3857
rect 801 3857 806 3862
rect 1337 3857 1342 3862
rect 801 3852 830 3857
rect 1025 3852 1198 3857
rect 1217 3852 1342 3857
rect 1513 3857 1518 3862
rect 1993 3862 2094 3867
rect 2481 3862 2774 3867
rect 2801 3862 2878 3867
rect 1993 3857 1998 3862
rect 1513 3852 1998 3857
rect 2089 3857 2094 3862
rect 2873 3857 2878 3862
rect 3385 3862 3414 3867
rect 3433 3862 3462 3867
rect 3481 3862 3830 3867
rect 4105 3862 4286 3867
rect 3385 3857 3390 3862
rect 2089 3852 2486 3857
rect 2873 3852 3390 3857
rect 625 3847 630 3852
rect 2481 3847 2486 3852
rect 4105 3847 4110 3862
rect 217 3842 630 3847
rect 753 3842 790 3847
rect 817 3842 1046 3847
rect 1121 3842 1158 3847
rect 2481 3842 2854 3847
rect 4081 3842 4110 3847
rect 4281 3847 4286 3862
rect 4689 3852 4726 3857
rect 4281 3842 4334 3847
rect 809 3832 910 3837
rect 1057 3832 2078 3837
rect 2153 3832 2206 3837
rect 2305 3832 2478 3837
rect 3153 3832 3246 3837
rect 3873 3832 4062 3837
rect 4073 3832 4174 3837
rect 4249 3832 4270 3837
rect 905 3827 1062 3832
rect 3153 3827 3158 3832
rect 169 3822 278 3827
rect 641 3822 886 3827
rect 1089 3822 1134 3827
rect 1945 3822 1966 3827
rect 2177 3822 2326 3827
rect 2473 3822 2598 3827
rect 2641 3822 2686 3827
rect 2969 3822 3086 3827
rect 3129 3822 3158 3827
rect 3241 3827 3246 3832
rect 3241 3822 3318 3827
rect 3449 3822 3494 3827
rect 3857 3822 3910 3827
rect 4105 3822 4238 3827
rect 4297 3822 4326 3827
rect 4401 3822 4438 3827
rect 881 3817 886 3822
rect 1985 3817 2158 3822
rect 2345 3817 2454 3822
rect 4233 3817 4302 3822
rect 881 3812 1078 3817
rect 1145 3812 1934 3817
rect 1961 3812 1990 3817
rect 2153 3812 2214 3817
rect 2265 3812 2350 3817
rect 2449 3812 2534 3817
rect 2545 3812 2814 3817
rect 3417 3812 3486 3817
rect 4065 3812 4126 3817
rect 649 3807 798 3812
rect 1073 3807 1150 3812
rect 273 3802 302 3807
rect 337 3802 654 3807
rect 793 3802 918 3807
rect 1937 3802 2742 3807
rect 3145 3802 3230 3807
rect 3473 3802 3510 3807
rect 3537 3802 3582 3807
rect 3601 3802 3702 3807
rect 3905 3802 4166 3807
rect 4681 3802 4734 3807
rect 3601 3797 3606 3802
rect 137 3792 238 3797
rect 665 3792 782 3797
rect 857 3792 910 3797
rect 937 3792 1222 3797
rect 1281 3792 1326 3797
rect 1337 3792 1374 3797
rect 1497 3792 1542 3797
rect 1553 3792 1582 3797
rect 1689 3792 1718 3797
rect 1817 3792 1886 3797
rect 1969 3792 2022 3797
rect 2209 3792 2430 3797
rect 2561 3792 2590 3797
rect 2657 3792 2806 3797
rect 2985 3792 3206 3797
rect 3393 3792 3470 3797
rect 3569 3792 3606 3797
rect 2057 3787 2150 3792
rect 2209 3787 2214 3792
rect 2425 3787 2566 3792
rect 3697 3787 3702 3802
rect 3721 3792 3806 3797
rect 3841 3792 3910 3797
rect 4097 3792 4254 3797
rect 4361 3792 4638 3797
rect 3841 3787 3846 3792
rect 169 3782 294 3787
rect 889 3782 958 3787
rect 1209 3782 1286 3787
rect 1329 3782 1414 3787
rect 1729 3782 1846 3787
rect 1937 3782 2062 3787
rect 2145 3782 2214 3787
rect 2233 3782 2262 3787
rect 2689 3782 2974 3787
rect 785 3777 870 3782
rect 977 3777 1046 3782
rect 1937 3777 1942 3782
rect 2257 3777 2406 3782
rect 2969 3777 2974 3782
rect 3217 3782 3382 3787
rect 3481 3782 3678 3787
rect 3697 3782 3846 3787
rect 4753 3782 4790 3787
rect 3217 3777 3222 3782
rect 3377 3777 3486 3782
rect 3865 3777 3990 3782
rect 321 3772 358 3777
rect 545 3772 790 3777
rect 865 3772 982 3777
rect 1041 3772 1942 3777
rect 1953 3772 2134 3777
rect 2401 3772 2422 3777
rect 2441 3772 2670 3777
rect 2969 3772 3222 3777
rect 3633 3772 3870 3777
rect 3985 3772 4414 3777
rect 1953 3767 1958 3772
rect 2441 3767 2446 3772
rect 2665 3767 2798 3772
rect 201 3762 238 3767
rect 377 3762 526 3767
rect 801 3762 1030 3767
rect 1193 3762 1214 3767
rect 1249 3762 1670 3767
rect 1825 3762 1958 3767
rect 1985 3762 2030 3767
rect 2041 3762 2102 3767
rect 2185 3762 2246 3767
rect 2313 3762 2446 3767
rect 2793 3762 2822 3767
rect 3297 3762 3374 3767
rect 3449 3762 3574 3767
rect 3673 3762 3974 3767
rect 377 3757 382 3762
rect 313 3752 382 3757
rect 521 3757 526 3762
rect 3297 3757 3302 3762
rect 521 3752 710 3757
rect 937 3752 966 3757
rect 1241 3752 1358 3757
rect 1465 3752 1542 3757
rect 1777 3752 3302 3757
rect 3369 3757 3374 3762
rect 4001 3757 4094 3762
rect 3369 3752 3438 3757
rect 705 3747 710 3752
rect 809 3747 942 3752
rect 3433 3747 3438 3752
rect 3537 3752 4006 3757
rect 4089 3752 4230 3757
rect 4361 3752 4462 3757
rect 3537 3747 3542 3752
rect 153 3742 190 3747
rect 281 3742 334 3747
rect 361 3742 486 3747
rect 481 3737 486 3742
rect 657 3742 686 3747
rect 705 3742 814 3747
rect 1089 3742 1150 3747
rect 1249 3742 1382 3747
rect 1393 3742 1486 3747
rect 1529 3742 1574 3747
rect 1689 3742 1718 3747
rect 1729 3742 1966 3747
rect 2089 3742 2174 3747
rect 2225 3742 2294 3747
rect 2377 3742 2406 3747
rect 2505 3742 2606 3747
rect 2617 3742 2686 3747
rect 3073 3742 3134 3747
rect 3313 3742 3358 3747
rect 3433 3742 3542 3747
rect 3561 3742 3598 3747
rect 3721 3742 3758 3747
rect 3785 3742 3902 3747
rect 4017 3742 4134 3747
rect 4241 3742 4270 3747
rect 4281 3742 4406 3747
rect 4673 3742 4702 3747
rect 657 3737 662 3742
rect 1729 3737 1734 3742
rect 481 3732 662 3737
rect 833 3732 1078 3737
rect 1073 3727 1078 3732
rect 1161 3732 1238 3737
rect 1161 3727 1166 3732
rect 1073 3722 1166 3727
rect 1233 3727 1238 3732
rect 1353 3732 1734 3737
rect 1769 3732 1830 3737
rect 1921 3732 2110 3737
rect 2161 3732 2414 3737
rect 2425 3732 2494 3737
rect 2561 3732 2638 3737
rect 2713 3732 2758 3737
rect 3033 3732 3110 3737
rect 4089 3732 4126 3737
rect 4201 3732 4294 3737
rect 4513 3732 4694 3737
rect 1353 3727 1358 3732
rect 1233 3722 1358 3727
rect 1377 3722 1470 3727
rect 1529 3722 1798 3727
rect 2073 3722 2318 3727
rect 2593 3722 2670 3727
rect 2729 3722 2958 3727
rect 4041 3722 4350 3727
rect 1793 3717 1798 3722
rect 2409 3717 2478 3722
rect 4345 3717 4350 3722
rect 4417 3722 4510 3727
rect 4417 3717 4422 3722
rect 409 3712 462 3717
rect 1417 3712 1502 3717
rect 1513 3712 1566 3717
rect 1609 3712 1782 3717
rect 1793 3712 2414 3717
rect 2473 3712 2766 3717
rect 2761 3707 2766 3712
rect 2897 3712 3022 3717
rect 2897 3707 2902 3712
rect 3017 3707 3022 3712
rect 3097 3712 3126 3717
rect 3361 3712 3470 3717
rect 4113 3712 4214 3717
rect 4265 3712 4326 3717
rect 4345 3712 4422 3717
rect 3097 3707 3102 3712
rect 441 3702 846 3707
rect 937 3702 1358 3707
rect 1393 3702 1438 3707
rect 1993 3702 2086 3707
rect 2097 3702 2342 3707
rect 2425 3702 2462 3707
rect 2641 3702 2742 3707
rect 2761 3702 2902 3707
rect 2921 3702 2974 3707
rect 3017 3702 3102 3707
rect 937 3697 942 3702
rect 913 3692 942 3697
rect 1353 3697 1358 3702
rect 1633 3697 1974 3702
rect 1353 3692 1382 3697
rect 1449 3692 1638 3697
rect 1969 3692 2374 3697
rect 2585 3692 2662 3697
rect 961 3687 1246 3692
rect 1377 3687 1454 3692
rect 881 3682 966 3687
rect 1241 3682 1270 3687
rect 1649 3682 2654 3687
rect 3305 3682 4126 3687
rect 193 3672 1206 3677
rect 1281 3672 1478 3677
rect 1201 3667 1286 3672
rect 1473 3667 1478 3672
rect 1633 3672 1782 3677
rect 1633 3667 1638 3672
rect 825 3662 942 3667
rect 977 3662 1182 3667
rect 1177 3657 1182 3662
rect 1425 3662 1454 3667
rect 1473 3662 1638 3667
rect 1777 3667 1782 3672
rect 1865 3672 1966 3677
rect 1993 3672 2366 3677
rect 2409 3672 2438 3677
rect 1865 3667 1870 3672
rect 2433 3667 2438 3672
rect 2673 3672 2750 3677
rect 2857 3672 2942 3677
rect 2961 3672 3030 3677
rect 3049 3672 3158 3677
rect 3177 3672 3286 3677
rect 2673 3667 2678 3672
rect 2857 3667 2862 3672
rect 1777 3662 1870 3667
rect 2057 3662 2086 3667
rect 2281 3662 2390 3667
rect 2433 3662 2678 3667
rect 2833 3662 2862 3667
rect 2937 3667 2942 3672
rect 3049 3667 3054 3672
rect 2937 3662 3054 3667
rect 3153 3667 3158 3672
rect 3305 3667 3310 3682
rect 4121 3667 4126 3682
rect 3153 3662 3310 3667
rect 3329 3662 3806 3667
rect 4121 3662 4198 3667
rect 4425 3662 4550 3667
rect 1425 3657 1430 3662
rect 2081 3657 2286 3662
rect 3329 3657 3334 3662
rect 337 3652 406 3657
rect 337 3647 342 3652
rect 217 3642 342 3647
rect 401 3647 406 3652
rect 513 3652 614 3657
rect 1041 3652 1102 3657
rect 1177 3652 1430 3657
rect 1889 3652 1942 3657
rect 2001 3652 2054 3657
rect 3201 3652 3334 3657
rect 3801 3657 3806 3662
rect 4425 3657 4430 3662
rect 3801 3652 4110 3657
rect 4377 3652 4430 3657
rect 4545 3657 4550 3662
rect 4545 3652 4574 3657
rect 4681 3652 4758 3657
rect 513 3647 518 3652
rect 3065 3647 3182 3652
rect 3553 3647 3766 3652
rect 4681 3647 4686 3652
rect 401 3642 518 3647
rect 537 3642 782 3647
rect 873 3642 1158 3647
rect 1657 3642 1758 3647
rect 1921 3642 1958 3647
rect 2161 3642 2286 3647
rect 2841 3642 2926 3647
rect 3009 3642 3070 3647
rect 3177 3642 3262 3647
rect 3273 3642 3558 3647
rect 3761 3642 3790 3647
rect 4113 3642 4142 3647
rect 4441 3642 4534 3647
rect 4657 3642 4686 3647
rect 4753 3647 4758 3652
rect 4753 3642 4798 3647
rect 1657 3637 1662 3642
rect 353 3632 534 3637
rect 1025 3632 1110 3637
rect 1193 3632 1318 3637
rect 1633 3632 1662 3637
rect 1753 3637 1758 3642
rect 3009 3637 3014 3642
rect 3809 3637 3910 3642
rect 4017 3637 4094 3642
rect 1753 3632 1798 3637
rect 1833 3632 1998 3637
rect 2105 3632 2278 3637
rect 2537 3632 2574 3637
rect 2761 3632 2830 3637
rect 2921 3632 3014 3637
rect 3081 3632 3134 3637
rect 3145 3632 3198 3637
rect 3569 3632 3814 3637
rect 3905 3632 4022 3637
rect 4089 3632 4302 3637
rect 4481 3632 4526 3637
rect 2825 3627 2926 3632
rect 3377 3627 3486 3632
rect 137 3622 182 3627
rect 249 3622 278 3627
rect 297 3622 366 3627
rect 441 3622 486 3627
rect 505 3622 550 3627
rect 561 3622 654 3627
rect 481 3617 486 3622
rect 561 3617 566 3622
rect 89 3612 118 3617
rect 193 3612 462 3617
rect 481 3612 566 3617
rect 649 3617 654 3622
rect 737 3622 918 3627
rect 1089 3622 1134 3627
rect 1681 3622 1734 3627
rect 1785 3622 1838 3627
rect 1873 3622 1902 3627
rect 1953 3622 2094 3627
rect 2153 3622 2254 3627
rect 2569 3622 2622 3627
rect 2945 3622 3182 3627
rect 3257 3622 3382 3627
rect 3481 3622 3510 3627
rect 3585 3622 3678 3627
rect 3785 3622 3894 3627
rect 4033 3622 4134 3627
rect 4209 3622 4238 3627
rect 4313 3622 4462 3627
rect 4481 3622 4742 3627
rect 737 3617 742 3622
rect 4233 3617 4318 3622
rect 649 3612 742 3617
rect 865 3612 910 3617
rect 1065 3612 1254 3617
rect 1385 3612 1478 3617
rect 1497 3612 1630 3617
rect 1713 3612 2118 3617
rect 2361 3612 2390 3617
rect 2409 3612 2518 3617
rect 113 3607 198 3612
rect 1473 3607 1478 3612
rect 2161 3607 2310 3612
rect 2409 3607 2414 3612
rect 257 3602 374 3607
rect 761 3602 854 3607
rect 921 3602 1062 3607
rect 849 3597 926 3602
rect 1121 3597 1126 3607
rect 1137 3602 1174 3607
rect 1329 3602 1358 3607
rect 1425 3602 1462 3607
rect 1473 3602 2014 3607
rect 2129 3602 2166 3607
rect 2305 3602 2414 3607
rect 2513 3607 2518 3612
rect 2641 3612 2742 3617
rect 2897 3612 3094 3617
rect 3121 3612 3246 3617
rect 3393 3612 3454 3617
rect 4393 3612 4534 3617
rect 4609 3612 4654 3617
rect 2641 3607 2646 3612
rect 2513 3602 2646 3607
rect 2737 3607 2742 3612
rect 3241 3607 3398 3612
rect 2737 3602 3102 3607
rect 3417 3602 3462 3607
rect 3521 3602 4022 3607
rect 2009 3597 2134 3602
rect 4017 3597 4022 3602
rect 4089 3602 4422 3607
rect 4529 3602 4534 3612
rect 4089 3597 4094 3602
rect 169 3592 302 3597
rect 457 3592 510 3597
rect 577 3592 630 3597
rect 1121 3592 1318 3597
rect 1497 3592 1846 3597
rect 1945 3592 1990 3597
rect 2177 3592 2214 3597
rect 2225 3592 2294 3597
rect 2905 3592 2942 3597
rect 3009 3592 3110 3597
rect 3121 3592 3366 3597
rect 4017 3592 4094 3597
rect 4425 3592 4470 3597
rect 4649 3592 4726 3597
rect 1313 3587 1414 3592
rect 1497 3587 1502 3592
rect 2177 3587 2182 3592
rect 2409 3587 2846 3592
rect 3121 3587 3126 3592
rect 801 3582 886 3587
rect 1057 3582 1086 3587
rect 1169 3582 1198 3587
rect 1409 3582 1502 3587
rect 1521 3582 1558 3587
rect 1809 3582 2182 3587
rect 2201 3582 2238 3587
rect 2385 3582 2414 3587
rect 2841 3582 2870 3587
rect 2913 3582 2934 3587
rect 2945 3582 3126 3587
rect 3385 3582 3470 3587
rect 3505 3582 3606 3587
rect 4113 3582 4246 3587
rect 4433 3582 4518 3587
rect 1081 3577 1174 3582
rect 2945 3577 2950 3582
rect 3385 3577 3390 3582
rect 185 3572 350 3577
rect 553 3572 646 3577
rect 889 3572 1046 3577
rect 1673 3572 1710 3577
rect 1729 3572 1886 3577
rect 2201 3572 2950 3577
rect 3017 3572 3390 3577
rect 3465 3577 3470 3582
rect 4241 3577 4246 3582
rect 3465 3572 3758 3577
rect 3793 3572 3822 3577
rect 3833 3572 3862 3577
rect 4241 3572 4606 3577
rect 1881 3567 2206 3572
rect 81 3552 190 3557
rect 273 3552 326 3557
rect 161 3542 230 3547
rect 337 3537 342 3567
rect 609 3562 822 3567
rect 1097 3562 1254 3567
rect 1313 3562 1414 3567
rect 1785 3562 1862 3567
rect 2225 3562 2262 3567
rect 2377 3562 2478 3567
rect 2545 3562 3006 3567
rect 3025 3562 3150 3567
rect 3361 3562 3694 3567
rect 3761 3562 3886 3567
rect 4121 3562 4214 3567
rect 4345 3562 4638 3567
rect 1313 3557 1318 3562
rect 449 3552 486 3557
rect 601 3552 670 3557
rect 801 3552 1030 3557
rect 1073 3552 1134 3557
rect 1289 3552 1318 3557
rect 1409 3557 1414 3562
rect 4121 3557 4126 3562
rect 1409 3552 1438 3557
rect 1465 3552 1606 3557
rect 1905 3552 2022 3557
rect 2097 3552 2190 3557
rect 2313 3552 2838 3557
rect 2881 3552 3222 3557
rect 3449 3552 3598 3557
rect 3641 3552 3774 3557
rect 3825 3552 4126 3557
rect 1465 3547 1470 3552
rect 409 3542 582 3547
rect 593 3542 622 3547
rect 921 3542 950 3547
rect 1073 3542 1246 3547
rect 1409 3542 1470 3547
rect 1601 3547 1606 3552
rect 1785 3547 1886 3552
rect 4209 3547 4214 3562
rect 4257 3552 4326 3557
rect 4353 3552 4462 3557
rect 4497 3552 4518 3557
rect 4593 3552 4614 3557
rect 4257 3547 4262 3552
rect 1601 3542 1790 3547
rect 1881 3542 2390 3547
rect 2513 3542 2718 3547
rect 2977 3542 3110 3547
rect 3329 3542 3430 3547
rect 3545 3542 3630 3547
rect 3721 3542 3854 3547
rect 4137 3542 4190 3547
rect 4209 3542 4262 3547
rect 4321 3547 4326 3552
rect 4321 3542 4390 3547
rect 4425 3542 4494 3547
rect 2713 3537 2982 3542
rect 4513 3537 4518 3552
rect 4609 3547 4614 3552
rect 4545 3542 4590 3547
rect 4609 3542 4638 3547
rect 313 3532 342 3537
rect 569 3532 830 3537
rect 1225 3532 1366 3537
rect 361 3527 454 3532
rect 1361 3527 1366 3532
rect 1489 3532 1590 3537
rect 1801 3532 2542 3537
rect 2633 3532 2694 3537
rect 3001 3532 3166 3537
rect 3353 3532 3478 3537
rect 3873 3532 3910 3537
rect 4273 3532 4342 3537
rect 4497 3532 4518 3537
rect 4537 3532 4558 3537
rect 1489 3527 1494 3532
rect 2537 3527 2638 3532
rect 209 3522 366 3527
rect 449 3522 598 3527
rect 1361 3522 1494 3527
rect 2025 3522 2094 3527
rect 2169 3522 2350 3527
rect 2409 3522 2518 3527
rect 2657 3522 2806 3527
rect 2833 3522 2894 3527
rect 2961 3522 3062 3527
rect 3233 3522 3422 3527
rect 3505 3522 3790 3527
rect 4137 3522 4294 3527
rect 4497 3522 4502 3532
rect 4625 3527 4630 3537
rect 4601 3522 4630 3527
rect 1841 3517 2006 3522
rect 3121 3517 3214 3522
rect 129 3512 174 3517
rect 377 3512 422 3517
rect 521 3512 574 3517
rect 641 3512 1342 3517
rect 1609 3512 1702 3517
rect 1721 3512 1846 3517
rect 2001 3512 2206 3517
rect 2369 3512 2438 3517
rect 2521 3512 2574 3517
rect 2673 3512 2830 3517
rect 2841 3512 2886 3517
rect 3017 3512 3046 3517
rect 3081 3512 3126 3517
rect 3209 3512 3294 3517
rect 3337 3512 3438 3517
rect 3713 3512 3758 3517
rect 3769 3512 3982 3517
rect 1609 3507 1614 3512
rect 233 3502 366 3507
rect 361 3497 366 3502
rect 433 3502 614 3507
rect 1569 3502 1614 3507
rect 1697 3507 1702 3512
rect 2225 3507 2350 3512
rect 2905 3507 2998 3512
rect 4289 3507 4294 3522
rect 4353 3512 4438 3517
rect 4481 3512 4542 3517
rect 4617 3512 4710 3517
rect 4353 3507 4358 3512
rect 1697 3502 1758 3507
rect 1857 3502 2230 3507
rect 2345 3502 2910 3507
rect 2993 3502 3038 3507
rect 3161 3502 3190 3507
rect 3201 3502 3486 3507
rect 3505 3502 3694 3507
rect 3729 3502 3830 3507
rect 4153 3502 4238 3507
rect 4289 3502 4358 3507
rect 4441 3502 4654 3507
rect 433 3497 438 3502
rect 1753 3497 1862 3502
rect 3033 3497 3166 3502
rect 3505 3497 3510 3502
rect 289 3492 318 3497
rect 361 3492 438 3497
rect 513 3492 694 3497
rect 721 3492 742 3497
rect 761 3492 830 3497
rect 921 3492 1102 3497
rect 1225 3492 1262 3497
rect 1321 3492 1422 3497
rect 1545 3492 1734 3497
rect 1881 3492 2566 3497
rect 2689 3492 3014 3497
rect 3281 3492 3510 3497
rect 3689 3497 3694 3502
rect 3849 3497 4054 3502
rect 4649 3497 4654 3502
rect 4721 3502 4782 3507
rect 4721 3497 4726 3502
rect 3689 3492 3750 3497
rect 3777 3492 3854 3497
rect 4049 3492 4078 3497
rect 4505 3492 4558 3497
rect 4649 3492 4726 3497
rect 313 3477 318 3492
rect 513 3477 518 3492
rect 761 3487 766 3492
rect 545 3482 686 3487
rect 713 3482 766 3487
rect 825 3487 830 3492
rect 2585 3487 2694 3492
rect 825 3482 870 3487
rect 1065 3482 1110 3487
rect 1457 3482 1534 3487
rect 1841 3482 1918 3487
rect 1993 3482 2406 3487
rect 2449 3482 2590 3487
rect 2721 3482 4126 3487
rect 1241 3477 1438 3482
rect 1553 3477 1822 3482
rect 313 3472 518 3477
rect 537 3472 582 3477
rect 721 3472 814 3477
rect 1089 3472 1246 3477
rect 1433 3472 1558 3477
rect 1817 3472 2734 3477
rect 2857 3472 2942 3477
rect 3673 3472 3942 3477
rect 4041 3472 4070 3477
rect 2729 3467 2862 3472
rect 2937 3467 3678 3472
rect 3937 3467 4046 3472
rect 889 3462 1046 3467
rect 1257 3462 2710 3467
rect 2881 3462 2918 3467
rect 3697 3462 3726 3467
rect 3833 3462 3918 3467
rect 889 3457 894 3462
rect 1041 3457 1238 3462
rect 705 3452 758 3457
rect 793 3452 894 3457
rect 1233 3452 1678 3457
rect 1801 3452 2454 3457
rect 2561 3452 2638 3457
rect 2713 3452 2870 3457
rect 2929 3452 3646 3457
rect 945 3447 1022 3452
rect 2865 3447 2934 3452
rect 3641 3447 3646 3452
rect 3785 3452 4158 3457
rect 4177 3452 4270 3457
rect 3785 3447 3790 3452
rect 4177 3447 4182 3452
rect 153 3442 214 3447
rect 809 3442 950 3447
rect 1017 3442 1838 3447
rect 2057 3442 2646 3447
rect 3641 3442 3790 3447
rect 4145 3442 4182 3447
rect 4265 3447 4270 3452
rect 4265 3442 4430 3447
rect 4489 3442 4534 3447
rect 673 3437 790 3442
rect 1857 3437 1974 3442
rect 3265 3437 3382 3442
rect 3433 3437 3518 3442
rect 3881 3437 4022 3442
rect 649 3432 678 3437
rect 785 3432 862 3437
rect 857 3427 862 3432
rect 961 3432 1014 3437
rect 1113 3432 1862 3437
rect 1969 3432 1998 3437
rect 2009 3432 2110 3437
rect 2217 3432 2382 3437
rect 2401 3432 2494 3437
rect 2505 3432 2606 3437
rect 2729 3432 2774 3437
rect 2897 3432 2926 3437
rect 3241 3432 3270 3437
rect 3377 3432 3438 3437
rect 3513 3432 3622 3437
rect 3857 3432 3886 3437
rect 4017 3432 4046 3437
rect 961 3427 966 3432
rect 1009 3427 1118 3432
rect 4041 3427 4046 3432
rect 4113 3432 4222 3437
rect 4513 3432 4614 3437
rect 4113 3427 4118 3432
rect 4609 3427 4614 3432
rect 185 3422 230 3427
rect 265 3422 286 3427
rect 473 3422 518 3427
rect 625 3422 838 3427
rect 857 3422 966 3427
rect 1153 3422 1254 3427
rect 1265 3422 1350 3427
rect 273 3397 278 3417
rect 729 3412 750 3417
rect 441 3407 542 3412
rect 617 3407 702 3412
rect 833 3407 838 3422
rect 1265 3417 1270 3422
rect 985 3412 1270 3417
rect 1345 3417 1350 3422
rect 1465 3422 1998 3427
rect 2137 3422 2406 3427
rect 2441 3422 3366 3427
rect 1465 3417 1470 3422
rect 1993 3417 2142 3422
rect 3361 3417 3366 3422
rect 3449 3422 3486 3427
rect 3809 3422 4022 3427
rect 4041 3422 4118 3427
rect 4177 3422 4254 3427
rect 4385 3422 4438 3427
rect 4505 3422 4590 3427
rect 4609 3422 4662 3427
rect 3449 3417 3454 3422
rect 1345 3412 1470 3417
rect 1489 3412 1518 3417
rect 1777 3412 1806 3417
rect 1825 3412 1878 3417
rect 985 3407 990 3412
rect 1513 3407 1686 3412
rect 1777 3407 1782 3412
rect 377 3402 446 3407
rect 537 3402 622 3407
rect 697 3402 726 3407
rect 833 3402 990 3407
rect 1681 3402 1782 3407
rect 1873 3407 1878 3412
rect 1945 3412 1974 3417
rect 2617 3412 2670 3417
rect 3361 3412 3454 3417
rect 3905 3412 3990 3417
rect 1945 3407 1950 3412
rect 2457 3407 2598 3412
rect 1873 3402 1950 3407
rect 2089 3402 2142 3407
rect 2345 3402 2462 3407
rect 2593 3402 2894 3407
rect 3145 3402 3174 3407
rect 3193 3402 3302 3407
rect 3473 3402 3518 3407
rect 4457 3402 4582 3407
rect 3193 3397 3198 3402
rect 273 3392 294 3397
rect 321 3392 526 3397
rect 633 3392 678 3397
rect 713 3392 814 3397
rect 1009 3392 1166 3397
rect 1161 3387 1166 3392
rect 1265 3392 1326 3397
rect 1513 3392 1558 3397
rect 1265 3387 1270 3392
rect 217 3382 278 3387
rect 1161 3382 1270 3387
rect 1553 3387 1558 3392
rect 1633 3392 1662 3397
rect 1825 3392 1854 3397
rect 1633 3387 1638 3392
rect 1553 3382 1638 3387
rect 1849 3387 1854 3392
rect 1985 3392 2062 3397
rect 2473 3392 2534 3397
rect 2561 3392 2662 3397
rect 2969 3392 3198 3397
rect 3297 3397 3302 3402
rect 4457 3397 4462 3402
rect 3297 3392 3342 3397
rect 3801 3392 3934 3397
rect 4433 3392 4462 3397
rect 4577 3397 4582 3402
rect 4577 3392 4662 3397
rect 1985 3387 1990 3392
rect 1849 3382 1990 3387
rect 2329 3382 2366 3387
rect 2433 3382 2518 3387
rect 2577 3382 2750 3387
rect 2769 3382 2950 3387
rect 3097 3382 3286 3387
rect 3361 3382 3454 3387
rect 4353 3382 4566 3387
rect 2769 3377 2774 3382
rect 225 3372 286 3377
rect 297 3372 342 3377
rect 481 3372 622 3377
rect 337 3362 342 3372
rect 617 3367 622 3372
rect 729 3372 1142 3377
rect 1345 3372 1494 3377
rect 1665 3372 1750 3377
rect 2401 3372 2550 3377
rect 2633 3372 2774 3377
rect 2945 3377 2950 3382
rect 3361 3377 3366 3382
rect 2945 3372 3206 3377
rect 729 3367 734 3372
rect 1345 3367 1350 3372
rect 361 3362 454 3367
rect 617 3362 734 3367
rect 1289 3362 1350 3367
rect 1489 3367 1494 3372
rect 2545 3367 2638 3372
rect 3201 3367 3206 3372
rect 3297 3372 3366 3377
rect 3449 3377 3454 3382
rect 3449 3372 3494 3377
rect 3753 3372 3838 3377
rect 4417 3372 4574 3377
rect 4617 3372 4678 3377
rect 3297 3367 3302 3372
rect 3753 3367 3758 3372
rect 1489 3362 1534 3367
rect 2113 3362 2166 3367
rect 2497 3362 2526 3367
rect 361 3357 366 3362
rect 257 3352 366 3357
rect 449 3357 454 3362
rect 2521 3357 2526 3362
rect 2657 3362 2934 3367
rect 3201 3362 3302 3367
rect 3361 3362 3494 3367
rect 3729 3362 3758 3367
rect 3833 3367 3838 3372
rect 3833 3362 3862 3367
rect 4281 3362 4350 3367
rect 4561 3362 4678 3367
rect 2657 3357 2662 3362
rect 2929 3357 3182 3362
rect 449 3352 478 3357
rect 489 3352 590 3357
rect 1553 3352 1646 3357
rect 1889 3352 1926 3357
rect 2297 3352 2414 3357
rect 2521 3352 2662 3357
rect 2681 3352 2710 3357
rect 1553 3347 1558 3352
rect 169 3342 270 3347
rect 345 3342 430 3347
rect 513 3342 574 3347
rect 753 3342 1558 3347
rect 1641 3347 1646 3352
rect 3177 3347 3182 3357
rect 3361 3347 3366 3362
rect 3657 3352 3822 3357
rect 3873 3352 3902 3357
rect 4465 3352 4486 3357
rect 1641 3342 1774 3347
rect 1913 3342 2494 3347
rect 2809 3342 2838 3347
rect 2961 3342 3158 3347
rect 3177 3342 3366 3347
rect 3409 3342 3438 3347
rect 3585 3342 3670 3347
rect 3737 3342 3814 3347
rect 3873 3342 4110 3347
rect 4401 3342 4422 3347
rect 4537 3342 4654 3347
rect 2681 3337 2782 3342
rect 313 3332 334 3337
rect 473 3332 550 3337
rect 609 3332 734 3337
rect 1753 3332 1782 3337
rect 2129 3332 2150 3337
rect 2281 3332 2326 3337
rect 2409 3332 2438 3337
rect 353 3327 454 3332
rect 609 3327 614 3332
rect 249 3322 358 3327
rect 449 3322 614 3327
rect 729 3327 734 3332
rect 1393 3327 1486 3332
rect 729 3322 926 3327
rect 1281 3322 1398 3327
rect 1481 3322 1630 3327
rect 1801 3322 1846 3327
rect 2097 3322 2126 3327
rect 2145 3322 2150 3332
rect 2433 3327 2438 3332
rect 2505 3332 2686 3337
rect 2777 3332 2806 3337
rect 3385 3332 3438 3337
rect 3521 3332 3550 3337
rect 3633 3332 3662 3337
rect 4273 3332 4318 3337
rect 4329 3332 4398 3337
rect 2505 3327 2510 3332
rect 3545 3327 3638 3332
rect 2433 3322 2510 3327
rect 2697 3322 2846 3327
rect 2889 3322 2974 3327
rect 3481 3322 3502 3327
rect 4025 3322 4110 3327
rect 4025 3317 4030 3322
rect 137 3312 182 3317
rect 201 3312 318 3317
rect 353 3312 390 3317
rect 433 3312 486 3317
rect 569 3312 670 3317
rect 857 3312 918 3317
rect 1409 3312 1470 3317
rect 1825 3312 1870 3317
rect 1985 3312 2078 3317
rect 2185 3312 2238 3317
rect 2329 3312 2390 3317
rect 2553 3312 2598 3317
rect 2681 3312 2870 3317
rect 3049 3312 3262 3317
rect 3345 3312 3422 3317
rect 3505 3312 4030 3317
rect 4105 3317 4110 3322
rect 4129 3322 4222 3327
rect 4385 3322 4406 3327
rect 4417 3322 4422 3342
rect 4465 3332 4510 3337
rect 4561 3332 4702 3337
rect 4569 3322 4622 3327
rect 4129 3317 4134 3322
rect 4105 3312 4134 3317
rect 4217 3317 4222 3322
rect 4217 3312 4374 3317
rect 4441 3312 4470 3317
rect 4481 3312 4582 3317
rect 1985 3307 1990 3312
rect 329 3302 398 3307
rect 393 3297 398 3302
rect 497 3302 558 3307
rect 497 3297 502 3302
rect 305 3292 374 3297
rect 393 3292 502 3297
rect 553 3297 558 3302
rect 681 3302 806 3307
rect 817 3302 846 3307
rect 681 3297 686 3302
rect 553 3292 686 3297
rect 841 3297 846 3302
rect 937 3302 1238 3307
rect 1361 3302 1518 3307
rect 1801 3302 1990 3307
rect 2073 3307 2078 3312
rect 4369 3307 4446 3312
rect 2073 3302 2174 3307
rect 937 3297 942 3302
rect 2169 3297 2174 3302
rect 2249 3302 2318 3307
rect 2249 3297 2254 3302
rect 841 3292 942 3297
rect 1825 3292 1878 3297
rect 2001 3292 2070 3297
rect 2169 3292 2254 3297
rect 2313 3297 2318 3302
rect 2401 3302 2430 3307
rect 2561 3302 2662 3307
rect 3393 3302 3422 3307
rect 2401 3297 2406 3302
rect 2313 3292 2406 3297
rect 2473 3292 2510 3297
rect 3073 3292 3262 3297
rect 3417 3287 3422 3302
rect 3641 3302 3670 3307
rect 4041 3302 4094 3307
rect 4153 3302 4206 3307
rect 3641 3297 3646 3302
rect 3545 3292 3646 3297
rect 4393 3292 4518 3297
rect 4529 3292 4558 3297
rect 3545 3287 3550 3292
rect 1289 3282 1374 3287
rect 2817 3282 3054 3287
rect 3145 3282 3166 3287
rect 3321 3282 3366 3287
rect 3417 3282 3550 3287
rect 4289 3282 4350 3287
rect 4633 3282 4766 3287
rect 2817 3277 2822 3282
rect 425 3272 750 3277
rect 425 3267 430 3272
rect 257 3262 430 3267
rect 745 3267 750 3272
rect 1153 3272 1270 3277
rect 1153 3267 1158 3272
rect 745 3262 1158 3267
rect 1265 3267 1270 3272
rect 1401 3272 1526 3277
rect 1761 3272 2822 3277
rect 3049 3277 3054 3282
rect 3049 3272 3110 3277
rect 3569 3272 4278 3277
rect 1401 3267 1406 3272
rect 1265 3262 1406 3267
rect 1521 3267 1526 3272
rect 4273 3267 4278 3272
rect 4337 3272 4630 3277
rect 4337 3267 4342 3272
rect 1521 3262 1790 3267
rect 2073 3262 2134 3267
rect 2857 3262 3030 3267
rect 3177 3262 3246 3267
rect 3297 3262 3358 3267
rect 3377 3262 3470 3267
rect 4273 3262 4342 3267
rect 2857 3257 2862 3262
rect 3025 3257 3158 3262
rect 3377 3257 3382 3262
rect 265 3252 326 3257
rect 489 3252 662 3257
rect 1169 3252 1238 3257
rect 2025 3252 2126 3257
rect 2289 3252 2470 3257
rect 2833 3252 2862 3257
rect 3153 3252 3382 3257
rect 3465 3257 3470 3262
rect 3465 3252 3494 3257
rect 3649 3252 3694 3257
rect 3713 3252 3806 3257
rect 489 3247 494 3252
rect 441 3242 494 3247
rect 657 3247 662 3252
rect 2289 3247 2294 3252
rect 657 3242 734 3247
rect 1273 3242 1302 3247
rect 529 3237 622 3242
rect 1297 3237 1302 3242
rect 1417 3242 1510 3247
rect 1417 3237 1422 3242
rect 345 3232 438 3237
rect 433 3227 438 3232
rect 505 3232 534 3237
rect 617 3232 646 3237
rect 921 3232 1046 3237
rect 1113 3232 1150 3237
rect 1297 3232 1422 3237
rect 1505 3237 1510 3242
rect 1697 3242 2294 3247
rect 2465 3247 2470 3252
rect 2881 3247 2950 3252
rect 3713 3247 3718 3252
rect 2465 3242 2886 3247
rect 2945 3242 3422 3247
rect 3465 3242 3542 3247
rect 3673 3242 3718 3247
rect 3801 3247 3806 3252
rect 4481 3252 4670 3257
rect 3801 3242 3830 3247
rect 4361 3242 4382 3247
rect 1697 3237 1702 3242
rect 3561 3237 3654 3242
rect 4481 3237 4486 3252
rect 4633 3242 4678 3247
rect 1505 3232 1702 3237
rect 1721 3232 1758 3237
rect 2065 3232 2086 3237
rect 2305 3232 2454 3237
rect 2849 3232 2934 3237
rect 3193 3232 3238 3237
rect 3497 3232 3566 3237
rect 3649 3232 3742 3237
rect 3769 3232 3830 3237
rect 3977 3232 4118 3237
rect 4377 3232 4486 3237
rect 4505 3232 4710 3237
rect 505 3227 510 3232
rect 921 3227 926 3232
rect 113 3222 166 3227
rect 313 3222 358 3227
rect 433 3222 510 3227
rect 561 3222 614 3227
rect 689 3222 774 3227
rect 897 3222 926 3227
rect 1041 3227 1046 3232
rect 2953 3227 3174 3232
rect 3257 3227 3470 3232
rect 1041 3222 1070 3227
rect 2025 3222 2094 3227
rect 2273 3222 2318 3227
rect 2345 3222 2374 3227
rect 2465 3222 2630 3227
rect 2913 3222 2958 3227
rect 3169 3222 3262 3227
rect 3465 3222 3566 3227
rect 3609 3222 3654 3227
rect 3785 3222 3814 3227
rect 3841 3222 3958 3227
rect 2369 3217 2470 3222
rect 3649 3217 3790 3222
rect 3977 3217 3982 3232
rect 97 3212 270 3217
rect 529 3212 574 3217
rect 905 3212 1022 3217
rect 1041 3212 1110 3217
rect 1129 3212 1182 3217
rect 1441 3212 1486 3217
rect 2129 3212 2206 3217
rect 2521 3212 2566 3217
rect 2857 3212 2934 3217
rect 2945 3212 3342 3217
rect 3361 3212 3454 3217
rect 3609 3212 3630 3217
rect 3881 3212 3982 3217
rect 4113 3217 4118 3232
rect 4369 3222 4398 3227
rect 4113 3212 4174 3217
rect 1993 3207 2086 3212
rect 2129 3207 2134 3212
rect 857 3202 1190 3207
rect 1457 3202 1494 3207
rect 1529 3202 1590 3207
rect 1769 3202 1950 3207
rect 1969 3202 1998 3207
rect 2081 3202 2134 3207
rect 2201 3207 2206 3212
rect 4433 3207 4438 3227
rect 4657 3222 4702 3227
rect 4465 3212 4502 3217
rect 2201 3202 2358 3207
rect 2377 3202 2422 3207
rect 2649 3202 2758 3207
rect 2801 3202 2838 3207
rect 2985 3202 3022 3207
rect 3113 3202 3182 3207
rect 3201 3202 3254 3207
rect 3265 3202 3294 3207
rect 1769 3197 1774 3202
rect 113 3192 230 3197
rect 521 3192 574 3197
rect 625 3192 830 3197
rect 1001 3192 1070 3197
rect 1089 3192 1158 3197
rect 1169 3192 1254 3197
rect 1337 3192 1366 3197
rect 1521 3192 1598 3197
rect 1745 3192 1774 3197
rect 1945 3197 1950 3202
rect 2481 3197 2654 3202
rect 2753 3197 2758 3202
rect 3289 3197 3294 3202
rect 3465 3202 3630 3207
rect 3721 3202 3870 3207
rect 3921 3202 4102 3207
rect 4393 3202 4438 3207
rect 4505 3202 4598 3207
rect 3465 3197 3470 3202
rect 1945 3192 2486 3197
rect 2753 3192 2774 3197
rect 2769 3187 2774 3192
rect 2849 3192 2886 3197
rect 2849 3187 2854 3192
rect 137 3182 486 3187
rect 761 3182 814 3187
rect 1073 3182 1174 3187
rect 1385 3182 1502 3187
rect 1617 3182 1702 3187
rect 1745 3182 1766 3187
rect 1793 3182 1926 3187
rect 2041 3182 2294 3187
rect 2321 3182 2350 3187
rect 2385 3182 2422 3187
rect 2497 3182 2606 3187
rect 2617 3182 2742 3187
rect 2769 3182 2854 3187
rect 2881 3187 2886 3192
rect 3049 3192 3222 3197
rect 3289 3192 3470 3197
rect 3641 3192 3726 3197
rect 3761 3192 3982 3197
rect 4273 3192 4390 3197
rect 4425 3192 4694 3197
rect 3049 3187 3054 3192
rect 2881 3182 3054 3187
rect 3073 3182 3230 3187
rect 3625 3182 3654 3187
rect 3865 3182 3894 3187
rect 3985 3182 4046 3187
rect 4057 3182 4262 3187
rect 4521 3182 4598 3187
rect 4681 3182 4710 3187
rect 1273 3177 1390 3182
rect 1497 3177 1622 3182
rect 1697 3177 1702 3182
rect 1793 3177 1798 3182
rect 1921 3177 2022 3182
rect 3649 3177 3870 3182
rect 4257 3177 4526 3182
rect 4593 3177 4686 3182
rect 793 3172 894 3177
rect 953 3172 1278 3177
rect 1697 3172 1798 3177
rect 2017 3172 2182 3177
rect 2329 3172 2502 3177
rect 2513 3172 2702 3177
rect 3161 3172 3214 3177
rect 3361 3172 3606 3177
rect 4545 3172 4574 3177
rect 2177 3167 2334 3172
rect 2497 3167 2502 3172
rect 2721 3167 2790 3172
rect 3361 3167 3366 3172
rect 241 3162 286 3167
rect 505 3162 654 3167
rect 881 3162 942 3167
rect 1025 3162 1182 3167
rect 1289 3162 1686 3167
rect 1769 3162 2054 3167
rect 2497 3162 2726 3167
rect 2785 3162 2862 3167
rect 3289 3162 3366 3167
rect 3601 3167 3606 3172
rect 3601 3162 3702 3167
rect 3713 3162 3846 3167
rect 3857 3162 4118 3167
rect 4129 3162 4662 3167
rect 505 3157 510 3162
rect 417 3152 510 3157
rect 649 3157 654 3162
rect 937 3157 1030 3162
rect 2353 3157 2446 3162
rect 649 3152 678 3157
rect 777 3152 918 3157
rect 1049 3152 1070 3157
rect 1385 3152 1518 3157
rect 1537 3152 1598 3157
rect 1833 3152 2046 3157
rect 2065 3152 2174 3157
rect 2241 3152 2358 3157
rect 2441 3152 2774 3157
rect 1617 3147 1718 3152
rect 2065 3147 2070 3152
rect 2769 3147 2774 3152
rect 2857 3152 2886 3157
rect 3689 3152 3766 3157
rect 2857 3147 2862 3152
rect 3785 3147 4038 3152
rect 4129 3147 4134 3162
rect 4577 3152 4662 3157
rect 4209 3147 4302 3152
rect 265 3142 318 3147
rect 545 3142 646 3147
rect 665 3142 838 3147
rect 881 3142 982 3147
rect 1009 3142 1110 3147
rect 1153 3142 1190 3147
rect 1249 3142 1622 3147
rect 1713 3142 1870 3147
rect 2033 3142 2070 3147
rect 2217 3142 2270 3147
rect 2369 3142 2430 3147
rect 2505 3142 2582 3147
rect 2601 3142 2726 3147
rect 2769 3142 2862 3147
rect 3025 3142 3238 3147
rect 3377 3142 3790 3147
rect 4033 3142 4062 3147
rect 4105 3142 4134 3147
rect 4185 3142 4214 3147
rect 4297 3142 4326 3147
rect 4449 3142 4590 3147
rect 4673 3142 4734 3147
rect 3233 3137 3238 3142
rect 209 3132 254 3137
rect 249 3127 254 3132
rect 329 3132 534 3137
rect 609 3132 1046 3137
rect 1137 3132 1222 3137
rect 1441 3132 1574 3137
rect 1593 3132 1702 3137
rect 1857 3132 1974 3137
rect 2065 3132 2086 3137
rect 2121 3132 2142 3137
rect 2537 3132 2622 3137
rect 2705 3132 2750 3137
rect 3017 3132 3094 3137
rect 3233 3132 3286 3137
rect 3409 3132 3446 3137
rect 329 3127 334 3132
rect 529 3127 614 3132
rect 1041 3127 1142 3132
rect 1273 3127 1358 3132
rect 1769 3127 1838 3132
rect 2273 3127 2518 3132
rect 3441 3127 3446 3132
rect 3521 3132 3550 3137
rect 3633 3132 3686 3137
rect 3769 3132 3894 3137
rect 3913 3132 4486 3137
rect 3521 3127 3526 3132
rect 249 3122 334 3127
rect 633 3122 670 3127
rect 681 3122 750 3127
rect 873 3122 974 3127
rect 985 3122 1022 3127
rect 1161 3122 1278 3127
rect 1353 3122 1430 3127
rect 1425 3117 1430 3122
rect 1569 3122 1646 3127
rect 1713 3122 1774 3127
rect 1833 3122 2278 3127
rect 2513 3122 2838 3127
rect 2929 3122 3038 3127
rect 3361 3122 3422 3127
rect 3441 3122 3526 3127
rect 3729 3122 4126 3127
rect 4161 3122 4198 3127
rect 4281 3122 4582 3127
rect 1569 3117 1574 3122
rect 1641 3117 1718 3122
rect 4193 3117 4286 3122
rect 145 3112 174 3117
rect 473 3112 566 3117
rect 577 3112 606 3117
rect 601 3107 606 3112
rect 761 3112 822 3117
rect 985 3112 1190 3117
rect 1289 3112 1342 3117
rect 1425 3112 1574 3117
rect 1593 3112 1622 3117
rect 761 3107 766 3112
rect 1617 3107 1622 3112
rect 1785 3112 2030 3117
rect 2289 3112 2918 3117
rect 3049 3112 3270 3117
rect 3553 3112 3678 3117
rect 3745 3112 3822 3117
rect 3873 3112 3990 3117
rect 4097 3112 4174 3117
rect 4313 3112 4350 3117
rect 4401 3112 4454 3117
rect 4513 3112 4558 3117
rect 4569 3112 4606 3117
rect 4657 3112 4686 3117
rect 1785 3107 1790 3112
rect 2025 3107 2294 3112
rect 2913 3107 3054 3112
rect 241 3102 462 3107
rect 457 3097 462 3102
rect 521 3102 566 3107
rect 601 3102 766 3107
rect 1001 3102 1030 3107
rect 1161 3102 1278 3107
rect 1617 3102 1790 3107
rect 1809 3102 1862 3107
rect 1929 3102 2006 3107
rect 2313 3102 2582 3107
rect 2641 3102 2670 3107
rect 521 3097 526 3102
rect 1025 3097 1166 3102
rect 2665 3097 2670 3102
rect 2777 3102 2806 3107
rect 3665 3102 3734 3107
rect 2777 3097 2782 3102
rect 3729 3097 3734 3102
rect 3849 3102 3926 3107
rect 3849 3097 3854 3102
rect 457 3092 526 3097
rect 841 3092 926 3097
rect 1185 3092 1214 3097
rect 1249 3092 1318 3097
rect 1361 3092 1574 3097
rect 1953 3092 2078 3097
rect 2201 3092 2382 3097
rect 2401 3092 2494 3097
rect 2665 3092 2782 3097
rect 2817 3092 2910 3097
rect 2969 3092 3038 3097
rect 3729 3092 3854 3097
rect 841 3087 846 3092
rect 785 3082 846 3087
rect 921 3087 926 3092
rect 921 3082 950 3087
rect 961 3082 1022 3087
rect 1041 3082 1118 3087
rect 1153 3082 1174 3087
rect 1361 3082 1366 3092
rect 1569 3087 1574 3092
rect 1569 3082 1750 3087
rect 1041 3077 1046 3082
rect 673 3072 774 3077
rect 945 3072 1046 3077
rect 1113 3077 1118 3082
rect 1257 3077 1366 3082
rect 1745 3077 1750 3082
rect 1793 3082 1934 3087
rect 2049 3082 2078 3087
rect 1793 3077 1798 3082
rect 1113 3072 1262 3077
rect 1417 3072 1550 3077
rect 1745 3072 1798 3077
rect 1929 3077 1934 3082
rect 2121 3077 2230 3082
rect 2273 3077 2390 3082
rect 2489 3077 2494 3092
rect 2817 3077 2822 3092
rect 3921 3087 3926 3102
rect 4073 3102 4166 3107
rect 4073 3087 4078 3102
rect 4161 3097 4166 3102
rect 4249 3102 4278 3107
rect 4529 3102 4582 3107
rect 4249 3097 4254 3102
rect 4097 3092 4142 3097
rect 4161 3092 4254 3097
rect 4545 3092 4574 3097
rect 1929 3072 2126 3077
rect 2225 3072 2278 3077
rect 2385 3072 2414 3077
rect 2489 3072 2822 3077
rect 3233 3082 3390 3087
rect 3409 3082 3518 3087
rect 3873 3082 3902 3087
rect 3921 3082 4078 3087
rect 4649 3082 4790 3087
rect 769 3067 774 3072
rect 857 3067 950 3072
rect 1417 3067 1422 3072
rect 769 3062 862 3067
rect 969 3062 1102 3067
rect 1097 3057 1102 3062
rect 1273 3062 1302 3067
rect 1393 3062 1422 3067
rect 1545 3067 1550 3072
rect 1593 3067 1710 3072
rect 3233 3067 3238 3082
rect 1545 3062 1598 3067
rect 1705 3062 1734 3067
rect 1809 3062 1918 3067
rect 2137 3062 2318 3067
rect 2353 3062 2414 3067
rect 2977 3062 3238 3067
rect 3385 3067 3390 3082
rect 3385 3062 3854 3067
rect 4049 3062 4646 3067
rect 1273 3057 1278 3062
rect 1729 3057 1814 3062
rect 1913 3057 2142 3062
rect 4641 3057 4646 3062
rect 4801 3062 4870 3067
rect 4801 3057 4806 3062
rect 217 3052 382 3057
rect 1001 3052 1078 3057
rect 1097 3052 1278 3057
rect 1329 3052 1622 3057
rect 1665 3052 1694 3057
rect 2161 3052 2470 3057
rect 2665 3052 2774 3057
rect 3249 3052 3382 3057
rect 3753 3052 3782 3057
rect 4641 3052 4806 3057
rect 217 3037 222 3052
rect 177 3032 222 3037
rect 377 3037 382 3052
rect 2665 3047 2670 3052
rect 729 3042 830 3047
rect 929 3042 1054 3047
rect 1313 3042 1750 3047
rect 1769 3042 1846 3047
rect 1769 3037 1774 3042
rect 377 3032 406 3037
rect 993 3032 1550 3037
rect 1745 3032 1774 3037
rect 1841 3037 1846 3042
rect 1881 3042 2142 3047
rect 2321 3042 2422 3047
rect 2489 3042 2622 3047
rect 2641 3042 2670 3047
rect 2769 3047 2774 3052
rect 2769 3042 2862 3047
rect 3417 3042 3486 3047
rect 4481 3042 4526 3047
rect 1881 3037 1886 3042
rect 2137 3037 2302 3042
rect 2489 3037 2494 3042
rect 1841 3032 1886 3037
rect 2297 3032 2494 3037
rect 2617 3037 2622 3042
rect 3417 3037 3422 3042
rect 2617 3032 2766 3037
rect 2873 3032 3342 3037
rect 3369 3032 3422 3037
rect 3481 3037 3486 3042
rect 4521 3037 4526 3042
rect 4593 3042 4622 3047
rect 4593 3037 4598 3042
rect 3481 3032 3950 3037
rect 4193 3032 4222 3037
rect 4521 3032 4598 3037
rect 1545 3027 1750 3032
rect 2761 3027 2878 3032
rect 233 3022 294 3027
rect 409 3022 462 3027
rect 513 3022 582 3027
rect 633 3022 678 3027
rect 897 3022 966 3027
rect 1153 3022 1182 3027
rect 1377 3022 1406 3027
rect 1497 3022 1526 3027
rect 1777 3022 1830 3027
rect 1897 3022 1950 3027
rect 1985 3022 2622 3027
rect 2697 3022 2742 3027
rect 3433 3022 3478 3027
rect 3489 3022 3558 3027
rect 4105 3022 4230 3027
rect 4337 3022 4398 3027
rect 4673 3022 4734 3027
rect 1401 3017 1502 3022
rect 193 3012 254 3017
rect 697 3012 878 3017
rect 1521 3012 1782 3017
rect 2081 3012 2830 3017
rect 3217 3012 3342 3017
rect 3641 3012 3982 3017
rect 4073 3012 4214 3017
rect 4225 3012 4270 3017
rect 4369 3012 4502 3017
rect 697 3007 702 3012
rect 873 3007 966 3012
rect 1145 3007 1214 3012
rect 1521 3007 1526 3012
rect 121 3002 222 3007
rect 281 3002 702 3007
rect 961 3002 1150 3007
rect 1209 3002 1526 3007
rect 1785 3002 2062 3007
rect 2089 3002 2174 3007
rect 2217 3002 2382 3007
rect 2393 3002 2422 3007
rect 2897 3002 3198 3007
rect 3473 3002 3526 3007
rect 3937 3002 4150 3007
rect 2441 2997 2542 3002
rect 2633 2997 2750 3002
rect 897 2992 950 2997
rect 1161 2992 1198 2997
rect 1561 2992 1670 2997
rect 2065 2992 2446 2997
rect 2537 2992 2638 2997
rect 2745 2992 2878 2997
rect 625 2987 774 2992
rect 2897 2987 2902 3002
rect 3193 2987 3198 3002
rect 4145 2997 4150 3002
rect 3289 2992 3366 2997
rect 3489 2992 3542 2997
rect 3657 2992 3742 2997
rect 3785 2992 3838 2997
rect 4017 2992 4126 2997
rect 4145 2992 4166 2997
rect 4193 2992 4294 2997
rect 4329 2992 4390 2997
rect 4465 2992 4502 2997
rect 4681 2992 4710 2997
rect 273 2982 630 2987
rect 769 2982 1030 2987
rect 1121 2982 1166 2987
rect 1297 2982 1518 2987
rect 1721 2982 1790 2987
rect 1969 2982 2078 2987
rect 2137 2982 2198 2987
rect 2305 2982 2358 2987
rect 2457 2982 2526 2987
rect 2649 2982 2734 2987
rect 2841 2982 2902 2987
rect 2921 2982 3078 2987
rect 3193 2982 3742 2987
rect 1537 2977 1638 2982
rect 2353 2977 2462 2982
rect 2921 2977 2926 2982
rect 641 2972 758 2977
rect 897 2972 918 2977
rect 1153 2972 1206 2977
rect 1313 2972 1350 2977
rect 233 2967 310 2972
rect 1313 2967 1318 2972
rect 209 2962 238 2967
rect 305 2962 486 2967
rect 545 2962 670 2967
rect 729 2962 806 2967
rect 817 2962 1318 2967
rect 1345 2967 1350 2972
rect 1513 2972 1542 2977
rect 1633 2972 1710 2977
rect 1801 2972 1990 2977
rect 2313 2972 2334 2977
rect 2729 2972 2926 2977
rect 3073 2977 3078 2982
rect 3737 2977 3742 2982
rect 3833 2982 4006 2987
rect 4249 2982 4286 2987
rect 4329 2982 4462 2987
rect 3833 2977 3838 2982
rect 3073 2972 3182 2977
rect 3273 2972 3334 2977
rect 3497 2972 3718 2977
rect 3737 2972 3838 2977
rect 3857 2972 3886 2977
rect 4017 2972 4462 2977
rect 1513 2967 1518 2972
rect 1705 2967 1806 2972
rect 3177 2967 3182 2972
rect 3881 2967 4022 2972
rect 1345 2962 1518 2967
rect 1537 2962 1622 2967
rect 1961 2962 2166 2967
rect 2177 2962 2270 2967
rect 2297 2962 2326 2967
rect 2353 2962 2470 2967
rect 2601 2962 2822 2967
rect 2897 2962 3062 2967
rect 3177 2962 3374 2967
rect 2353 2957 2358 2962
rect 265 2952 294 2957
rect 921 2952 950 2957
rect 1217 2952 1326 2957
rect 1577 2952 1950 2957
rect 2113 2952 2230 2957
rect 289 2947 294 2952
rect 625 2947 926 2952
rect 1945 2947 2118 2952
rect 2225 2947 2230 2952
rect 2337 2952 2358 2957
rect 2465 2957 2470 2962
rect 4305 2957 4382 2962
rect 2465 2952 2590 2957
rect 2689 2952 2918 2957
rect 2337 2947 2342 2952
rect 2585 2947 2694 2952
rect 2913 2947 2918 2952
rect 3017 2952 3046 2957
rect 3457 2952 4310 2957
rect 4377 2952 4406 2957
rect 3017 2947 3022 2952
rect 161 2942 222 2947
rect 289 2942 630 2947
rect 1361 2942 1422 2947
rect 2137 2942 2166 2947
rect 2225 2942 2342 2947
rect 2369 2942 2454 2947
rect 2713 2942 2870 2947
rect 2913 2942 3022 2947
rect 3057 2942 3174 2947
rect 3257 2942 3326 2947
rect 4321 2942 4358 2947
rect 4449 2942 4670 2947
rect 649 2932 1350 2937
rect 1433 2932 2206 2937
rect 2433 2932 2478 2937
rect 2569 2932 2614 2937
rect 3049 2932 3086 2937
rect 3185 2932 3302 2937
rect 3961 2932 4022 2937
rect 4065 2932 4118 2937
rect 4369 2932 4406 2937
rect 1345 2927 1438 2932
rect 3081 2927 3190 2932
rect 521 2922 566 2927
rect 2225 2922 2350 2927
rect 2369 2922 2406 2927
rect 2585 2922 2630 2927
rect 2649 2922 2774 2927
rect 2889 2922 2934 2927
rect 3033 2922 3062 2927
rect 3281 2922 3950 2927
rect 4137 2922 4166 2927
rect 4249 2922 4342 2927
rect 4401 2922 4406 2932
rect 4433 2922 4470 2927
rect 1841 2917 1966 2922
rect 2137 2917 2230 2922
rect 2345 2917 2350 2922
rect 2649 2917 2654 2922
rect 97 2912 206 2917
rect 361 2912 406 2917
rect 601 2912 646 2917
rect 697 2912 726 2917
rect 721 2907 726 2912
rect 849 2912 878 2917
rect 913 2912 950 2917
rect 1193 2912 1230 2917
rect 1257 2912 1350 2917
rect 1465 2912 1582 2917
rect 1641 2912 1670 2917
rect 849 2907 854 2912
rect 1665 2907 1670 2912
rect 1817 2912 1846 2917
rect 1961 2912 2142 2917
rect 2345 2912 2366 2917
rect 1817 2907 1822 2912
rect 2361 2907 2366 2912
rect 2489 2912 2654 2917
rect 2769 2917 2774 2922
rect 3281 2917 3286 2922
rect 3945 2917 4142 2922
rect 4161 2917 4166 2922
rect 2769 2912 3022 2917
rect 2489 2907 2494 2912
rect 3017 2907 3022 2912
rect 3081 2912 3286 2917
rect 4161 2912 4286 2917
rect 3081 2907 3086 2912
rect 4281 2907 4286 2912
rect 4369 2912 4422 2917
rect 4369 2907 4374 2912
rect 209 2902 246 2907
rect 393 2902 510 2907
rect 505 2897 510 2902
rect 569 2902 598 2907
rect 721 2902 854 2907
rect 873 2902 990 2907
rect 1009 2902 1134 2907
rect 1153 2902 1206 2907
rect 1457 2902 1534 2907
rect 1665 2902 1822 2907
rect 1841 2902 1950 2907
rect 2153 2902 2334 2907
rect 2361 2902 2494 2907
rect 2609 2902 2694 2907
rect 2729 2902 2758 2907
rect 569 2897 574 2902
rect 1009 2897 1014 2902
rect 505 2892 574 2897
rect 953 2892 1014 2897
rect 1129 2897 1134 2902
rect 1129 2892 1278 2897
rect 1873 2892 1990 2897
rect 2201 2892 2238 2897
rect 2081 2887 2158 2892
rect 2753 2887 2758 2902
rect 2921 2902 2950 2907
rect 3017 2902 3086 2907
rect 3305 2902 3518 2907
rect 3537 2902 3606 2907
rect 3921 2902 4262 2907
rect 4281 2902 4374 2907
rect 4417 2907 4422 2912
rect 4481 2912 4614 2917
rect 4481 2907 4486 2912
rect 4417 2902 4486 2907
rect 2921 2887 2926 2902
rect 3201 2897 3310 2902
rect 3513 2897 3518 2902
rect 3177 2892 3206 2897
rect 3513 2892 3902 2897
rect 3329 2887 3494 2892
rect 4177 2887 4254 2892
rect 233 2882 302 2887
rect 897 2882 1254 2887
rect 1289 2882 1390 2887
rect 1985 2882 2086 2887
rect 2153 2882 2182 2887
rect 2233 2882 2302 2887
rect 2753 2882 2926 2887
rect 3105 2882 3334 2887
rect 3489 2882 3654 2887
rect 3977 2882 4182 2887
rect 4249 2882 4326 2887
rect 4553 2882 4590 2887
rect 1817 2877 1934 2882
rect 801 2872 1014 2877
rect 1137 2872 1262 2877
rect 1401 2872 1822 2877
rect 1929 2872 1958 2877
rect 2097 2872 2150 2877
rect 2321 2872 2414 2877
rect 1257 2867 1406 2872
rect 1977 2867 2078 2872
rect 2169 2867 2326 2872
rect 2409 2867 2414 2872
rect 2457 2872 2598 2877
rect 3041 2872 3422 2877
rect 3473 2872 3502 2877
rect 3601 2872 3750 2877
rect 4193 2872 4238 2877
rect 2457 2867 2462 2872
rect 513 2862 782 2867
rect 825 2862 1198 2867
rect 1209 2862 1238 2867
rect 1833 2862 1982 2867
rect 2073 2862 2174 2867
rect 2409 2862 2462 2867
rect 2593 2867 2598 2872
rect 3497 2867 3606 2872
rect 4057 2867 4174 2872
rect 2593 2862 2622 2867
rect 2961 2862 3198 2867
rect 3761 2862 4062 2867
rect 4169 2862 4294 2867
rect 4441 2862 4558 2867
rect 513 2857 518 2862
rect 489 2852 518 2857
rect 777 2857 782 2862
rect 3193 2857 3326 2862
rect 3761 2857 3766 2862
rect 777 2852 1230 2857
rect 1257 2852 1814 2857
rect 1953 2852 2566 2857
rect 3145 2852 3174 2857
rect 3321 2852 3766 2857
rect 4073 2852 4206 2857
rect 1257 2847 1262 2852
rect 1809 2847 1878 2852
rect 2905 2847 2974 2852
rect 3025 2847 3126 2852
rect 3953 2847 4054 2852
rect 601 2842 758 2847
rect 1033 2842 1086 2847
rect 1169 2842 1262 2847
rect 1873 2842 2110 2847
rect 2577 2842 2910 2847
rect 2969 2842 3030 2847
rect 3121 2842 3302 2847
rect 3929 2842 3958 2847
rect 4049 2842 4134 2847
rect 4401 2842 4454 2847
rect 601 2837 606 2842
rect 753 2837 1014 2842
rect 1081 2837 1174 2842
rect 1465 2837 1622 2842
rect 2105 2837 2518 2842
rect 2577 2837 2582 2842
rect 297 2832 606 2837
rect 1009 2832 1062 2837
rect 1193 2832 1398 2837
rect 1441 2832 1470 2837
rect 1617 2832 1646 2837
rect 1681 2832 1862 2837
rect 1961 2832 2086 2837
rect 2513 2832 2582 2837
rect 2921 2832 2958 2837
rect 3041 2832 3358 2837
rect 3465 2832 3486 2837
rect 3529 2832 3606 2837
rect 3817 2832 4126 2837
rect 4177 2832 4278 2837
rect 4377 2832 4406 2837
rect 1441 2827 1446 2832
rect 153 2822 198 2827
rect 617 2822 710 2827
rect 817 2822 1446 2827
rect 1457 2822 1670 2827
rect 1745 2822 1806 2827
rect 1977 2822 2070 2827
rect 2105 2822 2430 2827
rect 2449 2822 2494 2827
rect 2673 2822 2702 2827
rect 3073 2822 3262 2827
rect 3345 2822 3454 2827
rect 3481 2822 3558 2827
rect 3625 2822 3742 2827
rect 3761 2822 3798 2827
rect 4017 2822 4222 2827
rect 4241 2822 4270 2827
rect 4657 2822 4710 2827
rect 721 2817 822 2822
rect 1849 2817 1958 2822
rect 2105 2817 2110 2822
rect 337 2812 422 2817
rect 489 2812 726 2817
rect 1009 2812 1038 2817
rect 1249 2812 1342 2817
rect 1361 2812 1470 2817
rect 1673 2812 1854 2817
rect 1953 2812 2110 2817
rect 2425 2817 2430 2822
rect 3625 2817 3630 2822
rect 2425 2812 3102 2817
rect 3265 2812 3286 2817
rect 3297 2812 3630 2817
rect 3737 2817 3742 2822
rect 3793 2817 3950 2822
rect 4017 2817 4022 2822
rect 3737 2812 3774 2817
rect 3945 2812 4022 2817
rect 4089 2812 4270 2817
rect 4633 2812 4662 2817
rect 337 2807 342 2812
rect 265 2802 342 2807
rect 417 2807 422 2812
rect 1033 2807 1134 2812
rect 1249 2807 1254 2812
rect 1361 2807 1366 2812
rect 3097 2807 3182 2812
rect 3265 2807 3270 2812
rect 417 2802 446 2807
rect 593 2802 622 2807
rect 809 2802 934 2807
rect 1129 2802 1254 2807
rect 1289 2802 1366 2807
rect 1489 2802 1614 2807
rect 1641 2802 2558 2807
rect 2713 2802 2742 2807
rect 2857 2802 2918 2807
rect 2961 2802 3078 2807
rect 3177 2802 3270 2807
rect 3281 2807 3286 2812
rect 3281 2802 3390 2807
rect 2609 2797 2694 2802
rect 3385 2797 3390 2802
rect 3481 2802 3926 2807
rect 4129 2802 4614 2807
rect 3481 2797 3486 2802
rect 153 2792 286 2797
rect 353 2792 470 2797
rect 625 2792 798 2797
rect 817 2792 886 2797
rect 937 2792 1046 2797
rect 1273 2792 1302 2797
rect 1297 2787 1302 2792
rect 1377 2792 1486 2797
rect 1529 2792 1558 2797
rect 1377 2787 1382 2792
rect 1553 2787 1558 2792
rect 1745 2792 2502 2797
rect 2569 2792 2614 2797
rect 2689 2792 2846 2797
rect 3065 2792 3158 2797
rect 3385 2792 3486 2797
rect 3577 2792 3606 2797
rect 3705 2792 3734 2797
rect 4073 2792 4102 2797
rect 4305 2792 4334 2797
rect 4681 2792 4710 2797
rect 1745 2787 1750 2792
rect 2497 2787 2574 2792
rect 2841 2787 2934 2792
rect 3177 2787 3294 2792
rect 3601 2787 3710 2792
rect 4097 2787 4310 2792
rect 577 2782 886 2787
rect 881 2777 886 2782
rect 1057 2782 1110 2787
rect 1297 2782 1382 2787
rect 1465 2782 1510 2787
rect 1553 2782 1750 2787
rect 1769 2782 2102 2787
rect 2169 2782 2350 2787
rect 2625 2782 2814 2787
rect 2929 2782 3182 2787
rect 3289 2782 3366 2787
rect 3505 2782 3542 2787
rect 3825 2782 4038 2787
rect 1057 2777 1062 2782
rect 2369 2777 2478 2782
rect 3825 2777 3830 2782
rect 881 2772 1062 2777
rect 2081 2772 2374 2777
rect 2473 2772 2686 2777
rect 2825 2772 2910 2777
rect 3193 2772 3278 2777
rect 3385 2772 3486 2777
rect 3505 2772 3670 2777
rect 3689 2772 3782 2777
rect 3801 2772 3830 2777
rect 4033 2777 4038 2782
rect 4033 2772 4246 2777
rect 4449 2772 4478 2777
rect 4689 2772 4718 2777
rect 2681 2767 2830 2772
rect 3385 2767 3390 2772
rect 345 2762 862 2767
rect 857 2757 862 2762
rect 1105 2762 2054 2767
rect 2097 2762 2198 2767
rect 2313 2762 2342 2767
rect 2401 2762 2462 2767
rect 2945 2762 3390 2767
rect 3481 2767 3486 2772
rect 3689 2767 3694 2772
rect 3481 2762 3694 2767
rect 3777 2767 3782 2772
rect 3777 2762 4022 2767
rect 4097 2762 4334 2767
rect 1105 2757 1110 2762
rect 2585 2757 2662 2762
rect 4017 2757 4102 2762
rect 857 2752 1110 2757
rect 2385 2752 2414 2757
rect 2473 2752 2590 2757
rect 2657 2752 2806 2757
rect 2825 2752 2870 2757
rect 3241 2752 3270 2757
rect 3417 2752 3814 2757
rect 3833 2752 3926 2757
rect 4121 2752 4198 2757
rect 657 2747 750 2752
rect 1729 2747 1934 2752
rect 2409 2747 2478 2752
rect 3809 2747 3814 2752
rect 81 2742 286 2747
rect 513 2742 662 2747
rect 745 2742 774 2747
rect 1129 2742 1158 2747
rect 1577 2742 1654 2747
rect 1705 2742 1734 2747
rect 1929 2742 2382 2747
rect 2601 2742 2646 2747
rect 769 2737 774 2742
rect 2641 2737 2646 2742
rect 2745 2742 2862 2747
rect 2953 2742 3014 2747
rect 3057 2742 3214 2747
rect 3305 2742 3502 2747
rect 3809 2742 4110 2747
rect 2745 2737 2750 2742
rect 3521 2737 3662 2742
rect 4105 2737 4110 2742
rect 4193 2742 4222 2747
rect 4657 2742 4734 2747
rect 4193 2737 4198 2742
rect 265 2732 310 2737
rect 465 2732 526 2737
rect 673 2732 710 2737
rect 769 2732 838 2737
rect 1153 2732 1214 2737
rect 1225 2732 1654 2737
rect 1745 2732 1814 2737
rect 1841 2732 1918 2737
rect 2361 2732 2486 2737
rect 2641 2732 2750 2737
rect 2913 2732 2998 2737
rect 3225 2732 3294 2737
rect 3457 2732 3526 2737
rect 3657 2732 3862 2737
rect 465 2727 470 2732
rect 1649 2727 1750 2732
rect 2913 2727 2918 2732
rect 2993 2727 3230 2732
rect 3289 2727 3462 2732
rect 3857 2727 3862 2732
rect 3953 2732 3982 2737
rect 4105 2732 4198 2737
rect 4305 2732 4390 2737
rect 3953 2727 3958 2732
rect 329 2722 470 2727
rect 1025 2722 1110 2727
rect 1937 2722 2182 2727
rect 1025 2717 1030 2722
rect 145 2712 190 2717
rect 249 2712 318 2717
rect 313 2707 318 2712
rect 385 2712 494 2717
rect 505 2712 1030 2717
rect 1105 2717 1110 2722
rect 1417 2717 1486 2722
rect 1937 2717 1942 2722
rect 1105 2712 1422 2717
rect 1481 2712 1686 2717
rect 1713 2712 1942 2717
rect 2177 2717 2182 2722
rect 2249 2722 2342 2727
rect 2601 2722 2622 2727
rect 2833 2722 2918 2727
rect 2929 2722 2974 2727
rect 3481 2722 3646 2727
rect 2249 2717 2254 2722
rect 2337 2717 2470 2722
rect 3641 2717 3646 2722
rect 3809 2722 3838 2727
rect 3857 2722 3958 2727
rect 3809 2717 3814 2722
rect 2177 2712 2254 2717
rect 2465 2712 2894 2717
rect 3073 2712 3158 2717
rect 3217 2712 3518 2717
rect 3585 2712 3622 2717
rect 3641 2712 3814 2717
rect 4017 2712 4086 2717
rect 4177 2712 4238 2717
rect 4361 2712 4430 2717
rect 4449 2712 4518 2717
rect 4577 2712 4774 2717
rect 385 2707 390 2712
rect 4017 2707 4022 2712
rect 177 2702 278 2707
rect 313 2702 390 2707
rect 497 2702 534 2707
rect 1433 2702 1470 2707
rect 1905 2702 2166 2707
rect 2265 2702 2454 2707
rect 2921 2702 2974 2707
rect 3073 2702 3110 2707
rect 3985 2702 4022 2707
rect 4081 2707 4086 2712
rect 4449 2707 4454 2712
rect 4081 2702 4454 2707
rect 4513 2707 4518 2712
rect 4513 2702 4542 2707
rect 169 2692 254 2697
rect 273 2687 278 2702
rect 497 2687 502 2702
rect 1065 2697 1350 2702
rect 1489 2697 1574 2702
rect 2673 2697 2902 2702
rect 3129 2697 3662 2702
rect 521 2692 566 2697
rect 737 2692 1022 2697
rect 1041 2692 1070 2697
rect 1345 2692 1494 2697
rect 1569 2692 2678 2697
rect 2897 2692 3134 2697
rect 3657 2692 3750 2697
rect 3785 2692 3934 2697
rect 4033 2692 4070 2697
rect 4177 2692 4206 2697
rect 737 2687 742 2692
rect 273 2682 502 2687
rect 593 2682 694 2687
rect 713 2682 742 2687
rect 1017 2687 1022 2692
rect 4201 2687 4206 2692
rect 4289 2692 4318 2697
rect 4433 2692 4478 2697
rect 4513 2692 4574 2697
rect 4289 2687 4294 2692
rect 1017 2682 1046 2687
rect 1073 2682 1334 2687
rect 1457 2682 1558 2687
rect 1849 2682 1902 2687
rect 2689 2682 2718 2687
rect 2761 2682 3350 2687
rect 3393 2682 3438 2687
rect 3489 2682 3646 2687
rect 4201 2682 4294 2687
rect 593 2677 598 2682
rect 569 2672 598 2677
rect 689 2677 694 2682
rect 1945 2677 2502 2682
rect 689 2672 1022 2677
rect 1153 2672 1254 2677
rect 1337 2672 1366 2677
rect 1433 2672 1566 2677
rect 1729 2672 1830 2677
rect 1921 2672 1950 2677
rect 2497 2672 2526 2677
rect 2537 2672 2678 2677
rect 2961 2672 3414 2677
rect 3481 2672 3542 2677
rect 3553 2672 3646 2677
rect 3689 2672 3766 2677
rect 1041 2667 1134 2672
rect 1249 2667 1342 2672
rect 1729 2667 1734 2672
rect 561 2662 678 2667
rect 961 2662 1046 2667
rect 1129 2662 1230 2667
rect 1617 2662 1734 2667
rect 1825 2667 1830 2672
rect 2673 2667 2966 2672
rect 1825 2662 2558 2667
rect 2985 2662 3126 2667
rect 3185 2662 3254 2667
rect 3377 2662 3478 2667
rect 3521 2662 3774 2667
rect 3793 2662 4054 2667
rect 673 2657 966 2662
rect 3793 2657 3798 2662
rect 281 2652 430 2657
rect 985 2652 1430 2657
rect 1449 2652 1478 2657
rect 1745 2652 1926 2657
rect 2137 2652 2390 2657
rect 2489 2652 2782 2657
rect 2873 2652 3550 2657
rect 3697 2652 3798 2657
rect 4049 2657 4054 2662
rect 4505 2662 4598 2667
rect 4505 2657 4510 2662
rect 4049 2652 4078 2657
rect 4217 2652 4510 2657
rect 4593 2657 4598 2662
rect 4593 2652 4622 2657
rect 281 2647 286 2652
rect 257 2642 286 2647
rect 425 2647 430 2652
rect 1425 2647 1430 2652
rect 1945 2647 2118 2652
rect 2385 2647 2494 2652
rect 3545 2647 3702 2652
rect 3817 2647 3990 2652
rect 425 2642 1262 2647
rect 1425 2642 1574 2647
rect 1809 2642 1950 2647
rect 2113 2642 2270 2647
rect 3033 2642 3086 2647
rect 3441 2642 3526 2647
rect 3721 2642 3822 2647
rect 3985 2642 4110 2647
rect 2297 2637 2366 2642
rect 2513 2637 3014 2642
rect 3105 2637 3286 2642
rect 161 2632 198 2637
rect 225 2632 294 2637
rect 441 2632 502 2637
rect 921 2632 1110 2637
rect 1233 2632 2302 2637
rect 2361 2632 2518 2637
rect 3009 2632 3110 2637
rect 3281 2632 3974 2637
rect 4057 2632 4086 2637
rect 4137 2632 4206 2637
rect 4521 2632 4614 2637
rect 1105 2627 1238 2632
rect 3969 2627 4062 2632
rect 129 2622 174 2627
rect 281 2622 438 2627
rect 457 2622 494 2627
rect 1257 2622 1286 2627
rect 1369 2622 1590 2627
rect 433 2617 438 2622
rect 849 2617 974 2622
rect 1017 2617 1086 2622
rect 1281 2617 1374 2622
rect 193 2612 302 2617
rect 361 2612 398 2617
rect 433 2612 574 2617
rect 673 2612 710 2617
rect 825 2612 854 2617
rect 969 2612 1022 2617
rect 1081 2612 1110 2617
rect 1177 2612 1222 2617
rect 1393 2612 1438 2617
rect 1521 2612 1550 2617
rect 1585 2607 1590 2622
rect 1753 2622 1814 2627
rect 1825 2622 1998 2627
rect 2105 2622 2222 2627
rect 2313 2622 2350 2627
rect 2529 2622 3270 2627
rect 3417 2622 3502 2627
rect 3529 2622 3550 2627
rect 3697 2622 3798 2627
rect 3897 2622 3950 2627
rect 4201 2622 4318 2627
rect 4337 2622 4374 2627
rect 4545 2622 4702 2627
rect 1753 2607 1758 2622
rect 1809 2617 1814 2622
rect 2377 2617 2486 2622
rect 4105 2617 4182 2622
rect 1809 2612 1854 2617
rect 2041 2612 2070 2617
rect 2353 2612 2382 2617
rect 2481 2612 2518 2617
rect 2689 2612 3398 2617
rect 3457 2612 3718 2617
rect 3769 2612 3910 2617
rect 4041 2612 4110 2617
rect 4177 2612 4438 2617
rect 4601 2612 4694 2617
rect 2065 2607 2182 2612
rect 2353 2607 2358 2612
rect 2513 2607 2678 2612
rect 3393 2607 3398 2612
rect 177 2602 230 2607
rect 561 2602 662 2607
rect 657 2597 662 2602
rect 721 2602 958 2607
rect 1033 2602 1070 2607
rect 1305 2602 1462 2607
rect 1585 2602 1758 2607
rect 1833 2602 2038 2607
rect 2177 2602 2358 2607
rect 2377 2602 2470 2607
rect 2673 2602 2838 2607
rect 2889 2602 3302 2607
rect 3345 2602 3374 2607
rect 3393 2602 3422 2607
rect 3505 2602 3574 2607
rect 3857 2602 3934 2607
rect 4121 2602 4806 2607
rect 721 2597 726 2602
rect 3297 2597 3302 2602
rect 209 2592 238 2597
rect 345 2592 502 2597
rect 657 2592 726 2597
rect 857 2592 934 2597
rect 1057 2592 1102 2597
rect 1217 2592 1286 2597
rect 1345 2592 1374 2597
rect 1473 2592 1566 2597
rect 1777 2592 1846 2597
rect 2113 2592 2158 2597
rect 2489 2592 2654 2597
rect 2737 2592 2806 2597
rect 2841 2592 2886 2597
rect 2969 2592 3110 2597
rect 3121 2592 3174 2597
rect 3249 2592 3286 2597
rect 3297 2592 3446 2597
rect 3761 2592 3814 2597
rect 3873 2592 3910 2597
rect 3921 2592 3998 2597
rect 4553 2592 4726 2597
rect 1369 2587 1478 2592
rect 2489 2587 2494 2592
rect 65 2582 166 2587
rect 161 2577 166 2582
rect 233 2582 262 2587
rect 1873 2582 1902 2587
rect 2457 2582 2494 2587
rect 2649 2587 2654 2592
rect 4081 2587 4270 2592
rect 4313 2587 4430 2592
rect 2649 2582 2758 2587
rect 2913 2582 3262 2587
rect 3369 2582 3414 2587
rect 3545 2582 3590 2587
rect 3609 2582 3742 2587
rect 3793 2582 3902 2587
rect 4001 2582 4086 2587
rect 4265 2582 4318 2587
rect 4425 2582 4454 2587
rect 233 2577 238 2582
rect 2513 2577 2630 2582
rect 2777 2577 2894 2582
rect 3257 2577 3374 2582
rect 3609 2577 3614 2582
rect 161 2572 238 2577
rect 305 2572 1838 2577
rect 1849 2572 2278 2577
rect 2361 2572 2518 2577
rect 2625 2572 2782 2577
rect 2889 2572 2910 2577
rect 2993 2572 3110 2577
rect 3393 2572 3614 2577
rect 3737 2577 3742 2582
rect 3737 2572 3806 2577
rect 3849 2572 3990 2577
rect 4097 2572 4254 2577
rect 4329 2572 4430 2577
rect 4537 2572 4614 2577
rect 2905 2567 2998 2572
rect 3105 2567 3238 2572
rect 3393 2567 3398 2572
rect 3985 2567 4102 2572
rect 2441 2562 2622 2567
rect 2785 2562 2878 2567
rect 3233 2562 3398 2567
rect 3785 2562 3822 2567
rect 337 2557 454 2562
rect 593 2557 686 2562
rect 849 2557 950 2562
rect 1113 2557 1334 2562
rect 1977 2557 2150 2562
rect 2617 2557 2790 2562
rect 3017 2557 3086 2562
rect 3441 2557 3742 2562
rect 4305 2557 4438 2562
rect 313 2552 342 2557
rect 449 2552 478 2557
rect 473 2547 478 2552
rect 569 2552 598 2557
rect 681 2552 798 2557
rect 825 2552 854 2557
rect 945 2552 974 2557
rect 1089 2552 1118 2557
rect 1329 2552 1358 2557
rect 1593 2552 1702 2557
rect 1721 2552 1782 2557
rect 1849 2552 1982 2557
rect 2145 2552 2174 2557
rect 2257 2552 2350 2557
rect 2385 2552 2478 2557
rect 2561 2552 2598 2557
rect 2809 2552 3022 2557
rect 3081 2552 3214 2557
rect 3417 2552 3446 2557
rect 3737 2552 3798 2557
rect 3825 2552 4310 2557
rect 4433 2552 4462 2557
rect 569 2547 574 2552
rect 1593 2547 1598 2552
rect 313 2542 334 2547
rect 353 2542 446 2547
rect 473 2542 574 2547
rect 593 2542 670 2547
rect 665 2537 670 2542
rect 753 2542 1478 2547
rect 1489 2542 1534 2547
rect 1569 2542 1598 2547
rect 1697 2547 1702 2552
rect 1697 2542 1886 2547
rect 1993 2542 2142 2547
rect 2241 2542 2302 2547
rect 2329 2542 2470 2547
rect 2617 2542 2782 2547
rect 3033 2542 3070 2547
rect 3281 2542 3726 2547
rect 4321 2542 4398 2547
rect 4681 2542 4718 2547
rect 753 2537 758 2542
rect 1473 2537 1478 2542
rect 1881 2537 1998 2542
rect 2273 2537 2278 2542
rect 2497 2537 2622 2542
rect 2777 2537 2782 2542
rect 3089 2537 3214 2542
rect 217 2532 350 2537
rect 409 2532 454 2537
rect 665 2532 758 2537
rect 777 2532 798 2537
rect 841 2532 902 2537
rect 961 2532 990 2537
rect 1057 2532 1238 2537
rect 1473 2532 1566 2537
rect 1609 2532 1694 2537
rect 2017 2532 2078 2537
rect 2273 2532 2502 2537
rect 2777 2532 2798 2537
rect 1257 2527 1454 2532
rect 1785 2527 1862 2532
rect 2793 2527 2798 2532
rect 2865 2532 3094 2537
rect 3209 2532 3238 2537
rect 3393 2532 3886 2537
rect 4081 2532 4150 2537
rect 4161 2532 4358 2537
rect 4409 2532 4550 2537
rect 4561 2532 4582 2537
rect 4673 2532 4726 2537
rect 2865 2527 2870 2532
rect 1089 2522 1262 2527
rect 1449 2522 1638 2527
rect 1705 2522 1790 2527
rect 1857 2522 2358 2527
rect 2513 2522 2542 2527
rect 2561 2522 2742 2527
rect 2793 2522 2870 2527
rect 2889 2522 2910 2527
rect 3017 2522 3198 2527
rect 3561 2522 3638 2527
rect 3737 2522 3766 2527
rect 3897 2522 4046 2527
rect 1633 2517 1710 2522
rect 2353 2517 2518 2522
rect 3345 2517 3438 2522
rect 3761 2517 3902 2522
rect 313 2512 382 2517
rect 425 2512 454 2517
rect 537 2512 662 2517
rect 777 2512 838 2517
rect 1081 2512 1118 2517
rect 1201 2512 1534 2517
rect 1545 2512 1614 2517
rect 1801 2512 1846 2517
rect 1977 2512 2022 2517
rect 2265 2512 2334 2517
rect 2545 2512 2590 2517
rect 2649 2512 2694 2517
rect 3089 2512 3350 2517
rect 3433 2512 3558 2517
rect 4313 2512 4414 2517
rect 4521 2512 4566 2517
rect 537 2507 542 2512
rect 241 2502 542 2507
rect 657 2507 662 2512
rect 2105 2507 2246 2512
rect 657 2502 822 2507
rect 1017 2502 1070 2507
rect 1441 2502 1854 2507
rect 1953 2502 2062 2507
rect 2081 2502 2110 2507
rect 2241 2502 2390 2507
rect 2417 2502 2446 2507
rect 2889 2502 2926 2507
rect 3057 2502 3158 2507
rect 3249 2502 3278 2507
rect 3361 2502 3454 2507
rect 3649 2502 4350 2507
rect 4393 2502 4438 2507
rect 4577 2502 4582 2532
rect 345 2492 374 2497
rect 369 2477 374 2492
rect 553 2492 646 2497
rect 553 2477 558 2492
rect 1065 2487 1070 2502
rect 1257 2497 1446 2502
rect 1257 2487 1262 2497
rect 1465 2492 1502 2497
rect 1521 2492 1582 2497
rect 1753 2492 2254 2497
rect 2273 2492 2318 2497
rect 2633 2492 2782 2497
rect 3065 2492 3246 2497
rect 4289 2492 4318 2497
rect 1577 2487 1758 2492
rect 2337 2487 2486 2492
rect 2633 2487 2638 2492
rect 673 2482 750 2487
rect 905 2482 1014 2487
rect 1065 2482 1262 2487
rect 1281 2482 1342 2487
rect 1529 2482 1558 2487
rect 2017 2482 2342 2487
rect 2481 2482 2638 2487
rect 2777 2487 2782 2492
rect 2777 2482 3190 2487
rect 673 2477 678 2482
rect 369 2472 558 2477
rect 577 2472 678 2477
rect 745 2477 750 2482
rect 1553 2477 1558 2482
rect 1777 2477 2022 2482
rect 3185 2477 3190 2482
rect 3257 2482 3350 2487
rect 3257 2477 3262 2482
rect 745 2472 862 2477
rect 1553 2472 1782 2477
rect 2041 2472 2470 2477
rect 2649 2472 2766 2477
rect 3049 2472 3086 2477
rect 3121 2472 3166 2477
rect 3185 2472 3262 2477
rect 3345 2477 3350 2482
rect 3465 2482 4238 2487
rect 3465 2477 3470 2482
rect 3345 2472 3470 2477
rect 4313 2477 4318 2492
rect 4449 2492 4534 2497
rect 4585 2492 4670 2497
rect 4449 2477 4454 2492
rect 4313 2472 4454 2477
rect 689 2462 734 2467
rect 1433 2462 1526 2467
rect 1801 2462 2190 2467
rect 2273 2462 2366 2467
rect 3577 2462 3910 2467
rect 2185 2457 2278 2462
rect 3577 2457 3582 2462
rect 153 2452 174 2457
rect 2049 2452 2166 2457
rect 2297 2452 2422 2457
rect 2473 2452 3326 2457
rect 3553 2452 3582 2457
rect 3905 2457 3910 2462
rect 3953 2462 4086 2467
rect 4105 2462 4246 2467
rect 3953 2457 3958 2462
rect 3905 2452 3958 2457
rect 4081 2457 4086 2462
rect 4081 2452 4174 2457
rect 1433 2447 1550 2452
rect 1929 2447 2030 2452
rect 3601 2447 3774 2452
rect 1017 2442 1326 2447
rect 1345 2442 1438 2447
rect 1545 2442 1574 2447
rect 1713 2442 1806 2447
rect 1905 2442 1934 2447
rect 2025 2442 2118 2447
rect 2153 2442 2390 2447
rect 3513 2442 3542 2447
rect 3569 2442 3606 2447
rect 3769 2442 4142 2447
rect 4457 2442 4502 2447
rect 1017 2437 1022 2442
rect 993 2432 1022 2437
rect 1321 2437 1326 2442
rect 2625 2437 2806 2442
rect 2977 2437 3094 2442
rect 1321 2432 2630 2437
rect 2801 2432 2982 2437
rect 3089 2432 3310 2437
rect 3497 2432 3758 2437
rect 3849 2432 3878 2437
rect 3953 2432 3982 2437
rect 4241 2432 4318 2437
rect 3753 2427 3854 2432
rect 4241 2427 4246 2432
rect 161 2422 606 2427
rect 625 2422 798 2427
rect 1057 2422 1126 2427
rect 1297 2422 1366 2427
rect 1441 2422 1510 2427
rect 1545 2422 1598 2427
rect 1945 2422 2398 2427
rect 2641 2422 2718 2427
rect 2745 2422 2790 2427
rect 2993 2422 3078 2427
rect 3161 2422 3182 2427
rect 3449 2422 3526 2427
rect 3601 2422 3734 2427
rect 3921 2422 4150 2427
rect 4217 2422 4246 2427
rect 4313 2427 4318 2432
rect 4313 2422 4342 2427
rect 1057 2417 1062 2422
rect 81 2412 158 2417
rect 825 2412 1062 2417
rect 1121 2417 1126 2422
rect 1689 2417 1918 2422
rect 2553 2417 2622 2422
rect 2865 2417 2974 2422
rect 4497 2417 4502 2442
rect 4529 2422 4622 2427
rect 1121 2412 1278 2417
rect 1369 2412 1510 2417
rect 1665 2412 1694 2417
rect 1913 2412 2558 2417
rect 2617 2412 2686 2417
rect 2801 2412 2870 2417
rect 2969 2412 3094 2417
rect 3201 2412 3350 2417
rect 3369 2412 3398 2417
rect 3713 2412 3782 2417
rect 3889 2412 3982 2417
rect 4161 2412 4366 2417
rect 4497 2412 4526 2417
rect 2681 2407 2806 2412
rect 3201 2407 3206 2412
rect 1073 2402 1110 2407
rect 1233 2402 1422 2407
rect 1457 2402 1510 2407
rect 1673 2402 1902 2407
rect 1969 2402 2150 2407
rect 2169 2402 2214 2407
rect 2313 2402 2350 2407
rect 2569 2402 2662 2407
rect 2881 2402 3206 2407
rect 3345 2407 3350 2412
rect 3345 2402 3446 2407
rect 3465 2402 3558 2407
rect 3593 2402 3662 2407
rect 3889 2402 3894 2412
rect 3977 2407 4166 2412
rect 3921 2402 3958 2407
rect 4217 2402 4270 2407
rect 4641 2402 4726 2407
rect 2145 2397 2150 2402
rect 225 2392 374 2397
rect 433 2392 566 2397
rect 609 2392 646 2397
rect 961 2392 1014 2397
rect 1073 2392 1134 2397
rect 1193 2392 1214 2397
rect 1297 2392 1326 2397
rect 1609 2392 1718 2397
rect 1801 2392 1838 2397
rect 1929 2392 1966 2397
rect 2145 2392 2334 2397
rect 2393 2392 2438 2397
rect 2465 2392 2582 2397
rect 2761 2392 2814 2397
rect 2881 2392 2886 2402
rect 3465 2397 3470 2402
rect 2937 2392 3038 2397
rect 3057 2392 3110 2397
rect 3177 2392 3246 2397
rect 3257 2392 3470 2397
rect 3553 2397 3558 2402
rect 3921 2397 3926 2402
rect 3553 2392 3582 2397
rect 3857 2392 3926 2397
rect 3937 2392 4054 2397
rect 4113 2392 4262 2397
rect 4289 2392 4438 2397
rect 4505 2392 4606 2397
rect 4665 2392 4742 2397
rect 2601 2387 2742 2392
rect 4289 2387 4294 2392
rect 129 2382 182 2387
rect 505 2382 558 2387
rect 393 2377 486 2382
rect 553 2377 558 2382
rect 657 2382 862 2387
rect 1113 2382 1142 2387
rect 1225 2382 1422 2387
rect 657 2377 662 2382
rect 1137 2377 1230 2382
rect 1417 2377 1422 2382
rect 1521 2382 1598 2387
rect 1729 2382 1918 2387
rect 1977 2382 2326 2387
rect 2409 2382 2606 2387
rect 2737 2382 2886 2387
rect 3481 2382 3846 2387
rect 3961 2382 4294 2387
rect 4433 2387 4438 2392
rect 4433 2382 4462 2387
rect 4497 2382 4638 2387
rect 1521 2377 1526 2382
rect 1593 2377 1734 2382
rect 1913 2377 1982 2382
rect 2321 2377 2414 2382
rect 2881 2377 2886 2382
rect 3121 2377 3486 2382
rect 3841 2377 3966 2382
rect 4497 2377 4502 2382
rect 161 2372 398 2377
rect 481 2372 534 2377
rect 553 2372 662 2377
rect 1361 2372 1398 2377
rect 1417 2372 1526 2377
rect 1817 2372 1862 2377
rect 2153 2372 2302 2377
rect 2433 2372 2862 2377
rect 2881 2372 3126 2377
rect 3505 2372 3630 2377
rect 4073 2372 4502 2377
rect 4513 2372 4558 2377
rect 3649 2367 3782 2372
rect 3985 2367 4078 2372
rect 409 2362 486 2367
rect 849 2362 1158 2367
rect 1281 2362 1390 2367
rect 1673 2362 2142 2367
rect 2313 2362 2550 2367
rect 2649 2362 2686 2367
rect 2705 2362 2846 2367
rect 3209 2362 3422 2367
rect 3553 2362 3654 2367
rect 3777 2362 3846 2367
rect 3929 2362 3990 2367
rect 4097 2362 4134 2367
rect 4169 2362 4382 2367
rect 4465 2362 4662 2367
rect 2137 2357 2142 2362
rect 2225 2357 2318 2362
rect 2545 2357 2654 2362
rect 3209 2357 3214 2362
rect 313 2352 454 2357
rect 633 2352 726 2357
rect 1137 2352 1158 2357
rect 2137 2352 2230 2357
rect 2673 2352 3214 2357
rect 3417 2357 3422 2362
rect 4377 2357 4470 2362
rect 3417 2352 3446 2357
rect 3513 2352 3766 2357
rect 3857 2352 4174 2357
rect 4241 2352 4310 2357
rect 4329 2352 4358 2357
rect 1833 2347 1950 2352
rect 2337 2347 2526 2352
rect 2673 2347 2678 2352
rect 3761 2347 3862 2352
rect 4353 2347 4358 2352
rect 4489 2352 4630 2357
rect 4489 2347 4494 2352
rect 217 2342 334 2347
rect 433 2342 494 2347
rect 721 2342 846 2347
rect 881 2342 926 2347
rect 1809 2342 1838 2347
rect 1945 2342 2070 2347
rect 2249 2342 2342 2347
rect 2521 2342 2678 2347
rect 3225 2342 3286 2347
rect 3297 2342 3422 2347
rect 3505 2342 3606 2347
rect 3665 2342 3742 2347
rect 3889 2342 3982 2347
rect 4105 2342 4134 2347
rect 1721 2332 1742 2337
rect 1785 2332 1846 2337
rect 1905 2332 1934 2337
rect 2081 2332 2238 2337
rect 2353 2332 2382 2337
rect 2409 2332 2510 2337
rect 2681 2332 2870 2337
rect 2913 2332 2990 2337
rect 3409 2332 3518 2337
rect 3537 2332 3670 2337
rect 3753 2332 3934 2337
rect 1929 2327 2086 2332
rect 2233 2327 2358 2332
rect 441 2322 502 2327
rect 985 2322 1654 2327
rect 2137 2322 2158 2327
rect 2385 2322 2414 2327
rect 2505 2322 2582 2327
rect 985 2317 990 2322
rect 265 2312 310 2317
rect 377 2312 422 2317
rect 489 2312 518 2317
rect 537 2312 614 2317
rect 753 2312 990 2317
rect 1649 2317 1654 2322
rect 2409 2317 2510 2322
rect 2641 2317 2838 2322
rect 2913 2317 2918 2332
rect 2985 2327 2990 2332
rect 3537 2327 3542 2332
rect 3665 2327 3758 2332
rect 4145 2327 4150 2347
rect 4193 2342 4254 2347
rect 4353 2342 4494 2347
rect 4537 2342 4654 2347
rect 4177 2332 4302 2337
rect 4569 2332 4702 2337
rect 2985 2322 3150 2327
rect 3161 2322 3366 2327
rect 3505 2322 3542 2327
rect 3577 2322 3646 2327
rect 3849 2322 3886 2327
rect 4129 2322 4150 2327
rect 4513 2322 4566 2327
rect 4617 2322 4758 2327
rect 1649 2312 1678 2317
rect 1817 2312 1870 2317
rect 1881 2312 2358 2317
rect 2529 2312 2646 2317
rect 2833 2312 2918 2317
rect 2929 2312 2974 2317
rect 3193 2312 3230 2317
rect 3353 2312 3414 2317
rect 3489 2312 3606 2317
rect 3689 2312 3742 2317
rect 3913 2312 3966 2317
rect 4161 2312 4246 2317
rect 4281 2312 4366 2317
rect 4617 2312 4646 2317
rect 4641 2307 4646 2312
rect 4769 2312 4798 2317
rect 4769 2307 4774 2312
rect 297 2302 462 2307
rect 585 2302 678 2307
rect 689 2302 750 2307
rect 1473 2302 1630 2307
rect 1473 2297 1478 2302
rect 433 2292 598 2297
rect 705 2292 798 2297
rect 1001 2292 1478 2297
rect 1625 2297 1630 2302
rect 1697 2302 1798 2307
rect 2393 2302 2438 2307
rect 2617 2302 2822 2307
rect 2905 2302 2958 2307
rect 3529 2302 3878 2307
rect 4457 2302 4534 2307
rect 4641 2302 4774 2307
rect 1697 2297 1702 2302
rect 1793 2297 1934 2302
rect 2289 2297 2374 2302
rect 1625 2292 1702 2297
rect 1929 2292 2294 2297
rect 2369 2292 2606 2297
rect 2833 2292 2894 2297
rect 2969 2292 3382 2297
rect 3513 2292 3542 2297
rect 3657 2292 3686 2297
rect 4017 2292 4142 2297
rect 2601 2287 2838 2292
rect 2889 2287 2974 2292
rect 3537 2287 3662 2292
rect 4017 2287 4022 2292
rect 201 2282 286 2287
rect 281 2277 286 2282
rect 481 2282 534 2287
rect 481 2277 486 2282
rect 281 2272 486 2277
rect 529 2267 534 2282
rect 657 2282 718 2287
rect 817 2282 990 2287
rect 657 2267 662 2282
rect 985 2277 990 2282
rect 1489 2282 1774 2287
rect 1849 2282 1918 2287
rect 2305 2282 2350 2287
rect 2409 2282 2454 2287
rect 3769 2282 3798 2287
rect 3993 2282 4022 2287
rect 4137 2287 4142 2292
rect 4137 2282 4350 2287
rect 1489 2277 1494 2282
rect 985 2272 1494 2277
rect 1513 2272 1542 2277
rect 1641 2272 1726 2277
rect 1769 2272 2046 2277
rect 2065 2272 2550 2277
rect 2569 2272 3206 2277
rect 3377 2272 3790 2277
rect 1537 2267 1646 2272
rect 2569 2267 2574 2272
rect 529 2262 662 2267
rect 1665 2262 1694 2267
rect 2465 2262 2574 2267
rect 3201 2267 3206 2272
rect 3201 2262 3230 2267
rect 3921 2262 4550 2267
rect 681 2252 1198 2257
rect 681 2247 686 2252
rect 313 2242 406 2247
rect 425 2242 526 2247
rect 657 2242 686 2247
rect 1193 2247 1198 2252
rect 1265 2252 1446 2257
rect 1465 2252 1582 2257
rect 1265 2247 1270 2252
rect 1193 2242 1270 2247
rect 1441 2247 1446 2252
rect 1689 2247 1694 2262
rect 2177 2257 2470 2262
rect 2593 2257 2966 2262
rect 3025 2257 3126 2262
rect 3561 2257 3726 2262
rect 1905 2252 2182 2257
rect 2489 2252 2598 2257
rect 2961 2252 2990 2257
rect 3001 2252 3030 2257
rect 3121 2252 3190 2257
rect 3537 2252 3566 2257
rect 3721 2252 3750 2257
rect 1905 2247 1910 2252
rect 1441 2242 1622 2247
rect 1689 2242 1910 2247
rect 2201 2242 2294 2247
rect 2369 2242 3110 2247
rect 3433 2242 3766 2247
rect 3865 2242 3950 2247
rect 4289 2242 4334 2247
rect 4449 2242 4478 2247
rect 313 2237 318 2242
rect 161 2232 318 2237
rect 401 2237 406 2242
rect 1305 2237 1406 2242
rect 3865 2237 3870 2242
rect 401 2232 502 2237
rect 929 2232 966 2237
rect 1281 2232 1310 2237
rect 1401 2232 1526 2237
rect 1937 2232 2166 2237
rect 2185 2232 2230 2237
rect 2297 2232 2406 2237
rect 2825 2232 2854 2237
rect 3057 2232 3126 2237
rect 3361 2232 3534 2237
rect 3825 2232 3870 2237
rect 3945 2237 3950 2242
rect 3945 2232 3974 2237
rect 4121 2232 4166 2237
rect 1521 2227 1526 2232
rect 2161 2227 2166 2232
rect 2425 2227 2502 2232
rect 2609 2227 2798 2232
rect 2849 2227 3062 2232
rect 3553 2227 3678 2232
rect 129 2222 174 2227
rect 465 2222 542 2227
rect 625 2222 1182 2227
rect 1297 2222 1486 2227
rect 1521 2222 1662 2227
rect 1929 2222 1966 2227
rect 2161 2222 2430 2227
rect 2497 2222 2614 2227
rect 2793 2222 2822 2227
rect 3217 2222 3270 2227
rect 3313 2222 3558 2227
rect 3673 2222 3718 2227
rect 3737 2222 3790 2227
rect 3881 2222 3958 2227
rect 4049 2222 4158 2227
rect 4185 2222 4438 2227
rect 4537 2222 4766 2227
rect 2073 2217 2142 2222
rect 3081 2217 3198 2222
rect 4185 2217 4190 2222
rect 81 2212 110 2217
rect 209 2212 238 2217
rect 329 2212 638 2217
rect 921 2212 998 2217
rect 1121 2212 1270 2217
rect 1457 2212 1926 2217
rect 105 2207 214 2212
rect 1265 2207 1270 2212
rect 1377 2207 1462 2212
rect 1921 2207 1926 2212
rect 2017 2212 2078 2217
rect 2137 2212 2214 2217
rect 2369 2212 2486 2217
rect 2625 2212 3086 2217
rect 3193 2212 4190 2217
rect 4433 2217 4438 2222
rect 4433 2212 4462 2217
rect 4601 2212 4742 2217
rect 2017 2207 2022 2212
rect 2209 2207 2374 2212
rect 2481 2207 2630 2212
rect 417 2202 622 2207
rect 649 2202 758 2207
rect 1265 2202 1382 2207
rect 1481 2202 1598 2207
rect 1921 2202 2022 2207
rect 2089 2202 2190 2207
rect 2393 2202 2462 2207
rect 2649 2202 2814 2207
rect 3097 2202 3422 2207
rect 3473 2202 3638 2207
rect 3657 2202 4558 2207
rect 3633 2197 3638 2202
rect 177 2192 238 2197
rect 481 2192 662 2197
rect 777 2192 902 2197
rect 937 2192 1062 2197
rect 1137 2192 1182 2197
rect 1401 2192 1494 2197
rect 1617 2192 1902 2197
rect 2169 2192 2534 2197
rect 2665 2192 2734 2197
rect 2865 2192 2966 2197
rect 2985 2192 3046 2197
rect 3241 2192 3382 2197
rect 3489 2192 3598 2197
rect 3633 2192 3710 2197
rect 3785 2192 3814 2197
rect 3833 2192 3950 2197
rect 4145 2192 4230 2197
rect 4521 2192 4678 2197
rect 777 2187 782 2192
rect 545 2182 574 2187
rect 569 2177 574 2182
rect 649 2182 782 2187
rect 897 2187 902 2192
rect 1617 2187 1622 2192
rect 897 2182 1014 2187
rect 1441 2182 1622 2187
rect 1897 2187 1902 2192
rect 2553 2187 2646 2192
rect 2865 2187 2870 2192
rect 1897 2182 2078 2187
rect 2217 2182 2254 2187
rect 2441 2182 2470 2187
rect 2529 2182 2558 2187
rect 2641 2182 2830 2187
rect 2841 2182 2870 2187
rect 2961 2187 2966 2192
rect 3065 2187 3222 2192
rect 3969 2187 4126 2192
rect 2961 2182 3070 2187
rect 3217 2182 3446 2187
rect 3737 2182 3974 2187
rect 4121 2182 4278 2187
rect 4377 2182 4622 2187
rect 649 2177 654 2182
rect 217 2172 438 2177
rect 569 2172 654 2177
rect 881 2172 1006 2177
rect 1001 2167 1006 2172
rect 1073 2172 1542 2177
rect 1633 2172 1886 2177
rect 2089 2172 3566 2177
rect 3585 2172 3686 2177
rect 3705 2172 4214 2177
rect 4233 2172 4390 2177
rect 1073 2167 1078 2172
rect 1537 2167 1638 2172
rect 3585 2167 3590 2172
rect 673 2162 718 2167
rect 745 2162 974 2167
rect 1001 2162 1078 2167
rect 1457 2162 1518 2167
rect 1761 2162 1782 2167
rect 2433 2162 2710 2167
rect 2721 2162 2950 2167
rect 3353 2162 3382 2167
rect 3505 2162 3590 2167
rect 3681 2167 3686 2172
rect 4209 2167 4214 2172
rect 3681 2162 3886 2167
rect 4033 2162 4062 2167
rect 4129 2162 4174 2167
rect 4209 2162 4238 2167
rect 4401 2162 4598 2167
rect 2193 2157 2414 2162
rect 2945 2157 3254 2162
rect 3353 2157 3358 2162
rect 3881 2157 4038 2162
rect 4233 2157 4406 2162
rect 393 2152 542 2157
rect 553 2152 582 2157
rect 657 2152 742 2157
rect 849 2152 966 2157
rect 1465 2152 1694 2157
rect 1905 2152 2062 2157
rect 2169 2152 2198 2157
rect 2409 2152 2926 2157
rect 3249 2152 3358 2157
rect 3385 2152 3494 2157
rect 209 2142 342 2147
rect 433 2142 566 2147
rect 697 2142 830 2147
rect 849 2137 854 2152
rect 961 2142 982 2147
rect 1121 2142 1158 2147
rect 1449 2142 1550 2147
rect 1545 2137 1550 2142
rect 1681 2142 1710 2147
rect 1681 2137 1686 2142
rect 1905 2137 1910 2152
rect 169 2132 222 2137
rect 329 2132 526 2137
rect 537 2132 574 2137
rect 609 2132 854 2137
rect 1305 2132 1390 2137
rect 1505 2132 1526 2137
rect 1545 2132 1686 2137
rect 1713 2132 1790 2137
rect 1873 2132 1910 2137
rect 2057 2137 2062 2152
rect 3489 2147 3494 2152
rect 3561 2152 3718 2157
rect 3833 2152 3862 2157
rect 3561 2147 3566 2152
rect 3713 2147 3838 2152
rect 4121 2147 4198 2152
rect 2081 2142 2806 2147
rect 2993 2142 3102 2147
rect 3137 2142 3230 2147
rect 3489 2142 3566 2147
rect 3585 2142 3694 2147
rect 3937 2142 4022 2147
rect 4097 2142 4126 2147
rect 4193 2142 4414 2147
rect 4569 2142 4598 2147
rect 4097 2137 4102 2142
rect 2057 2132 2454 2137
rect 2505 2132 2606 2137
rect 2697 2132 2726 2137
rect 2905 2132 3310 2137
rect 3713 2132 3822 2137
rect 225 2122 318 2127
rect 417 2122 534 2127
rect 545 2122 742 2127
rect 857 2122 1086 2127
rect 313 2117 422 2122
rect 737 2117 838 2122
rect 137 2112 182 2117
rect 193 2112 222 2117
rect 233 2112 286 2117
rect 441 2112 478 2117
rect 665 2112 726 2117
rect 833 2112 902 2117
rect 1153 2112 1254 2117
rect 1489 2112 1510 2117
rect 921 2107 1134 2112
rect 1521 2107 1526 2132
rect 2601 2127 2702 2132
rect 3713 2127 3718 2132
rect 1889 2122 2582 2127
rect 2577 2117 2582 2122
rect 2737 2122 3006 2127
rect 3129 2122 3182 2127
rect 3321 2122 3430 2127
rect 3449 2122 3502 2127
rect 3601 2122 3718 2127
rect 3817 2127 3822 2132
rect 3889 2132 4102 2137
rect 4145 2132 4182 2137
rect 3889 2127 3894 2132
rect 4273 2127 4278 2137
rect 4393 2132 4470 2137
rect 4641 2132 4726 2137
rect 3817 2122 3894 2127
rect 3937 2122 4230 2127
rect 4273 2122 4302 2127
rect 2737 2117 2742 2122
rect 3001 2117 3134 2122
rect 3177 2117 3326 2122
rect 3425 2117 3430 2122
rect 1913 2112 1942 2117
rect 1937 2107 1942 2112
rect 2049 2112 2302 2117
rect 2529 2112 2558 2117
rect 2577 2112 2742 2117
rect 2881 2112 2982 2117
rect 3425 2112 4254 2117
rect 2049 2107 2054 2112
rect 2297 2107 2534 2112
rect 4297 2107 4302 2122
rect 4481 2122 4606 2127
rect 4481 2107 4486 2122
rect 377 2102 614 2107
rect 625 2102 926 2107
rect 1129 2102 1222 2107
rect 1273 2102 1470 2107
rect 1505 2102 1526 2107
rect 1545 2102 1702 2107
rect 1937 2102 2054 2107
rect 2145 2102 2278 2107
rect 3097 2102 3302 2107
rect 3361 2102 3406 2107
rect 3481 2102 3606 2107
rect 3697 2102 3790 2107
rect 1273 2097 1278 2102
rect 201 2092 366 2097
rect 433 2092 486 2097
rect 617 2092 1278 2097
rect 1465 2097 1470 2102
rect 1545 2097 1550 2102
rect 1465 2092 1550 2097
rect 1697 2097 1702 2102
rect 3097 2097 3102 2102
rect 1697 2092 1870 2097
rect 2073 2092 2134 2097
rect 361 2087 438 2092
rect 481 2087 598 2092
rect 2129 2087 2134 2092
rect 2193 2092 3102 2097
rect 3297 2097 3302 2102
rect 3785 2097 3790 2102
rect 3865 2102 3894 2107
rect 3945 2102 4094 2107
rect 4113 2102 4278 2107
rect 4297 2102 4486 2107
rect 3865 2097 3870 2102
rect 3297 2092 3326 2097
rect 3409 2092 3438 2097
rect 3561 2092 3590 2097
rect 3785 2092 3870 2097
rect 3913 2092 3934 2097
rect 2193 2087 2198 2092
rect 3321 2087 3414 2092
rect 593 2082 758 2087
rect 913 2082 1454 2087
rect 1561 2082 1686 2087
rect 2129 2082 2198 2087
rect 2273 2082 2438 2087
rect 2969 2082 2998 2087
rect 3113 2082 3286 2087
rect 777 2077 918 2082
rect 1449 2077 1566 2082
rect 2993 2077 3118 2082
rect 3281 2077 3286 2082
rect 3449 2082 3502 2087
rect 3449 2077 3454 2082
rect 0 2072 782 2077
rect 1009 2072 1038 2077
rect 1081 2072 1270 2077
rect 2217 2072 2366 2077
rect 2457 2072 2558 2077
rect 3281 2072 3454 2077
rect 3585 2077 3590 2092
rect 3913 2077 3918 2092
rect 3929 2087 3934 2092
rect 4057 2092 4086 2097
rect 4057 2087 4062 2092
rect 3929 2082 4062 2087
rect 3585 2072 3918 2077
rect 2457 2067 2462 2072
rect 497 2062 550 2067
rect 601 2062 1630 2067
rect 1737 2062 1830 2067
rect 1921 2062 2126 2067
rect 2425 2062 2462 2067
rect 2553 2067 2558 2072
rect 2553 2062 2582 2067
rect 2617 2062 2662 2067
rect 2777 2062 3262 2067
rect 3937 2062 4110 2067
rect 497 2057 502 2062
rect 1921 2057 1926 2062
rect 249 2052 502 2057
rect 553 2052 662 2057
rect 777 2052 1310 2057
rect 1641 2052 1926 2057
rect 2121 2057 2126 2062
rect 2121 2052 2150 2057
rect 2361 2052 2390 2057
rect 2481 2052 2510 2057
rect 2521 2052 2550 2057
rect 2673 2052 2766 2057
rect 657 2047 782 2052
rect 1305 2047 1502 2052
rect 1641 2047 1646 2052
rect 2385 2047 2486 2052
rect 2545 2047 2678 2052
rect 2761 2047 2766 2052
rect 3225 2052 3414 2057
rect 3225 2047 3230 2052
rect 337 2042 638 2047
rect 801 2042 854 2047
rect 969 2042 1286 2047
rect 1497 2042 1646 2047
rect 1961 2042 2038 2047
rect 1961 2037 1966 2042
rect 169 2032 262 2037
rect 257 2027 262 2032
rect 345 2032 630 2037
rect 745 2032 806 2037
rect 969 2032 1478 2037
rect 1937 2032 1966 2037
rect 2033 2037 2038 2042
rect 2193 2042 2278 2047
rect 2761 2042 3230 2047
rect 3433 2042 3598 2047
rect 2193 2037 2198 2042
rect 2033 2032 2198 2037
rect 2273 2037 2278 2042
rect 3273 2037 3366 2042
rect 3433 2037 3438 2042
rect 2273 2032 2438 2037
rect 2553 2032 2686 2037
rect 3249 2032 3278 2037
rect 3361 2032 3438 2037
rect 3593 2037 3598 2042
rect 3593 2032 3622 2037
rect 345 2027 350 2032
rect 857 2027 950 2032
rect 137 2022 182 2027
rect 201 2022 238 2027
rect 257 2022 350 2027
rect 385 2022 422 2027
rect 521 2022 566 2027
rect 681 2022 750 2027
rect 769 2022 862 2027
rect 945 2022 998 2027
rect 1033 2022 1142 2027
rect 1233 2022 1278 2027
rect 1457 2022 1494 2027
rect 1529 2022 1766 2027
rect 1969 2022 1998 2027
rect 2121 2022 2190 2027
rect 2273 2022 2318 2027
rect 2505 2022 2606 2027
rect 2641 2022 2742 2027
rect 2777 2022 2806 2027
rect 3065 2022 3142 2027
rect 3265 2022 3350 2027
rect 3473 2022 3574 2027
rect 3761 2022 3814 2027
rect 4329 2022 4518 2027
rect 4569 2022 4630 2027
rect 1529 2017 1534 2022
rect 545 2012 614 2017
rect 641 2012 686 2017
rect 721 2012 934 2017
rect 1153 2012 1222 2017
rect 1289 2012 1446 2017
rect 1505 2012 1534 2017
rect 1761 2017 1766 2022
rect 1993 2017 2126 2022
rect 2337 2017 2430 2022
rect 3473 2017 3478 2022
rect 3569 2017 3670 2022
rect 1761 2012 1958 2017
rect 929 2007 1158 2012
rect 1217 2007 1294 2012
rect 1441 2007 1510 2012
rect 1953 2007 1958 2012
rect 2201 2012 2342 2017
rect 2425 2012 3238 2017
rect 3305 2012 3478 2017
rect 3665 2012 3782 2017
rect 2201 2007 2206 2012
rect 3233 2007 3238 2012
rect 369 2002 430 2007
rect 617 2002 910 2007
rect 1953 2002 2206 2007
rect 2265 2002 2374 2007
rect 2385 2002 2414 2007
rect 3097 2002 3158 2007
rect 3233 2002 3326 2007
rect 3489 2002 3654 2007
rect 3921 2002 4006 2007
rect 4457 2002 4502 2007
rect 2369 1997 2374 2002
rect 2433 1997 2550 2002
rect 2617 1997 2758 2002
rect 89 1992 286 1997
rect 417 1992 574 1997
rect 665 1992 1158 1997
rect 1233 1992 1254 1997
rect 1273 1992 1526 1997
rect 1545 1992 1750 1997
rect 2249 1992 2310 1997
rect 2369 1992 2438 1997
rect 2545 1992 2622 1997
rect 2753 1992 2782 1997
rect 3009 1992 3078 1997
rect 3561 1992 3662 1997
rect 4073 1992 4110 1997
rect 4425 1992 4542 1997
rect 4625 1992 4734 1997
rect 1153 1987 1158 1992
rect 1273 1987 1278 1992
rect 305 1982 358 1987
rect 353 1977 358 1982
rect 417 1982 446 1987
rect 545 1982 846 1987
rect 1153 1982 1278 1987
rect 1521 1987 1526 1992
rect 3897 1987 4014 1992
rect 1521 1982 1566 1987
rect 1769 1982 1950 1987
rect 417 1977 422 1982
rect 921 1977 1134 1982
rect 1297 1977 1446 1982
rect 1769 1977 1774 1982
rect 353 1972 422 1977
rect 545 1972 582 1977
rect 681 1972 710 1977
rect 857 1972 926 1977
rect 1129 1972 1302 1977
rect 1441 1972 1774 1977
rect 1945 1977 1950 1982
rect 2049 1982 2190 1987
rect 2209 1982 2534 1987
rect 2633 1982 2718 1987
rect 2793 1982 3422 1987
rect 3585 1982 3718 1987
rect 3833 1982 3902 1987
rect 4009 1982 4102 1987
rect 2049 1977 2054 1982
rect 1945 1972 1974 1977
rect 2025 1972 2054 1977
rect 2185 1977 2190 1982
rect 2529 1977 2638 1982
rect 2713 1977 2798 1982
rect 2185 1972 2510 1977
rect 2657 1972 2694 1977
rect 2945 1972 3142 1977
rect 3641 1972 3678 1977
rect 3713 1972 3822 1977
rect 3913 1972 3942 1977
rect 3969 1972 3998 1977
rect 4113 1972 4430 1977
rect 4449 1972 4558 1977
rect 705 1967 862 1972
rect 1793 1967 1926 1972
rect 3817 1967 3918 1972
rect 3993 1967 4118 1972
rect 4449 1967 4454 1972
rect 937 1962 1798 1967
rect 1921 1962 2174 1967
rect 2521 1962 2646 1967
rect 2705 1962 3206 1967
rect 3369 1962 3566 1967
rect 4393 1962 4454 1967
rect 4553 1967 4558 1972
rect 4553 1962 4606 1967
rect 2169 1957 2462 1962
rect 2521 1957 2526 1962
rect 2641 1957 2710 1962
rect 3369 1957 3374 1962
rect 3561 1957 3734 1962
rect 737 1952 766 1957
rect 761 1947 766 1952
rect 881 1952 958 1957
rect 1057 1952 1166 1957
rect 1257 1952 2078 1957
rect 2457 1952 2526 1957
rect 3001 1952 3078 1957
rect 3185 1952 3374 1957
rect 3729 1952 3902 1957
rect 3913 1952 4150 1957
rect 4361 1952 4646 1957
rect 881 1947 886 1952
rect 953 1947 1046 1952
rect 265 1942 302 1947
rect 329 1942 606 1947
rect 665 1942 686 1947
rect 761 1942 886 1947
rect 905 1942 934 1947
rect 1041 1937 1046 1947
rect 1129 1942 1422 1947
rect 1457 1942 1518 1947
rect 1881 1942 2022 1947
rect 2241 1942 2294 1947
rect 2369 1942 2438 1947
rect 2577 1942 2606 1947
rect 2625 1942 2782 1947
rect 3009 1942 3054 1947
rect 3385 1942 3430 1947
rect 3473 1942 3718 1947
rect 3841 1942 3950 1947
rect 4209 1942 4310 1947
rect 4433 1942 4478 1947
rect 4673 1942 4710 1947
rect 1129 1937 1134 1942
rect 1625 1937 1862 1942
rect 2625 1937 2630 1942
rect 2777 1937 2886 1942
rect 553 1932 646 1937
rect 977 1932 1006 1937
rect 1041 1932 1134 1937
rect 1313 1932 1342 1937
rect 1529 1932 1630 1937
rect 1857 1932 2230 1937
rect 2305 1932 2358 1937
rect 2449 1932 2630 1937
rect 2881 1932 2998 1937
rect 3065 1932 3190 1937
rect 3481 1932 3558 1937
rect 3865 1932 4070 1937
rect 4089 1932 4142 1937
rect 2225 1927 2310 1932
rect 2353 1927 2454 1932
rect 2657 1927 2742 1932
rect 2993 1927 3070 1932
rect 3665 1927 3766 1932
rect 4321 1927 4502 1932
rect 1369 1922 1390 1927
rect 1641 1922 1846 1927
rect 1865 1922 1958 1927
rect 2585 1922 2662 1927
rect 2737 1922 2766 1927
rect 2841 1922 2870 1927
rect 3641 1922 3670 1927
rect 3761 1922 4046 1927
rect 4241 1922 4326 1927
rect 4497 1922 4678 1927
rect 1473 1917 1606 1922
rect 137 1912 182 1917
rect 777 1912 838 1917
rect 1153 1912 1198 1917
rect 1305 1912 1334 1917
rect 1401 1912 1478 1917
rect 1601 1912 2126 1917
rect 2145 1912 2246 1917
rect 2265 1912 2310 1917
rect 2329 1912 2382 1917
rect 2409 1912 2462 1917
rect 2673 1912 2718 1917
rect 2889 1912 3206 1917
rect 3225 1912 3334 1917
rect 3353 1912 3462 1917
rect 3689 1912 3878 1917
rect 3897 1912 3950 1917
rect 4161 1912 4262 1917
rect 4337 1912 4390 1917
rect 4433 1912 4486 1917
rect 4641 1912 4702 1917
rect 1329 1907 1406 1912
rect 2145 1907 2150 1912
rect 169 1902 502 1907
rect 625 1902 1310 1907
rect 1489 1902 1590 1907
rect 2081 1902 2150 1907
rect 2241 1907 2246 1912
rect 2481 1907 2574 1912
rect 2817 1907 2894 1912
rect 3201 1907 3206 1912
rect 3353 1907 3358 1912
rect 2241 1902 2486 1907
rect 2569 1902 2662 1907
rect 1609 1897 1982 1902
rect 2657 1897 2662 1902
rect 2729 1902 2822 1907
rect 3201 1902 3358 1907
rect 3457 1907 3462 1912
rect 3457 1902 3486 1907
rect 3513 1902 3870 1907
rect 4041 1902 4174 1907
rect 4617 1902 4646 1907
rect 2729 1897 2734 1902
rect 3089 1897 3182 1902
rect 4641 1897 4646 1902
rect 4713 1902 4766 1907
rect 4713 1897 4718 1902
rect 825 1892 862 1897
rect 1129 1892 1174 1897
rect 1505 1892 1614 1897
rect 1977 1892 2070 1897
rect 2137 1892 2558 1897
rect 2657 1892 2734 1897
rect 2833 1892 3094 1897
rect 3177 1892 3374 1897
rect 3417 1892 3446 1897
rect 2065 1887 2142 1892
rect 3441 1887 3446 1892
rect 3825 1892 3854 1897
rect 4641 1892 4718 1897
rect 3825 1887 3830 1892
rect 481 1882 574 1887
rect 833 1882 894 1887
rect 1385 1882 1470 1887
rect 1521 1882 1966 1887
rect 2465 1882 2566 1887
rect 3105 1882 3278 1887
rect 3441 1882 3830 1887
rect 1073 1877 1150 1882
rect 1385 1877 1390 1882
rect 729 1872 846 1877
rect 993 1872 1078 1877
rect 1145 1872 1390 1877
rect 1465 1877 1470 1882
rect 2161 1877 2446 1882
rect 1465 1872 1622 1877
rect 1857 1872 2166 1877
rect 2441 1872 3094 1877
rect 3193 1872 3222 1877
rect 3249 1872 3294 1877
rect 1617 1867 1750 1872
rect 1857 1867 1862 1872
rect 3089 1867 3198 1872
rect 1089 1862 1134 1867
rect 1417 1862 1598 1867
rect 1745 1862 1862 1867
rect 1881 1862 1982 1867
rect 1977 1857 1982 1862
rect 2081 1862 2110 1867
rect 2177 1862 2574 1867
rect 2081 1857 2086 1862
rect 2817 1857 2974 1862
rect 161 1852 294 1857
rect 313 1852 470 1857
rect 721 1852 1302 1857
rect 1577 1852 1726 1857
rect 1977 1852 2086 1857
rect 2321 1852 2454 1857
rect 2585 1852 2822 1857
rect 2969 1852 2998 1857
rect 3017 1852 3182 1857
rect 3481 1852 3798 1857
rect 4577 1852 4654 1857
rect 313 1837 318 1852
rect 257 1832 318 1837
rect 465 1837 470 1852
rect 1297 1847 1302 1852
rect 1401 1847 1582 1852
rect 2153 1847 2278 1852
rect 2449 1847 2590 1852
rect 3017 1847 3022 1852
rect 1097 1842 1158 1847
rect 1297 1842 1406 1847
rect 1745 1842 1958 1847
rect 2129 1842 2158 1847
rect 2273 1842 2430 1847
rect 2833 1842 3022 1847
rect 3177 1847 3182 1852
rect 3177 1842 3246 1847
rect 4001 1842 4150 1847
rect 4601 1842 4630 1847
rect 1601 1837 1750 1842
rect 1953 1837 1958 1842
rect 2649 1837 2766 1842
rect 465 1832 494 1837
rect 585 1832 646 1837
rect 833 1832 902 1837
rect 1073 1832 1190 1837
rect 1241 1832 1278 1837
rect 1425 1832 1606 1837
rect 1953 1832 2510 1837
rect 2625 1832 2654 1837
rect 2761 1832 2790 1837
rect 2921 1832 3166 1837
rect 3433 1832 3550 1837
rect 3817 1832 3982 1837
rect 833 1827 838 1832
rect 145 1822 190 1827
rect 329 1822 374 1827
rect 417 1822 478 1827
rect 545 1822 734 1827
rect 745 1822 838 1827
rect 897 1827 902 1832
rect 897 1822 1078 1827
rect 1225 1822 1254 1827
rect 1617 1822 1942 1827
rect 2137 1822 2182 1827
rect 2345 1822 2534 1827
rect 2689 1822 2742 1827
rect 3281 1822 3406 1827
rect 1073 1817 1230 1822
rect 1977 1817 2118 1822
rect 2201 1817 2302 1822
rect 3441 1817 3446 1827
rect 3465 1822 3510 1827
rect 3529 1822 3566 1827
rect 3585 1822 3630 1827
rect 3817 1817 3822 1832
rect 3977 1817 3982 1832
rect 4001 1817 4006 1842
rect 4145 1837 4150 1842
rect 4145 1832 4334 1837
rect 4497 1832 4598 1837
rect 4673 1832 4758 1837
rect 4329 1827 4334 1832
rect 4673 1827 4678 1832
rect 4329 1822 4358 1827
rect 4425 1822 4550 1827
rect 4601 1822 4678 1827
rect 4753 1827 4758 1832
rect 4753 1822 4782 1827
rect 281 1812 430 1817
rect 849 1812 886 1817
rect 1033 1812 1054 1817
rect 1369 1812 1894 1817
rect 625 1807 758 1812
rect 905 1807 1014 1812
rect 1889 1807 1894 1812
rect 1953 1812 1982 1817
rect 2113 1812 2206 1817
rect 2297 1812 2326 1817
rect 2337 1812 2414 1817
rect 3337 1812 3390 1817
rect 3441 1812 3526 1817
rect 3641 1812 3822 1817
rect 3841 1812 3958 1817
rect 3977 1812 4006 1817
rect 4017 1812 4134 1817
rect 4401 1812 4462 1817
rect 4673 1812 4758 1817
rect 1953 1807 1958 1812
rect 3521 1807 3646 1812
rect 3841 1807 3846 1812
rect 81 1802 134 1807
rect 129 1797 134 1802
rect 193 1802 222 1807
rect 233 1802 270 1807
rect 193 1797 198 1802
rect 129 1792 198 1797
rect 265 1797 270 1802
rect 329 1802 630 1807
rect 753 1802 910 1807
rect 1009 1802 1270 1807
rect 1625 1802 1862 1807
rect 1889 1802 1958 1807
rect 2001 1802 2038 1807
rect 2057 1802 2110 1807
rect 2121 1802 2206 1807
rect 2241 1802 2318 1807
rect 2993 1802 3078 1807
rect 3473 1802 3502 1807
rect 3809 1802 3846 1807
rect 3953 1807 3958 1812
rect 3953 1802 3982 1807
rect 4145 1802 4638 1807
rect 4649 1802 4718 1807
rect 329 1797 334 1802
rect 1289 1797 1502 1802
rect 2993 1797 2998 1802
rect 265 1792 334 1797
rect 353 1792 462 1797
rect 641 1792 742 1797
rect 737 1787 742 1792
rect 873 1792 1110 1797
rect 873 1787 878 1792
rect 1105 1787 1110 1792
rect 1201 1792 1294 1797
rect 1497 1792 1526 1797
rect 1697 1792 1726 1797
rect 1841 1792 1870 1797
rect 2065 1792 2230 1797
rect 2409 1792 2454 1797
rect 2473 1792 2566 1797
rect 1201 1787 1206 1792
rect 1953 1787 2046 1792
rect 2249 1787 2390 1792
rect 2473 1787 2478 1792
rect 465 1782 574 1787
rect 737 1782 878 1787
rect 897 1782 926 1787
rect 1057 1782 1086 1787
rect 1105 1782 1206 1787
rect 1257 1782 1646 1787
rect 1705 1782 1734 1787
rect 1841 1782 1918 1787
rect 1929 1782 1958 1787
rect 2041 1782 2254 1787
rect 2385 1782 2478 1787
rect 2561 1787 2566 1792
rect 2689 1792 2774 1797
rect 2793 1792 2878 1797
rect 2969 1792 2998 1797
rect 3073 1797 3078 1802
rect 3977 1797 4150 1802
rect 3073 1792 3102 1797
rect 3121 1792 3238 1797
rect 3505 1792 3542 1797
rect 3609 1792 3646 1797
rect 3849 1792 3950 1797
rect 4393 1792 4414 1797
rect 4569 1792 4670 1797
rect 2689 1787 2694 1792
rect 2561 1782 2694 1787
rect 2769 1787 2774 1792
rect 2769 1782 3182 1787
rect 3249 1782 3486 1787
rect 3897 1782 4182 1787
rect 4281 1782 4558 1787
rect 4617 1782 4694 1787
rect 921 1777 1062 1782
rect 3177 1777 3254 1782
rect 4553 1777 4622 1782
rect 377 1772 486 1777
rect 689 1772 718 1777
rect 1385 1772 2046 1777
rect 2137 1772 2542 1777
rect 2705 1772 2758 1777
rect 2753 1767 2758 1772
rect 2825 1772 2854 1777
rect 3089 1772 3158 1777
rect 4641 1772 4742 1777
rect 2825 1767 2830 1772
rect 97 1762 158 1767
rect 329 1762 646 1767
rect 641 1757 646 1762
rect 737 1762 838 1767
rect 889 1762 1014 1767
rect 1225 1762 2022 1767
rect 2033 1762 2550 1767
rect 2753 1762 2830 1767
rect 2857 1762 2902 1767
rect 3225 1762 3382 1767
rect 4449 1762 4718 1767
rect 737 1757 742 1762
rect 177 1752 390 1757
rect 425 1752 550 1757
rect 641 1752 742 1757
rect 833 1757 838 1762
rect 2017 1757 2022 1762
rect 4449 1757 4454 1762
rect 833 1752 862 1757
rect 937 1752 990 1757
rect 1529 1752 1982 1757
rect 2017 1752 2222 1757
rect 2241 1752 2326 1757
rect 2929 1752 3254 1757
rect 3777 1752 3902 1757
rect 4001 1752 4246 1757
rect 4305 1752 4454 1757
rect 4561 1752 4670 1757
rect 1289 1747 1414 1752
rect 4561 1747 4566 1752
rect 361 1742 454 1747
rect 553 1742 654 1747
rect 769 1742 870 1747
rect 977 1742 1006 1747
rect 1097 1742 1294 1747
rect 1409 1742 1518 1747
rect 1593 1742 1622 1747
rect 1713 1742 1742 1747
rect 1929 1742 2094 1747
rect 2105 1742 2414 1747
rect 2569 1742 2838 1747
rect 2865 1742 2926 1747
rect 2977 1742 3062 1747
rect 1513 1737 1598 1742
rect 1737 1737 1934 1742
rect 2569 1737 2574 1742
rect 441 1732 758 1737
rect 753 1727 758 1732
rect 881 1732 1014 1737
rect 1305 1732 1374 1737
rect 881 1727 886 1732
rect 1393 1727 1398 1737
rect 1953 1732 2006 1737
rect 2169 1732 2222 1737
rect 2313 1732 2342 1737
rect 2025 1727 2150 1732
rect 2337 1727 2342 1732
rect 2409 1732 2574 1737
rect 2833 1737 2838 1742
rect 3057 1737 3062 1742
rect 3129 1742 3262 1747
rect 3313 1742 3342 1747
rect 3369 1742 3462 1747
rect 3593 1742 3702 1747
rect 3825 1742 4062 1747
rect 4385 1742 4566 1747
rect 4585 1742 4614 1747
rect 3129 1737 3134 1742
rect 2833 1732 2886 1737
rect 3057 1732 3134 1737
rect 3377 1732 3398 1737
rect 3665 1732 3814 1737
rect 3977 1732 4006 1737
rect 4081 1732 4206 1737
rect 2409 1727 2414 1732
rect 2681 1727 2790 1732
rect 217 1722 294 1727
rect 329 1722 422 1727
rect 513 1722 606 1727
rect 753 1722 886 1727
rect 1225 1722 1534 1727
rect 1601 1722 1638 1727
rect 1697 1722 1758 1727
rect 1777 1722 1934 1727
rect 217 1717 222 1722
rect 169 1712 222 1717
rect 289 1717 294 1722
rect 1777 1717 1782 1722
rect 289 1712 318 1717
rect 337 1712 446 1717
rect 497 1712 598 1717
rect 1033 1712 1206 1717
rect 1393 1712 1446 1717
rect 1561 1712 1782 1717
rect 1929 1717 1934 1722
rect 2001 1722 2030 1727
rect 2145 1722 2214 1727
rect 2337 1722 2414 1727
rect 2529 1722 2606 1727
rect 2657 1722 2686 1727
rect 2785 1722 2814 1727
rect 3153 1722 3238 1727
rect 2001 1717 2006 1722
rect 3665 1717 3670 1732
rect 3809 1727 3982 1732
rect 4081 1727 4086 1732
rect 3681 1722 3718 1727
rect 4049 1722 4086 1727
rect 4201 1727 4206 1732
rect 4297 1732 4366 1737
rect 4473 1732 4558 1737
rect 4641 1732 4662 1737
rect 4297 1727 4302 1732
rect 4201 1722 4302 1727
rect 4361 1727 4366 1732
rect 4361 1722 4654 1727
rect 1929 1712 2006 1717
rect 2025 1712 2246 1717
rect 2433 1712 2494 1717
rect 2537 1712 2758 1717
rect 2849 1712 2982 1717
rect 3017 1712 3046 1717
rect 3177 1712 3246 1717
rect 3417 1712 3462 1717
rect 3545 1712 3670 1717
rect 3689 1712 3854 1717
rect 3897 1712 3942 1717
rect 4017 1712 4046 1717
rect 4105 1712 4190 1717
rect 4313 1712 4350 1717
rect 4457 1712 4518 1717
rect 1033 1707 1038 1712
rect 233 1702 262 1707
rect 257 1697 262 1702
rect 361 1702 486 1707
rect 505 1702 534 1707
rect 361 1697 366 1702
rect 257 1692 366 1697
rect 481 1697 486 1702
rect 529 1697 534 1702
rect 617 1702 838 1707
rect 953 1702 1038 1707
rect 1201 1707 1206 1712
rect 1801 1707 1910 1712
rect 1201 1702 1382 1707
rect 1457 1702 1806 1707
rect 1905 1702 1934 1707
rect 2057 1702 2166 1707
rect 2601 1702 2718 1707
rect 3129 1702 3190 1707
rect 3393 1702 3478 1707
rect 3705 1702 3814 1707
rect 617 1697 622 1702
rect 1377 1697 1462 1702
rect 3809 1697 3814 1702
rect 3881 1702 4006 1707
rect 3881 1697 3886 1702
rect 481 1692 502 1697
rect 529 1692 622 1697
rect 1129 1692 1182 1697
rect 1609 1692 1942 1697
rect 2385 1692 2526 1697
rect 2545 1692 2582 1697
rect 2697 1692 2726 1697
rect 2745 1692 3110 1697
rect 3265 1692 3334 1697
rect 3809 1692 3886 1697
rect 4001 1697 4006 1702
rect 4121 1702 4374 1707
rect 4121 1697 4126 1702
rect 4001 1692 4126 1697
rect 4145 1692 4190 1697
rect 2385 1687 2390 1692
rect 985 1682 1598 1687
rect 1849 1682 2390 1687
rect 2521 1687 2526 1692
rect 2745 1687 2750 1692
rect 3105 1687 3270 1692
rect 3329 1687 3334 1692
rect 4185 1687 4190 1692
rect 4385 1692 4478 1697
rect 4385 1687 4390 1692
rect 2521 1682 2750 1687
rect 3329 1682 3358 1687
rect 3385 1682 3446 1687
rect 4185 1682 4390 1687
rect 1593 1677 1598 1682
rect 1697 1677 1854 1682
rect 937 1672 990 1677
rect 1593 1672 1702 1677
rect 1873 1672 1902 1677
rect 2017 1672 2046 1677
rect 2401 1672 2606 1677
rect 2761 1672 3454 1677
rect 3905 1672 4038 1677
rect 1081 1667 1230 1672
rect 1897 1667 2022 1672
rect 2601 1667 2766 1672
rect 3905 1667 3910 1672
rect 857 1662 926 1667
rect 1001 1662 1086 1667
rect 1225 1662 1254 1667
rect 1273 1662 1398 1667
rect 921 1657 1006 1662
rect 1273 1657 1278 1662
rect 1097 1652 1278 1657
rect 1393 1657 1398 1662
rect 1441 1662 1574 1667
rect 1441 1657 1446 1662
rect 1393 1652 1446 1657
rect 1569 1657 1574 1662
rect 1721 1662 1814 1667
rect 2385 1662 2414 1667
rect 3081 1662 3166 1667
rect 3417 1662 3494 1667
rect 3881 1662 3910 1667
rect 4033 1667 4038 1672
rect 4081 1672 4166 1677
rect 4081 1667 4086 1672
rect 4033 1662 4086 1667
rect 4161 1667 4166 1672
rect 4521 1672 4646 1677
rect 4521 1667 4526 1672
rect 4161 1662 4526 1667
rect 4641 1667 4646 1672
rect 4641 1662 4670 1667
rect 1721 1657 1726 1662
rect 1569 1652 1726 1657
rect 1809 1657 1814 1662
rect 2409 1657 2582 1662
rect 2961 1657 3086 1662
rect 3161 1657 3422 1662
rect 1809 1652 2102 1657
rect 2121 1652 2366 1657
rect 2577 1652 2966 1657
rect 3105 1652 3142 1657
rect 3441 1652 3510 1657
rect 3697 1652 3782 1657
rect 3809 1652 3902 1657
rect 4097 1652 4150 1657
rect 2121 1647 2126 1652
rect 185 1642 230 1647
rect 441 1642 1462 1647
rect 1737 1642 2126 1647
rect 2361 1647 2366 1652
rect 3697 1647 3702 1652
rect 2361 1642 2558 1647
rect 1457 1637 1558 1642
rect 329 1632 398 1637
rect 1193 1632 1358 1637
rect 1369 1632 1438 1637
rect 329 1627 334 1632
rect 161 1622 182 1627
rect 193 1622 334 1627
rect 393 1627 398 1632
rect 1001 1627 1078 1632
rect 1553 1627 1558 1637
rect 1737 1627 1742 1642
rect 2553 1637 2558 1642
rect 2985 1642 3310 1647
rect 3329 1642 3414 1647
rect 3457 1642 3518 1647
rect 3529 1642 3582 1647
rect 3617 1642 3702 1647
rect 3777 1647 3782 1652
rect 3921 1647 4054 1652
rect 4441 1647 4550 1652
rect 3777 1642 3806 1647
rect 3857 1642 3926 1647
rect 4049 1642 4446 1647
rect 4545 1642 4630 1647
rect 2985 1637 2990 1642
rect 1761 1632 1790 1637
rect 393 1622 510 1627
rect 833 1622 1006 1627
rect 1073 1622 1102 1627
rect 1233 1622 1350 1627
rect 1489 1622 1534 1627
rect 1553 1622 1742 1627
rect 1785 1627 1790 1632
rect 1913 1632 2094 1637
rect 2553 1632 2990 1637
rect 3097 1632 3134 1637
rect 3241 1632 3398 1637
rect 3473 1632 3574 1637
rect 3865 1632 3886 1637
rect 3937 1632 4534 1637
rect 1913 1627 1918 1632
rect 1785 1622 1918 1627
rect 1937 1622 1966 1627
rect 1121 1617 1214 1622
rect 1961 1617 1966 1622
rect 2049 1622 2390 1627
rect 2409 1622 2438 1627
rect 2465 1622 2534 1627
rect 3257 1622 3342 1627
rect 3449 1622 3566 1627
rect 3713 1622 3926 1627
rect 3937 1622 4118 1627
rect 4305 1622 4334 1627
rect 4489 1622 4606 1627
rect 4673 1622 4782 1627
rect 2049 1617 2054 1622
rect 4329 1617 4494 1622
rect 209 1612 286 1617
rect 321 1612 382 1617
rect 465 1612 574 1617
rect 1017 1612 1126 1617
rect 1209 1612 1366 1617
rect 1961 1612 2054 1617
rect 3009 1612 3046 1617
rect 3353 1612 3406 1617
rect 3609 1612 3710 1617
rect 3721 1612 3974 1617
rect 4033 1612 4094 1617
rect 4161 1612 4198 1617
rect 4577 1612 4622 1617
rect 2385 1607 2526 1612
rect 3969 1607 3974 1612
rect 297 1602 334 1607
rect 689 1602 734 1607
rect 801 1602 838 1607
rect 1089 1602 1238 1607
rect 1617 1602 1750 1607
rect 1257 1597 1366 1602
rect 1617 1597 1622 1602
rect 441 1592 470 1597
rect 545 1592 614 1597
rect 673 1592 1262 1597
rect 1361 1592 1622 1597
rect 1745 1597 1750 1602
rect 1761 1602 1918 1607
rect 1761 1597 1766 1602
rect 1745 1592 1766 1597
rect 1913 1597 1918 1602
rect 2121 1602 2318 1607
rect 2361 1602 2390 1607
rect 2521 1602 2646 1607
rect 3265 1602 3302 1607
rect 3361 1602 3470 1607
rect 3745 1602 3870 1607
rect 3969 1602 4310 1607
rect 4433 1602 4534 1607
rect 2121 1597 2126 1602
rect 1913 1592 2126 1597
rect 2313 1597 2318 1602
rect 2313 1592 2750 1597
rect 3273 1592 3326 1597
rect 3609 1592 3686 1597
rect 3705 1592 3822 1597
rect 3993 1592 4046 1597
rect 4145 1592 4254 1597
rect 4281 1592 4334 1597
rect 3889 1587 3974 1592
rect 681 1582 846 1587
rect 1081 1582 1110 1587
rect 1105 1577 1110 1582
rect 1185 1582 1350 1587
rect 1633 1582 1742 1587
rect 1785 1582 1894 1587
rect 2137 1582 2526 1587
rect 2657 1582 2782 1587
rect 3321 1582 3406 1587
rect 3641 1582 3894 1587
rect 3969 1582 4126 1587
rect 1185 1577 1190 1582
rect 1785 1577 1790 1582
rect 385 1572 662 1577
rect 721 1572 958 1577
rect 1105 1572 1190 1577
rect 1209 1572 1246 1577
rect 1417 1572 1518 1577
rect 1569 1572 1598 1577
rect 1593 1567 1598 1572
rect 1721 1572 1790 1577
rect 1889 1577 1894 1582
rect 2521 1577 2662 1582
rect 1889 1572 2126 1577
rect 1721 1567 1726 1572
rect 593 1562 806 1567
rect 1233 1562 1278 1567
rect 1593 1562 1726 1567
rect 1745 1562 1926 1567
rect 2121 1557 2126 1572
rect 2249 1572 2318 1577
rect 3073 1572 3166 1577
rect 3561 1572 3630 1577
rect 3905 1572 4182 1577
rect 2249 1557 2254 1572
rect 3073 1567 3078 1572
rect 2377 1562 2622 1567
rect 505 1552 582 1557
rect 577 1547 582 1552
rect 673 1552 750 1557
rect 793 1552 862 1557
rect 1129 1552 1278 1557
rect 1745 1552 1902 1557
rect 2121 1552 2254 1557
rect 2617 1557 2622 1562
rect 2793 1562 2838 1567
rect 3049 1562 3078 1567
rect 3161 1567 3166 1572
rect 3625 1567 3910 1572
rect 3161 1562 3206 1567
rect 3425 1562 3542 1567
rect 3929 1562 4326 1567
rect 2793 1557 2798 1562
rect 3425 1557 3430 1562
rect 2617 1552 2798 1557
rect 3017 1552 3150 1557
rect 3393 1552 3430 1557
rect 3537 1557 3542 1562
rect 3537 1552 3902 1557
rect 4201 1552 4238 1557
rect 673 1547 678 1552
rect 3921 1547 4166 1552
rect 4257 1547 4326 1552
rect 577 1542 678 1547
rect 697 1542 726 1547
rect 721 1537 726 1542
rect 793 1542 822 1547
rect 897 1542 950 1547
rect 1097 1542 1150 1547
rect 1465 1542 1502 1547
rect 1753 1542 1782 1547
rect 1873 1542 1918 1547
rect 1945 1542 2046 1547
rect 2481 1542 2526 1547
rect 2537 1542 2598 1547
rect 3329 1542 3398 1547
rect 3457 1542 3558 1547
rect 3569 1542 3598 1547
rect 793 1537 798 1542
rect 1945 1537 1950 1542
rect 289 1532 414 1537
rect 481 1532 534 1537
rect 721 1532 798 1537
rect 977 1532 998 1537
rect 1185 1532 1294 1537
rect 1481 1532 1534 1537
rect 1649 1532 1726 1537
rect 1889 1532 1950 1537
rect 2041 1537 2046 1542
rect 3593 1537 3598 1542
rect 3697 1542 3926 1547
rect 4161 1542 4190 1547
rect 4233 1542 4262 1547
rect 4321 1542 4398 1547
rect 4713 1542 4774 1547
rect 3697 1537 3702 1542
rect 2041 1532 2070 1537
rect 2473 1532 2550 1537
rect 3081 1532 3118 1537
rect 3185 1532 3214 1537
rect 3593 1532 3702 1537
rect 3721 1532 3766 1537
rect 3873 1532 4310 1537
rect 4545 1532 4646 1537
rect 1185 1527 1190 1532
rect 233 1522 358 1527
rect 465 1522 526 1527
rect 569 1522 662 1527
rect 1017 1522 1190 1527
rect 1289 1527 1294 1532
rect 1649 1527 1654 1532
rect 1721 1527 1870 1532
rect 3761 1527 3766 1532
rect 4329 1527 4438 1532
rect 4545 1527 4550 1532
rect 1289 1522 1326 1527
rect 1553 1522 1582 1527
rect 1625 1522 1654 1527
rect 1865 1522 1998 1527
rect 2153 1522 2246 1527
rect 2601 1522 2686 1527
rect 2913 1522 3062 1527
rect 3193 1522 3246 1527
rect 3393 1522 3470 1527
rect 3761 1522 3790 1527
rect 3809 1522 3990 1527
rect 4217 1522 4334 1527
rect 4433 1522 4462 1527
rect 4481 1522 4550 1527
rect 4641 1527 4646 1532
rect 4641 1522 4702 1527
rect 569 1517 574 1522
rect 129 1512 174 1517
rect 193 1512 238 1517
rect 257 1512 302 1517
rect 313 1512 334 1517
rect 361 1512 390 1517
rect 385 1507 390 1512
rect 505 1512 574 1517
rect 657 1517 662 1522
rect 2153 1517 2158 1522
rect 657 1512 686 1517
rect 785 1512 966 1517
rect 993 1512 1038 1517
rect 1073 1512 1158 1517
rect 1185 1512 1278 1517
rect 1345 1512 1590 1517
rect 1601 1512 1646 1517
rect 1665 1512 2158 1517
rect 2241 1517 2246 1522
rect 2241 1512 2270 1517
rect 2481 1512 2638 1517
rect 505 1507 510 1512
rect 249 1502 294 1507
rect 385 1502 510 1507
rect 905 1502 942 1507
rect 609 1497 774 1502
rect 961 1497 966 1512
rect 1345 1507 1350 1512
rect 1057 1502 1086 1507
rect 1137 1502 1166 1507
rect 1057 1497 1062 1502
rect 185 1492 254 1497
rect 585 1492 614 1497
rect 769 1492 798 1497
rect 961 1492 1062 1497
rect 1161 1497 1166 1502
rect 1289 1502 1350 1507
rect 1585 1507 1590 1512
rect 1585 1502 1630 1507
rect 1289 1497 1294 1502
rect 1161 1492 1294 1497
rect 793 1487 798 1492
rect 593 1482 774 1487
rect 793 1482 894 1487
rect 889 1477 894 1482
rect 1313 1482 1462 1487
rect 1313 1477 1318 1482
rect 889 1472 1318 1477
rect 1457 1477 1462 1482
rect 1665 1477 1670 1512
rect 2913 1507 2918 1522
rect 1713 1502 1758 1507
rect 1865 1502 1990 1507
rect 2169 1502 2246 1507
rect 2273 1502 2302 1507
rect 2889 1502 2918 1507
rect 3057 1507 3062 1522
rect 4081 1517 4198 1522
rect 4697 1517 4702 1522
rect 4777 1522 4806 1527
rect 4777 1517 4782 1522
rect 3113 1512 3206 1517
rect 3745 1512 3774 1517
rect 3769 1507 3774 1512
rect 3889 1512 3950 1517
rect 4057 1512 4086 1517
rect 4193 1512 4534 1517
rect 4697 1512 4782 1517
rect 3889 1507 3894 1512
rect 3057 1502 3118 1507
rect 2561 1497 2686 1502
rect 3113 1497 3118 1502
rect 3217 1502 3334 1507
rect 3449 1502 3526 1507
rect 3545 1502 3726 1507
rect 3769 1502 3894 1507
rect 3913 1502 4238 1507
rect 4249 1502 4398 1507
rect 4521 1502 4630 1507
rect 3217 1497 3222 1502
rect 1753 1492 1782 1497
rect 1457 1472 1670 1477
rect 1777 1477 1782 1492
rect 1929 1492 1974 1497
rect 2385 1492 2566 1497
rect 2681 1492 3094 1497
rect 3113 1492 3222 1497
rect 3945 1492 3974 1497
rect 3985 1492 4014 1497
rect 1929 1477 1934 1492
rect 2177 1487 2294 1492
rect 2073 1482 2182 1487
rect 2289 1482 2430 1487
rect 1777 1472 1934 1477
rect 1993 1472 2062 1477
rect 2057 1467 2062 1472
rect 2193 1472 2278 1477
rect 2193 1467 2198 1472
rect 689 1462 838 1467
rect 2057 1462 2198 1467
rect 2425 1467 2430 1482
rect 2577 1482 2670 1487
rect 2577 1467 2582 1482
rect 2425 1462 2582 1467
rect 2665 1467 2670 1482
rect 2833 1482 2862 1487
rect 2833 1467 2838 1482
rect 3089 1477 3094 1492
rect 3945 1487 3950 1492
rect 3737 1482 3950 1487
rect 4009 1487 4014 1492
rect 4081 1492 4166 1497
rect 4081 1487 4086 1492
rect 4009 1482 4086 1487
rect 4113 1482 4142 1487
rect 3737 1477 3742 1482
rect 3089 1472 3742 1477
rect 4137 1477 4142 1482
rect 4289 1482 4342 1487
rect 4289 1477 4294 1482
rect 4137 1472 4294 1477
rect 4337 1477 4342 1482
rect 4409 1482 4462 1487
rect 4409 1477 4414 1482
rect 4337 1472 4414 1477
rect 2665 1462 2838 1467
rect 473 1452 646 1457
rect 473 1447 478 1452
rect 265 1442 478 1447
rect 641 1447 646 1452
rect 689 1447 694 1462
rect 641 1442 694 1447
rect 833 1447 838 1462
rect 881 1452 974 1457
rect 1337 1452 1438 1457
rect 1641 1452 1742 1457
rect 2217 1452 2406 1457
rect 2601 1452 2646 1457
rect 2945 1452 3070 1457
rect 881 1447 886 1452
rect 833 1442 886 1447
rect 969 1447 974 1452
rect 1641 1447 1646 1452
rect 969 1442 1646 1447
rect 1737 1447 1742 1452
rect 1737 1442 1766 1447
rect 2001 1442 2254 1447
rect 2881 1442 2926 1447
rect 2945 1437 2950 1452
rect 145 1432 230 1437
rect 401 1432 430 1437
rect 489 1432 574 1437
rect 425 1427 494 1432
rect 569 1427 574 1432
rect 673 1432 958 1437
rect 1393 1432 1510 1437
rect 1657 1432 1742 1437
rect 1993 1432 2022 1437
rect 2537 1432 2598 1437
rect 2633 1432 2670 1437
rect 2761 1432 2950 1437
rect 3065 1437 3070 1452
rect 3065 1432 3118 1437
rect 3297 1432 3366 1437
rect 3585 1432 3710 1437
rect 673 1427 678 1432
rect 3585 1427 3590 1432
rect 65 1422 150 1427
rect 177 1422 246 1427
rect 569 1422 678 1427
rect 697 1422 750 1427
rect 801 1422 846 1427
rect 1217 1422 1262 1427
rect 1481 1422 1566 1427
rect 1625 1422 1670 1427
rect 1969 1422 2014 1427
rect 2625 1422 2662 1427
rect 2721 1422 2750 1427
rect 2745 1417 2750 1422
rect 2825 1422 3198 1427
rect 3537 1422 3590 1427
rect 3705 1427 3710 1432
rect 3969 1432 4038 1437
rect 3969 1427 3974 1432
rect 3705 1422 3822 1427
rect 3945 1422 3974 1427
rect 4033 1427 4038 1432
rect 4129 1432 4198 1437
rect 4129 1427 4134 1432
rect 4033 1422 4134 1427
rect 4193 1427 4198 1432
rect 4249 1432 4414 1437
rect 4193 1422 4222 1427
rect 2825 1417 2830 1422
rect 65 1412 86 1417
rect 425 1412 550 1417
rect 753 1412 822 1417
rect 921 1412 998 1417
rect 1025 1412 1070 1417
rect 1137 1412 1174 1417
rect 1281 1412 1374 1417
rect 1961 1412 2030 1417
rect 2745 1412 2830 1417
rect 1193 1407 1286 1412
rect 1369 1407 1374 1412
rect 369 1402 422 1407
rect 1033 1402 1198 1407
rect 1369 1402 1702 1407
rect 1945 1402 1974 1407
rect 81 1392 158 1397
rect 185 1392 382 1397
rect 409 1392 862 1397
rect 897 1392 1070 1397
rect 1081 1392 1142 1397
rect 1169 1392 1350 1397
rect 1753 1392 1790 1397
rect 1817 1392 1910 1397
rect 1993 1392 2126 1397
rect 2145 1392 2190 1397
rect 2465 1392 2766 1397
rect 2849 1392 2854 1422
rect 4249 1417 4254 1432
rect 3017 1412 3134 1417
rect 3561 1412 3694 1417
rect 4145 1412 4190 1417
rect 4217 1412 4254 1417
rect 4409 1417 4414 1432
rect 4433 1422 4542 1427
rect 4601 1422 4662 1427
rect 4409 1412 4598 1417
rect 4593 1407 4598 1412
rect 4665 1412 4710 1417
rect 4665 1407 4670 1412
rect 2873 1402 2902 1407
rect 2897 1397 2902 1402
rect 2985 1402 3014 1407
rect 3401 1402 3598 1407
rect 2985 1397 2990 1402
rect 2897 1392 2990 1397
rect 3593 1397 3598 1402
rect 3833 1402 4022 1407
rect 4265 1402 4334 1407
rect 4393 1402 4478 1407
rect 4593 1402 4670 1407
rect 3833 1397 3838 1402
rect 3593 1392 3838 1397
rect 1521 1387 1630 1392
rect 4449 1387 4542 1392
rect 217 1382 254 1387
rect 1025 1382 1070 1387
rect 1137 1382 1526 1387
rect 1625 1382 1710 1387
rect 2001 1382 2038 1387
rect 2601 1382 2638 1387
rect 2745 1382 2830 1387
rect 3089 1382 3150 1387
rect 4425 1382 4454 1387
rect 4537 1382 4566 1387
rect 4633 1382 4662 1387
rect 1785 1377 1982 1382
rect 209 1372 326 1377
rect 321 1367 326 1372
rect 441 1372 470 1377
rect 737 1372 822 1377
rect 1001 1372 1358 1377
rect 1553 1372 1614 1377
rect 1737 1372 1790 1377
rect 1977 1372 2054 1377
rect 3489 1372 3574 1377
rect 441 1367 446 1372
rect 737 1367 742 1372
rect 177 1362 206 1367
rect 321 1362 446 1367
rect 505 1362 742 1367
rect 817 1367 822 1372
rect 1353 1367 1558 1372
rect 3489 1367 3494 1372
rect 817 1362 846 1367
rect 1185 1362 1334 1367
rect 1577 1362 2022 1367
rect 2137 1362 2238 1367
rect 2889 1362 3070 1367
rect 2889 1357 2894 1362
rect 753 1352 822 1357
rect 865 1352 982 1357
rect 865 1347 870 1352
rect 233 1342 294 1347
rect 649 1342 750 1347
rect 841 1342 870 1347
rect 977 1347 982 1352
rect 993 1352 1102 1357
rect 1129 1352 1166 1357
rect 1257 1352 1526 1357
rect 1705 1352 1854 1357
rect 2065 1352 2262 1357
rect 2849 1352 2894 1357
rect 3065 1357 3070 1362
rect 3393 1362 3494 1367
rect 3569 1367 3574 1372
rect 3937 1372 4022 1377
rect 3937 1367 3942 1372
rect 3569 1362 3942 1367
rect 4017 1367 4022 1372
rect 4161 1372 4294 1377
rect 4313 1372 4566 1377
rect 4161 1367 4166 1372
rect 4017 1362 4046 1367
rect 4137 1362 4166 1367
rect 4289 1367 4294 1372
rect 4561 1367 4566 1372
rect 4289 1362 4318 1367
rect 4449 1362 4542 1367
rect 4561 1362 4774 1367
rect 3393 1357 3398 1362
rect 4313 1357 4454 1362
rect 3065 1352 3398 1357
rect 3513 1352 3558 1357
rect 3953 1352 4278 1357
rect 993 1347 998 1352
rect 977 1342 998 1347
rect 1097 1347 1102 1352
rect 1849 1347 1958 1352
rect 2065 1347 2070 1352
rect 4273 1347 4278 1352
rect 4473 1352 4502 1357
rect 4473 1347 4478 1352
rect 1097 1342 1142 1347
rect 1153 1342 1270 1347
rect 1745 1342 1830 1347
rect 1953 1342 2070 1347
rect 2145 1342 2366 1347
rect 2417 1342 2534 1347
rect 1625 1337 1702 1342
rect 2417 1337 2422 1342
rect 177 1332 230 1337
rect 289 1332 334 1337
rect 441 1332 598 1337
rect 617 1332 862 1337
rect 1009 1332 1326 1337
rect 1449 1332 1534 1337
rect 1601 1332 1630 1337
rect 1697 1332 1734 1337
rect 1841 1332 1934 1337
rect 2113 1332 2214 1337
rect 2297 1332 2342 1337
rect 2393 1332 2422 1337
rect 2529 1337 2534 1342
rect 2585 1342 2718 1347
rect 3025 1342 3102 1347
rect 3361 1342 3430 1347
rect 3441 1342 3534 1347
rect 4025 1342 4070 1347
rect 4273 1342 4478 1347
rect 4553 1342 4598 1347
rect 4689 1342 4750 1347
rect 2529 1332 2558 1337
rect 177 1322 182 1332
rect 441 1327 446 1332
rect 361 1322 446 1327
rect 593 1327 598 1332
rect 1449 1327 1454 1332
rect 593 1322 910 1327
rect 961 1322 1454 1327
rect 1529 1327 1534 1332
rect 1729 1327 1846 1332
rect 2585 1327 2590 1342
rect 1529 1322 1558 1327
rect 1649 1322 1686 1327
rect 2121 1322 2158 1327
rect 2361 1322 2590 1327
rect 2713 1327 2718 1342
rect 2905 1332 2966 1337
rect 3193 1332 3286 1337
rect 3305 1332 3366 1337
rect 3193 1327 3198 1332
rect 2713 1322 2742 1327
rect 2833 1322 2854 1327
rect 3137 1322 3198 1327
rect 3281 1327 3286 1332
rect 3361 1327 3366 1332
rect 3457 1332 3502 1337
rect 3593 1332 4054 1337
rect 4577 1332 4630 1337
rect 3457 1327 3462 1332
rect 3281 1322 3342 1327
rect 3361 1322 3462 1327
rect 3481 1322 3550 1327
rect 4057 1322 4230 1327
rect 4265 1322 4414 1327
rect 4713 1322 4734 1327
rect 457 1312 574 1317
rect 721 1312 766 1317
rect 801 1312 838 1317
rect 849 1312 902 1317
rect 961 1312 966 1322
rect 2833 1317 2838 1322
rect 977 1312 1046 1317
rect 1057 1312 1142 1317
rect 1249 1312 1358 1317
rect 1465 1312 1558 1317
rect 1601 1312 1638 1317
rect 1761 1312 1790 1317
rect 1817 1312 1862 1317
rect 2105 1312 2182 1317
rect 2201 1312 2222 1317
rect 2601 1312 2702 1317
rect 2801 1312 2838 1317
rect 3209 1312 3318 1317
rect 3337 1307 3342 1322
rect 3481 1307 3486 1322
rect 3577 1312 3614 1317
rect 3713 1312 3750 1317
rect 4033 1312 4054 1317
rect 4225 1312 4230 1322
rect 4377 1312 4438 1317
rect 4537 1312 4678 1317
rect 465 1297 470 1307
rect 497 1302 606 1307
rect 657 1302 766 1307
rect 881 1302 934 1307
rect 1017 1302 1062 1307
rect 1161 1302 1270 1307
rect 1345 1302 1486 1307
rect 2073 1302 2102 1307
rect 3065 1302 3294 1307
rect 3337 1302 3486 1307
rect 3593 1302 3630 1307
rect 3729 1302 3838 1307
rect 4033 1302 4086 1307
rect 4505 1302 4526 1307
rect 1513 1297 1638 1302
rect 465 1292 494 1297
rect 889 1292 918 1297
rect 1033 1292 1198 1297
rect 489 1287 694 1292
rect 689 1277 694 1287
rect 889 1277 894 1292
rect 1193 1287 1198 1292
rect 1281 1292 1374 1297
rect 1497 1292 1518 1297
rect 1633 1292 1742 1297
rect 1753 1292 1782 1297
rect 2313 1292 2582 1297
rect 1281 1287 1286 1292
rect 1369 1287 1502 1292
rect 1193 1282 1286 1287
rect 1305 1282 1350 1287
rect 1345 1277 1350 1282
rect 1521 1282 1750 1287
rect 1521 1277 1526 1282
rect 2313 1277 2318 1292
rect 2577 1287 2582 1292
rect 2857 1292 3046 1297
rect 3185 1292 3214 1297
rect 3569 1292 3710 1297
rect 2857 1287 2862 1292
rect 2577 1282 2862 1287
rect 3041 1287 3046 1292
rect 3041 1282 3142 1287
rect 409 1272 670 1277
rect 689 1272 894 1277
rect 1081 1272 1174 1277
rect 1345 1272 1526 1277
rect 2289 1272 2318 1277
rect 3137 1277 3142 1282
rect 3225 1277 3294 1282
rect 3137 1272 3230 1277
rect 3289 1272 3390 1277
rect 4433 1272 4518 1277
rect 4433 1267 4438 1272
rect 2249 1262 3126 1267
rect 3241 1262 3278 1267
rect 4409 1262 4438 1267
rect 4513 1267 4518 1272
rect 4513 1262 4702 1267
rect 513 1252 550 1257
rect 913 1252 1494 1257
rect 2665 1252 2686 1257
rect 2865 1252 2902 1257
rect 3233 1252 3278 1257
rect 3337 1252 3382 1257
rect 3609 1252 3774 1257
rect 2377 1247 2454 1252
rect 265 1242 358 1247
rect 553 1242 702 1247
rect 721 1242 838 1247
rect 2353 1242 2382 1247
rect 2449 1242 2758 1247
rect 2769 1242 3006 1247
rect 3033 1242 3062 1247
rect 3113 1242 3262 1247
rect 3329 1242 3366 1247
rect 3569 1242 3590 1247
rect 265 1237 270 1242
rect 161 1232 270 1237
rect 353 1237 358 1242
rect 721 1237 726 1242
rect 3609 1237 3614 1252
rect 353 1232 382 1237
rect 457 1232 726 1237
rect 801 1232 862 1237
rect 985 1232 1070 1237
rect 2329 1232 2438 1237
rect 2601 1232 2630 1237
rect 2785 1232 2870 1237
rect 2889 1232 2918 1237
rect 985 1227 990 1232
rect 129 1222 174 1227
rect 369 1222 406 1227
rect 521 1222 566 1227
rect 649 1222 686 1227
rect 793 1222 822 1227
rect 833 1222 990 1227
rect 1065 1227 1070 1232
rect 1065 1222 1470 1227
rect 1521 1222 1550 1227
rect 1569 1222 1614 1227
rect 2273 1222 2350 1227
rect 2409 1222 2510 1227
rect 2585 1222 2630 1227
rect 2649 1222 2718 1227
rect 161 1212 190 1217
rect 281 1212 326 1217
rect 465 1212 574 1217
rect 673 1212 726 1217
rect 761 1212 846 1217
rect 1001 1212 1054 1217
rect 2321 1212 2358 1217
rect 2865 1212 2870 1232
rect 2913 1227 2918 1232
rect 3049 1232 3086 1237
rect 3185 1232 3318 1237
rect 3353 1232 3414 1237
rect 3521 1232 3614 1237
rect 3769 1237 3774 1252
rect 3857 1252 4222 1257
rect 3857 1237 3862 1252
rect 4217 1237 4222 1252
rect 4241 1242 4342 1247
rect 4441 1242 4502 1247
rect 3769 1232 3798 1237
rect 3833 1232 3862 1237
rect 3961 1232 4062 1237
rect 4217 1232 4646 1237
rect 3049 1227 3054 1232
rect 3521 1227 3526 1232
rect 3961 1227 3966 1232
rect 2913 1222 3054 1227
rect 3073 1222 3102 1227
rect 3225 1222 3254 1227
rect 3345 1222 3526 1227
rect 3537 1222 3622 1227
rect 3633 1222 3966 1227
rect 4057 1227 4062 1232
rect 4057 1222 4086 1227
rect 4193 1222 4270 1227
rect 4369 1222 4422 1227
rect 4473 1222 4518 1227
rect 4633 1222 4726 1227
rect 3633 1217 3638 1222
rect 3561 1212 3638 1217
rect 3673 1212 3846 1217
rect 3865 1212 4182 1217
rect 4281 1212 4550 1217
rect 4561 1212 4614 1217
rect 161 1187 166 1212
rect 4177 1207 4286 1212
rect 257 1202 438 1207
rect 713 1202 750 1207
rect 849 1202 982 1207
rect 993 1202 1078 1207
rect 977 1197 982 1202
rect 1073 1197 1078 1202
rect 1185 1202 1326 1207
rect 2713 1202 3126 1207
rect 1185 1197 1190 1202
rect 3121 1197 3126 1202
rect 3217 1202 3286 1207
rect 3305 1202 3366 1207
rect 3481 1202 3542 1207
rect 3737 1202 3822 1207
rect 3969 1202 4134 1207
rect 3217 1197 3222 1202
rect 361 1192 390 1197
rect 385 1187 390 1192
rect 457 1192 630 1197
rect 721 1192 966 1197
rect 977 1192 1030 1197
rect 1073 1192 1190 1197
rect 1209 1192 1238 1197
rect 1529 1192 1582 1197
rect 1945 1192 2046 1197
rect 2273 1192 2310 1197
rect 2601 1192 2678 1197
rect 3121 1192 3222 1197
rect 3281 1197 3286 1202
rect 3601 1197 3670 1202
rect 4129 1197 4134 1202
rect 4305 1202 4438 1207
rect 4305 1197 4310 1202
rect 4481 1197 4630 1202
rect 3281 1192 3494 1197
rect 457 1187 462 1192
rect 3489 1187 3494 1192
rect 3577 1192 3606 1197
rect 3665 1192 3854 1197
rect 3913 1192 3966 1197
rect 4057 1192 4110 1197
rect 4129 1192 4310 1197
rect 4329 1192 4358 1197
rect 4449 1192 4486 1197
rect 4625 1192 4718 1197
rect 3577 1187 3582 1192
rect 4353 1187 4454 1192
rect 161 1182 206 1187
rect 385 1182 462 1187
rect 657 1182 926 1187
rect 1681 1182 1926 1187
rect 2137 1182 2246 1187
rect 2321 1182 2414 1187
rect 2577 1182 2614 1187
rect 2905 1182 3022 1187
rect 3233 1182 3342 1187
rect 3489 1182 3582 1187
rect 3601 1182 3654 1187
rect 3737 1182 3798 1187
rect 3841 1182 3934 1187
rect 4497 1182 4590 1187
rect 777 1172 1054 1177
rect 1441 1172 1510 1177
rect 1441 1167 1446 1172
rect 185 1162 214 1167
rect 481 1162 542 1167
rect 657 1162 806 1167
rect 833 1162 910 1167
rect 1289 1162 1406 1167
rect 1417 1162 1446 1167
rect 1505 1167 1510 1172
rect 1681 1167 1686 1182
rect 1921 1177 1926 1182
rect 2241 1177 2326 1182
rect 3649 1177 3742 1182
rect 4217 1177 4302 1182
rect 1921 1172 2118 1177
rect 2617 1172 2710 1177
rect 3233 1172 3286 1177
rect 3297 1172 3366 1177
rect 3921 1172 3958 1177
rect 3977 1172 4094 1177
rect 4193 1172 4222 1177
rect 4297 1172 4678 1177
rect 1505 1162 1558 1167
rect 1569 1162 1686 1167
rect 2113 1167 2118 1172
rect 3977 1167 3982 1172
rect 2113 1162 2230 1167
rect 2241 1162 2462 1167
rect 2625 1162 2662 1167
rect 2873 1162 2990 1167
rect 3721 1162 3982 1167
rect 4089 1167 4094 1172
rect 4089 1162 4182 1167
rect 2873 1157 2878 1162
rect 689 1152 718 1157
rect 713 1147 718 1152
rect 793 1152 894 1157
rect 793 1147 798 1152
rect 441 1142 486 1147
rect 561 1142 646 1147
rect 713 1142 798 1147
rect 889 1147 894 1152
rect 1065 1152 1614 1157
rect 1697 1152 2086 1157
rect 1065 1147 1070 1152
rect 1609 1147 1702 1152
rect 2081 1147 2086 1152
rect 2145 1152 2174 1157
rect 2401 1152 2494 1157
rect 2849 1152 2878 1157
rect 2985 1157 2990 1162
rect 4177 1157 4182 1162
rect 4257 1162 4286 1167
rect 4409 1162 4686 1167
rect 4257 1157 4262 1162
rect 2985 1152 3014 1157
rect 3105 1152 3150 1157
rect 3257 1152 3334 1157
rect 3553 1152 3590 1157
rect 3897 1152 4078 1157
rect 4177 1152 4262 1157
rect 4281 1152 4334 1157
rect 4393 1152 4598 1157
rect 4705 1152 4758 1157
rect 2145 1147 2150 1152
rect 889 1142 1070 1147
rect 1233 1142 1414 1147
rect 1409 1137 1414 1142
rect 1497 1142 1590 1147
rect 1921 1142 1990 1147
rect 2081 1142 2150 1147
rect 2225 1142 2382 1147
rect 2409 1142 2438 1147
rect 2521 1142 2734 1147
rect 2777 1142 2862 1147
rect 2889 1142 2974 1147
rect 3041 1142 3286 1147
rect 3329 1142 3350 1147
rect 3393 1142 3454 1147
rect 3577 1142 3670 1147
rect 3697 1142 3814 1147
rect 3929 1142 4046 1147
rect 4297 1142 4326 1147
rect 4449 1142 4510 1147
rect 4585 1142 4726 1147
rect 1497 1137 1502 1142
rect 1921 1137 1926 1142
rect 2433 1137 2526 1142
rect 2969 1137 3046 1142
rect 3281 1137 3286 1142
rect 529 1132 614 1137
rect 817 1132 870 1137
rect 1337 1132 1390 1137
rect 1409 1132 1502 1137
rect 1649 1132 1694 1137
rect 1721 1132 1926 1137
rect 1945 1132 2062 1137
rect 3185 1132 3246 1137
rect 3281 1132 3358 1137
rect 3353 1127 3358 1132
rect 3449 1132 3734 1137
rect 3449 1127 3454 1132
rect 2449 1122 2550 1127
rect 2617 1122 2646 1127
rect 2897 1122 2974 1127
rect 2993 1122 3022 1127
rect 3113 1122 3182 1127
rect 3353 1122 3454 1127
rect 3729 1127 3734 1132
rect 3801 1132 3830 1137
rect 3905 1132 3950 1137
rect 3801 1127 3806 1132
rect 3969 1127 3974 1137
rect 4457 1132 4486 1137
rect 3729 1122 3806 1127
rect 3929 1122 3974 1127
rect 4057 1122 4238 1127
rect 1665 1117 1758 1122
rect 2449 1117 2454 1122
rect 81 1112 110 1117
rect 585 1112 638 1117
rect 1081 1112 1198 1117
rect 1521 1112 1670 1117
rect 1753 1112 1894 1117
rect 2033 1112 2086 1117
rect 2329 1112 2390 1117
rect 2425 1112 2454 1117
rect 2545 1117 2550 1122
rect 2897 1117 2902 1122
rect 2545 1112 2638 1117
rect 2689 1112 2902 1117
rect 2969 1117 2974 1122
rect 2969 1112 3126 1117
rect 3137 1112 3246 1117
rect 3305 1112 3334 1117
rect 3121 1107 3126 1112
rect 3329 1107 3334 1112
rect 3473 1112 3574 1117
rect 3585 1112 3710 1117
rect 3905 1112 3942 1117
rect 4225 1112 4302 1117
rect 4313 1112 4358 1117
rect 4465 1112 4582 1117
rect 4625 1112 4678 1117
rect 4689 1112 4710 1117
rect 3473 1107 3478 1112
rect 577 1102 614 1107
rect 1057 1102 1086 1107
rect 1081 1097 1086 1102
rect 1193 1102 1222 1107
rect 1369 1102 1446 1107
rect 1465 1102 1510 1107
rect 1681 1102 1758 1107
rect 1969 1102 2054 1107
rect 2153 1102 2174 1107
rect 2433 1102 2478 1107
rect 2505 1102 2534 1107
rect 2617 1102 2654 1107
rect 2897 1102 3014 1107
rect 3081 1102 3102 1107
rect 3121 1102 3286 1107
rect 3329 1102 3478 1107
rect 3569 1107 3574 1112
rect 3569 1102 3702 1107
rect 4329 1102 4414 1107
rect 4497 1102 4590 1107
rect 1193 1097 1198 1102
rect 1969 1097 1974 1102
rect 865 1092 886 1097
rect 1081 1092 1198 1097
rect 1473 1092 1518 1097
rect 1513 1087 1518 1092
rect 1825 1092 1974 1097
rect 2401 1092 2470 1097
rect 3097 1092 3134 1097
rect 3537 1092 3670 1097
rect 3681 1092 3710 1097
rect 1825 1087 1830 1092
rect 3665 1087 3670 1092
rect 681 1082 910 1087
rect 1513 1082 1830 1087
rect 2417 1082 2502 1087
rect 3665 1082 3686 1087
rect 4257 1082 4350 1087
rect 4257 1077 4262 1082
rect 3953 1072 4070 1077
rect 809 1062 1062 1067
rect 1401 1062 1494 1067
rect 2761 1062 2942 1067
rect 1401 1057 1406 1062
rect 281 1052 798 1057
rect 793 1047 798 1052
rect 897 1052 926 1057
rect 1073 1052 1406 1057
rect 1489 1057 1494 1062
rect 3953 1057 3958 1072
rect 4065 1067 4070 1072
rect 4113 1072 4214 1077
rect 4233 1072 4262 1077
rect 4345 1077 4350 1082
rect 4345 1072 4430 1077
rect 4113 1067 4118 1072
rect 4065 1062 4118 1067
rect 4209 1067 4214 1072
rect 4209 1062 4334 1067
rect 1489 1052 1630 1057
rect 3041 1052 3078 1057
rect 3177 1052 3302 1057
rect 897 1047 902 1052
rect 3177 1047 3182 1052
rect 793 1042 902 1047
rect 1921 1042 2030 1047
rect 2049 1042 2150 1047
rect 2473 1042 2622 1047
rect 3081 1042 3182 1047
rect 3297 1047 3302 1052
rect 3705 1052 3790 1057
rect 3809 1052 3958 1057
rect 4081 1052 4214 1057
rect 4353 1052 4454 1057
rect 3705 1047 3710 1052
rect 3297 1042 3358 1047
rect 3681 1042 3710 1047
rect 3785 1047 3790 1052
rect 4353 1047 4358 1052
rect 3785 1042 4358 1047
rect 4449 1047 4454 1052
rect 4449 1042 4502 1047
rect 89 1032 182 1037
rect 1417 1032 1478 1037
rect 1593 1032 1678 1037
rect 1721 1032 1806 1037
rect 1921 1027 1926 1042
rect 2025 1037 2030 1042
rect 2473 1037 2478 1042
rect 2025 1032 2062 1037
rect 2313 1032 2358 1037
rect 2449 1032 2478 1037
rect 2617 1037 2622 1042
rect 2617 1032 2686 1037
rect 2769 1032 2870 1037
rect 73 1022 182 1027
rect 225 1022 254 1027
rect 289 1022 334 1027
rect 537 1022 734 1027
rect 801 1022 846 1027
rect 881 1022 910 1027
rect 921 1022 1078 1027
rect 1121 1022 1750 1027
rect 1825 1022 1926 1027
rect 1937 1022 1982 1027
rect 2129 1022 2198 1027
rect 2345 1022 2406 1027
rect 2497 1022 2582 1027
rect 2673 1022 2694 1027
rect 169 1012 382 1017
rect 401 1012 518 1017
rect 537 1007 542 1022
rect 729 1007 734 1022
rect 1825 1017 1830 1022
rect 2497 1017 2502 1022
rect 753 1012 902 1017
rect 1249 1012 1278 1017
rect 1273 1007 1278 1012
rect 1401 1012 1430 1017
rect 1641 1012 1830 1017
rect 1953 1012 2030 1017
rect 2217 1012 2502 1017
rect 2577 1017 2582 1022
rect 2913 1017 2918 1037
rect 3041 1032 3118 1037
rect 3793 1032 4262 1037
rect 4369 1032 4438 1037
rect 4433 1027 4438 1032
rect 4513 1032 4614 1037
rect 4697 1032 4734 1037
rect 4513 1027 4518 1032
rect 3193 1022 3286 1027
rect 3665 1022 4238 1027
rect 4257 1022 4342 1027
rect 4433 1022 4518 1027
rect 4545 1017 4550 1027
rect 2577 1012 2606 1017
rect 2873 1012 2918 1017
rect 3457 1012 3566 1017
rect 3729 1012 3822 1017
rect 3897 1012 3926 1017
rect 4049 1012 4198 1017
rect 4345 1012 4414 1017
rect 4545 1012 4582 1017
rect 4617 1012 4670 1017
rect 1401 1007 1406 1012
rect 1953 1007 1958 1012
rect 3457 1007 3462 1012
rect 145 1002 214 1007
rect 209 997 214 1002
rect 313 1002 342 1007
rect 369 1002 542 1007
rect 569 1002 710 1007
rect 729 1002 950 1007
rect 1273 1002 1406 1007
rect 1737 1002 1958 1007
rect 2505 1002 2598 1007
rect 2633 1002 2678 1007
rect 3401 1002 3462 1007
rect 3561 1007 3566 1012
rect 3921 1007 4054 1012
rect 4193 1007 4350 1012
rect 3561 1002 3622 1007
rect 4073 1002 4174 1007
rect 4369 1002 4422 1007
rect 4569 1002 4782 1007
rect 313 997 318 1002
rect 569 997 574 1002
rect 129 992 190 997
rect 209 992 318 997
rect 361 992 574 997
rect 705 997 710 1002
rect 705 992 926 997
rect 1193 992 1230 997
rect 1569 992 1694 997
rect 1857 992 1886 997
rect 2705 992 2790 997
rect 3025 992 3054 997
rect 3217 992 3302 997
rect 3473 992 3550 997
rect 3657 992 3742 997
rect 3961 992 4022 997
rect 4057 992 4270 997
rect 4537 992 4566 997
rect 2705 987 2710 992
rect 353 982 382 987
rect 377 977 382 982
rect 585 982 782 987
rect 793 982 1014 987
rect 1073 982 1182 987
rect 585 977 590 982
rect 1177 977 1182 982
rect 1241 982 2054 987
rect 2345 982 2486 987
rect 2513 982 2614 987
rect 1241 977 1246 982
rect 377 972 590 977
rect 609 972 646 977
rect 689 972 806 977
rect 849 972 950 977
rect 1137 972 1158 977
rect 1177 972 1246 977
rect 1609 972 1638 977
rect 1633 967 1638 972
rect 1841 972 1910 977
rect 1841 967 1846 972
rect 1633 962 1846 967
rect 1905 967 1910 972
rect 1993 972 2046 977
rect 1993 967 1998 972
rect 2345 967 2350 982
rect 1905 962 1998 967
rect 2249 962 2350 967
rect 2481 967 2486 982
rect 2609 977 2614 982
rect 2689 982 2710 987
rect 2785 987 2790 992
rect 2785 982 2814 987
rect 3641 982 3950 987
rect 4081 982 4454 987
rect 2689 977 2694 982
rect 3945 977 4086 982
rect 2609 972 2694 977
rect 2793 972 2854 977
rect 3417 972 3558 977
rect 3857 972 3886 977
rect 3417 967 3422 972
rect 2481 962 2518 967
rect 2713 962 2798 967
rect 2841 962 2870 967
rect 3273 962 3374 967
rect 3393 962 3422 967
rect 3553 967 3558 972
rect 3673 967 3790 972
rect 3881 967 3886 972
rect 4105 972 4214 977
rect 4105 967 4110 972
rect 3553 962 3678 967
rect 3785 962 3814 967
rect 3881 962 4110 967
rect 4209 967 4214 972
rect 4465 972 4638 977
rect 4465 967 4470 972
rect 4209 962 4470 967
rect 3273 957 3278 962
rect 505 952 590 957
rect 665 952 838 957
rect 1289 952 1406 957
rect 1865 952 1886 957
rect 2209 952 2238 957
rect 2361 952 2486 957
rect 2713 952 2822 957
rect 2881 952 2998 957
rect 3249 952 3278 957
rect 3369 957 3374 962
rect 3369 952 3478 957
rect 3489 952 3542 957
rect 3689 952 3766 957
rect 4129 952 4190 957
rect 505 947 510 952
rect 481 942 510 947
rect 585 947 590 952
rect 1289 947 1294 952
rect 585 942 654 947
rect 649 937 654 942
rect 729 942 758 947
rect 817 942 854 947
rect 977 942 1174 947
rect 1265 942 1294 947
rect 1401 947 1406 952
rect 1401 942 1430 947
rect 1561 942 1606 947
rect 1641 942 1702 947
rect 1785 942 1806 947
rect 1905 942 2054 947
rect 2185 942 2214 947
rect 2257 942 2310 947
rect 2321 942 2350 947
rect 3017 942 3198 947
rect 3273 942 3358 947
rect 3433 942 3486 947
rect 3753 942 4118 947
rect 4201 942 4454 947
rect 729 937 734 942
rect 873 937 982 942
rect 209 932 366 937
rect 649 932 734 937
rect 825 932 878 937
rect 209 917 214 932
rect 361 927 366 932
rect 1169 927 1174 942
rect 1905 937 1910 942
rect 1649 932 1910 937
rect 2049 937 2054 942
rect 3017 937 3022 942
rect 2049 932 2078 937
rect 2193 932 2350 937
rect 2825 932 3022 937
rect 3193 937 3198 942
rect 3353 937 3438 942
rect 4113 937 4206 942
rect 3193 932 3222 937
rect 3457 932 3502 937
rect 3585 932 3614 937
rect 3657 932 3686 937
rect 4465 932 4494 937
rect 1649 927 1654 932
rect 361 922 390 927
rect 465 922 582 927
rect 833 922 918 927
rect 1017 922 1150 927
rect 1169 922 1654 927
rect 1729 922 1790 927
rect 1929 922 1958 927
rect 2313 922 2542 927
rect 2585 922 2646 927
rect 3105 922 3150 927
rect 3345 922 3374 927
rect 3857 922 3894 927
rect 3953 922 4030 927
rect 4145 922 4254 927
rect 4393 922 4438 927
rect 97 912 214 917
rect 233 912 278 917
rect 337 912 502 917
rect 513 912 606 917
rect 625 912 702 917
rect 993 912 1038 917
rect 1217 912 1278 917
rect 1465 912 1502 917
rect 497 907 502 912
rect 625 907 630 912
rect 185 902 222 907
rect 265 902 350 907
rect 497 902 630 907
rect 697 907 702 912
rect 1497 907 1502 912
rect 1617 912 1646 917
rect 1753 912 1838 917
rect 1881 912 1926 917
rect 1937 912 1982 917
rect 2025 912 2046 917
rect 2529 912 2638 917
rect 2649 912 2758 917
rect 2817 912 2846 917
rect 1617 907 1622 912
rect 2841 907 2846 912
rect 2953 912 3254 917
rect 3353 912 3526 917
rect 3601 912 3670 917
rect 3929 912 4342 917
rect 4665 912 4718 917
rect 2953 907 2958 912
rect 697 902 822 907
rect 1161 902 1222 907
rect 1353 902 1478 907
rect 1497 902 1622 907
rect 1665 902 1870 907
rect 1865 897 1870 902
rect 1977 902 2086 907
rect 2353 902 2382 907
rect 1977 897 1982 902
rect 569 892 686 897
rect 1129 892 1246 897
rect 1681 892 1846 897
rect 1865 892 1982 897
rect 2377 897 2382 902
rect 2529 902 2662 907
rect 2841 902 2958 907
rect 3081 902 3182 907
rect 2529 897 2534 902
rect 3177 897 3182 902
rect 3265 902 3366 907
rect 3569 902 3614 907
rect 3785 902 3814 907
rect 3849 902 3942 907
rect 4065 902 4126 907
rect 4217 902 4246 907
rect 3265 897 3270 902
rect 4241 897 4246 902
rect 4329 902 4358 907
rect 4409 902 4454 907
rect 4713 902 4742 907
rect 4329 897 4334 902
rect 2377 892 2534 897
rect 2553 892 2614 897
rect 3137 892 3158 897
rect 3177 892 3270 897
rect 3329 892 3358 897
rect 3369 892 3414 897
rect 3561 892 3638 897
rect 3745 892 3790 897
rect 4241 892 4334 897
rect 1113 882 1406 887
rect 1497 882 1646 887
rect 1825 882 1830 892
rect 3313 882 3342 887
rect 1497 877 1502 882
rect 721 872 846 877
rect 1129 872 1182 877
rect 1225 872 1254 877
rect 1393 872 1502 877
rect 1641 877 1646 882
rect 3337 877 3342 882
rect 3425 882 4102 887
rect 3425 877 3430 882
rect 1641 872 1702 877
rect 2145 872 2222 877
rect 3337 872 3430 877
rect 3505 872 3998 877
rect 4113 872 4198 877
rect 721 867 726 872
rect 697 862 726 867
rect 841 867 846 872
rect 3993 867 4118 872
rect 841 862 1630 867
rect 1625 857 1630 862
rect 1713 862 2254 867
rect 3585 862 3974 867
rect 1713 857 1718 862
rect 233 852 318 857
rect 233 847 238 852
rect 209 842 238 847
rect 313 847 318 852
rect 593 852 678 857
rect 1161 852 1262 857
rect 1417 852 1502 857
rect 1625 852 1718 857
rect 1809 852 1838 857
rect 2265 852 2342 857
rect 3065 852 3206 857
rect 3633 852 3686 857
rect 3977 852 4054 857
rect 593 847 598 852
rect 313 842 342 847
rect 433 842 478 847
rect 529 842 598 847
rect 673 847 678 852
rect 673 842 830 847
rect 1217 842 1358 847
rect 1441 842 1526 847
rect 1785 842 1806 847
rect 1969 842 2046 847
rect 2241 842 2318 847
rect 2753 842 2830 847
rect 1969 837 1974 842
rect 297 832 486 837
rect 609 832 702 837
rect 769 832 806 837
rect 1177 832 1262 837
rect 1273 832 1310 837
rect 1369 832 1726 837
rect 1777 832 1878 837
rect 1945 832 1974 837
rect 2041 837 2046 842
rect 2753 837 2758 842
rect 2041 832 2070 837
rect 2105 832 2222 837
rect 2329 832 2534 837
rect 2729 832 2758 837
rect 2825 837 2830 842
rect 3065 837 3070 852
rect 2825 832 3070 837
rect 3201 837 3206 852
rect 3681 847 3982 852
rect 4049 847 4054 852
rect 4129 852 4158 857
rect 4129 847 4134 852
rect 3337 842 3462 847
rect 3601 842 3662 847
rect 4049 842 4134 847
rect 3201 832 3230 837
rect 1305 827 1374 832
rect 2217 827 2334 832
rect 3337 827 3342 842
rect 201 822 246 827
rect 305 822 334 827
rect 329 817 334 822
rect 433 822 462 827
rect 633 822 678 827
rect 737 822 814 827
rect 865 822 918 827
rect 1233 822 1286 827
rect 1449 822 1534 827
rect 1641 822 1670 827
rect 1785 822 1822 827
rect 1833 822 2078 827
rect 2137 822 2174 827
rect 2537 822 2566 827
rect 2673 822 2718 827
rect 433 817 438 822
rect 1121 817 1214 822
rect 2713 817 2718 822
rect 2833 822 2878 827
rect 3081 822 3118 827
rect 3209 822 3302 827
rect 3313 822 3342 827
rect 3457 827 3462 842
rect 3481 832 4030 837
rect 4497 832 4574 837
rect 3457 822 3566 827
rect 3641 822 3678 827
rect 4481 822 4534 827
rect 4625 822 4654 827
rect 2833 817 2838 822
rect 3297 817 3302 822
rect 3697 817 3822 822
rect 329 812 438 817
rect 593 812 750 817
rect 1097 812 1126 817
rect 1209 812 1230 817
rect 1297 812 1438 817
rect 1545 812 1694 817
rect 1705 812 1870 817
rect 2057 812 2150 817
rect 2161 812 2230 817
rect 2273 812 2334 817
rect 2465 812 2494 817
rect 2713 812 2838 817
rect 3057 812 3094 817
rect 3105 812 3182 817
rect 3297 812 3446 817
rect 3649 812 3702 817
rect 3817 812 3878 817
rect 1225 807 1302 812
rect 1433 807 1550 812
rect 1865 807 2062 812
rect 3441 807 3518 812
rect 3649 807 3654 812
rect 3873 807 3878 812
rect 4041 812 4222 817
rect 4305 812 4382 817
rect 4545 812 4582 817
rect 4041 807 4046 812
rect 625 802 1006 807
rect 1113 802 1198 807
rect 1825 802 1846 807
rect 2081 802 2166 807
rect 2337 802 2486 807
rect 3097 802 3126 807
rect 3513 802 3654 807
rect 3673 802 3694 807
rect 3745 802 3806 807
rect 3873 802 4046 807
rect 4297 802 4326 807
rect 4353 802 4406 807
rect 4481 802 4502 807
rect 4649 802 4678 807
rect 1825 797 1830 802
rect 3161 797 3270 802
rect 193 792 254 797
rect 561 792 678 797
rect 713 792 790 797
rect 1041 792 1286 797
rect 1473 792 1502 797
rect 1729 792 1830 797
rect 1897 792 2062 797
rect 2449 792 2478 797
rect 2857 792 2934 797
rect 2953 792 3014 797
rect 3081 792 3166 797
rect 3265 792 3294 797
rect 3329 792 3494 797
rect 3737 792 3854 797
rect 4177 792 4206 797
rect 4289 792 4334 797
rect 4545 792 4678 797
rect 809 787 958 792
rect 2857 787 2862 792
rect 217 782 262 787
rect 281 782 366 787
rect 465 782 638 787
rect 761 782 814 787
rect 953 782 982 787
rect 1049 782 1086 787
rect 1241 782 1302 787
rect 1321 782 1454 787
rect 1505 782 1526 787
rect 1545 782 1654 787
rect 1673 782 1966 787
rect 2145 782 2198 787
rect 2225 782 2326 787
rect 281 777 286 782
rect 145 772 286 777
rect 361 777 366 782
rect 1113 777 1222 782
rect 1321 777 1326 782
rect 361 772 414 777
rect 537 772 582 777
rect 689 772 1078 777
rect 1089 772 1118 777
rect 1217 772 1326 777
rect 1449 777 1454 782
rect 1545 777 1550 782
rect 1449 772 1550 777
rect 1649 777 1654 782
rect 2193 777 2198 782
rect 2321 777 2326 782
rect 2441 782 2718 787
rect 2833 782 2862 787
rect 2929 787 2934 792
rect 2929 782 2998 787
rect 3065 782 3102 787
rect 3177 782 3374 787
rect 3457 782 3486 787
rect 3649 782 3718 787
rect 3737 782 3782 787
rect 4185 782 4206 787
rect 4273 782 4318 787
rect 2441 777 2446 782
rect 3369 777 3462 782
rect 3649 777 3654 782
rect 1649 772 1838 777
rect 2193 772 2254 777
rect 2321 772 2446 777
rect 2697 772 2758 777
rect 2873 772 2918 777
rect 1089 767 1094 772
rect 2913 767 2918 772
rect 3009 772 3182 777
rect 3257 772 3350 777
rect 3513 772 3582 777
rect 3625 772 3654 777
rect 3713 777 3718 782
rect 3713 772 3758 777
rect 3009 767 3014 772
rect 3513 767 3518 772
rect 417 762 494 767
rect 825 762 942 767
rect 1049 762 1094 767
rect 1129 762 1342 767
rect 1369 762 1422 767
rect 1609 762 1662 767
rect 1873 762 1958 767
rect 2745 762 2774 767
rect 2913 762 3014 767
rect 3057 762 3094 767
rect 3161 762 3342 767
rect 3417 762 3518 767
rect 3577 767 3582 772
rect 3577 762 3606 767
rect 3769 762 3902 767
rect 937 757 1054 762
rect 1441 757 1542 762
rect 3601 757 3774 762
rect 273 752 350 757
rect 545 752 590 757
rect 777 752 918 757
rect 1073 752 1446 757
rect 1537 752 1598 757
rect 1633 752 1742 757
rect 3041 752 3190 757
rect 3201 752 3254 757
rect 4273 752 4310 757
rect 4337 752 4382 757
rect 4537 752 4614 757
rect 273 747 278 752
rect 3041 747 3046 752
rect 161 742 278 747
rect 289 742 318 747
rect 337 742 390 747
rect 449 742 662 747
rect 793 742 814 747
rect 961 742 998 747
rect 1089 742 1134 747
rect 1193 742 1246 747
rect 1321 742 1350 747
rect 1345 737 1350 742
rect 1449 742 1526 747
rect 1993 742 2014 747
rect 2201 742 2318 747
rect 2361 742 2462 747
rect 2809 742 3046 747
rect 3065 742 3222 747
rect 3241 742 3422 747
rect 3481 742 3566 747
rect 3657 742 3702 747
rect 1449 737 1454 742
rect 337 732 1014 737
rect 1185 732 1214 737
rect 1345 732 1454 737
rect 1521 737 1526 742
rect 3217 737 3222 742
rect 3793 737 3798 747
rect 3937 742 3982 747
rect 4089 742 4158 747
rect 4225 742 4334 747
rect 4369 742 4414 747
rect 4505 742 4694 747
rect 1521 732 1542 737
rect 1577 732 1886 737
rect 2521 732 2574 737
rect 3217 732 3246 737
rect 3241 727 3246 732
rect 3377 732 3454 737
rect 3377 727 3382 732
rect 241 722 302 727
rect 393 722 598 727
rect 833 722 854 727
rect 1473 722 1494 727
rect 1825 722 1878 727
rect 1993 722 2102 727
rect 2985 722 3054 727
rect 3241 722 3382 727
rect 3449 727 3454 732
rect 3561 732 3590 737
rect 3681 732 3750 737
rect 3793 732 3894 737
rect 3961 732 4046 737
rect 4249 732 4302 737
rect 3561 727 3566 732
rect 4321 727 4326 737
rect 4657 732 4742 737
rect 3449 722 3566 727
rect 3649 722 4574 727
rect 2873 717 2966 722
rect 129 712 174 717
rect 185 712 214 717
rect 321 712 374 717
rect 401 712 430 717
rect 529 712 574 717
rect 641 712 758 717
rect 801 712 862 717
rect 905 712 950 717
rect 1089 712 1166 717
rect 1529 712 1574 717
rect 1857 712 1950 717
rect 2521 712 2606 717
rect 2849 712 2878 717
rect 2961 712 2998 717
rect 3017 712 3134 717
rect 3193 712 3222 717
rect 3633 712 3654 717
rect 4233 712 4422 717
rect 4441 712 4534 717
rect 4721 712 4758 717
rect 1089 707 1094 712
rect 177 702 358 707
rect 817 702 838 707
rect 849 702 1094 707
rect 1161 707 1166 712
rect 3785 707 3926 712
rect 4417 707 4422 712
rect 1161 702 1462 707
rect 849 697 854 702
rect 1457 697 1462 702
rect 1585 702 1870 707
rect 1897 702 1974 707
rect 2273 702 2382 707
rect 2417 702 2502 707
rect 2553 702 2670 707
rect 2913 702 2942 707
rect 1585 697 1590 702
rect 337 692 398 697
rect 641 692 854 697
rect 873 692 982 697
rect 1105 692 1158 697
rect 1457 692 1590 697
rect 2937 697 2942 702
rect 3017 702 3046 707
rect 3065 702 3118 707
rect 3401 702 3494 707
rect 3521 702 3614 707
rect 3665 702 3790 707
rect 3921 702 4134 707
rect 4417 702 4494 707
rect 4593 702 4702 707
rect 3017 697 3022 702
rect 3401 697 3406 702
rect 2937 692 3022 697
rect 3073 692 3166 697
rect 3377 692 3406 697
rect 3489 697 3494 702
rect 4153 697 4398 702
rect 4513 697 4598 702
rect 4697 697 4702 702
rect 3489 692 3510 697
rect 641 687 646 692
rect 225 682 326 687
rect 409 682 646 687
rect 2145 682 2254 687
rect 321 677 414 682
rect 3505 677 3510 692
rect 3705 692 4158 697
rect 4393 692 4518 697
rect 4697 692 4870 697
rect 3705 677 3710 692
rect 3729 682 4654 687
rect 4713 682 4742 687
rect 2609 672 2806 677
rect 3409 672 3470 677
rect 3505 672 3710 677
rect 3745 672 4494 677
rect 4489 667 4494 672
rect 4577 672 4638 677
rect 4577 667 4582 672
rect 377 662 590 667
rect 377 657 382 662
rect 201 652 382 657
rect 585 657 590 662
rect 665 662 790 667
rect 3745 662 3774 667
rect 4017 662 4038 667
rect 4489 662 4582 667
rect 665 657 670 662
rect 585 652 670 657
rect 785 657 790 662
rect 785 652 1150 657
rect 3057 652 3246 657
rect 393 642 782 647
rect 2233 642 2398 647
rect 3057 637 3062 652
rect 553 632 646 637
rect 1185 632 1214 637
rect 1473 632 1494 637
rect 369 622 750 627
rect 865 622 918 627
rect 1129 622 1214 627
rect 1225 622 1310 627
rect 1481 622 1534 627
rect 1553 622 1710 627
rect 1745 622 1838 627
rect 1553 617 1558 622
rect 161 612 406 617
rect 633 612 742 617
rect 817 612 894 617
rect 1073 612 1558 617
rect 1705 617 1710 622
rect 1705 612 1734 617
rect 1873 612 1918 617
rect 425 607 614 612
rect 305 602 350 607
rect 393 602 430 607
rect 609 602 1006 607
rect 1089 602 1286 607
rect 1657 602 1710 607
rect 1481 597 1566 602
rect 361 592 518 597
rect 569 592 606 597
rect 625 592 694 597
rect 769 592 1038 597
rect 1145 592 1222 597
rect 1321 592 1350 597
rect 1457 592 1486 597
rect 1561 592 1646 597
rect 1713 592 1966 597
rect 225 582 358 587
rect 553 582 590 587
rect 617 582 646 587
rect 889 582 966 587
rect 1017 582 1550 587
rect 665 577 870 582
rect 1545 577 1550 582
rect 1641 582 1742 587
rect 2049 582 2054 637
rect 2329 632 2358 637
rect 3033 632 3062 637
rect 3241 637 3246 652
rect 3241 632 3270 637
rect 3505 632 3582 637
rect 4513 632 4590 637
rect 2537 622 2638 627
rect 2993 622 3046 627
rect 3097 622 3142 627
rect 3265 622 3294 627
rect 3561 622 3590 627
rect 4489 622 4542 627
rect 3049 612 3086 617
rect 3169 612 3230 617
rect 3465 612 3502 617
rect 3521 612 3558 617
rect 2345 602 2374 607
rect 3929 602 4030 607
rect 4305 602 4334 607
rect 4377 602 4446 607
rect 3049 597 3126 602
rect 2353 592 2478 597
rect 2513 592 2630 597
rect 2817 592 2862 597
rect 3025 592 3054 597
rect 3121 592 3254 597
rect 3329 592 3462 597
rect 3497 592 3534 597
rect 3817 592 3878 597
rect 4153 592 4198 597
rect 4281 592 4358 597
rect 4417 592 4550 597
rect 4561 592 4686 597
rect 4721 592 4758 597
rect 2513 587 2518 592
rect 2361 582 2406 587
rect 2425 582 2518 587
rect 2625 587 2630 592
rect 4545 587 4550 592
rect 2625 582 2758 587
rect 3081 582 3110 587
rect 3225 582 3350 587
rect 3761 582 3830 587
rect 4081 582 4166 587
rect 4449 582 4526 587
rect 4545 582 4582 587
rect 4609 582 4646 587
rect 1641 577 1646 582
rect 2401 577 2406 582
rect 81 572 230 577
rect 225 567 230 572
rect 401 572 430 577
rect 545 572 670 577
rect 865 572 982 577
rect 1113 572 1166 577
rect 1193 572 1334 577
rect 1545 572 1646 577
rect 2137 572 2182 577
rect 2401 572 2454 577
rect 401 567 406 572
rect 1377 567 1502 572
rect 2449 567 2454 572
rect 2529 572 2614 577
rect 3073 572 3110 577
rect 3601 572 3742 577
rect 2529 567 2534 572
rect 225 562 406 567
rect 577 562 990 567
rect 1305 562 1382 567
rect 1497 562 1526 567
rect 1985 562 2046 567
rect 2073 562 2102 567
rect 2217 562 2246 567
rect 2449 562 2534 567
rect 2097 557 2222 562
rect 3601 557 3606 572
rect 185 552 206 557
rect 593 552 630 557
rect 753 552 862 557
rect 897 552 1094 557
rect 1113 552 1286 557
rect 1393 552 1542 557
rect 1561 552 1638 557
rect 2897 552 3086 557
rect 3577 552 3606 557
rect 3737 557 3742 572
rect 3849 562 4062 567
rect 4145 562 4366 567
rect 4561 562 4694 567
rect 3849 557 3854 562
rect 3737 552 3854 557
rect 4057 557 4062 562
rect 4057 552 4238 557
rect 753 547 758 552
rect 1113 547 1118 552
rect 1281 547 1374 552
rect 1561 547 1566 552
rect 441 542 566 547
rect 633 542 758 547
rect 769 542 1006 547
rect 1033 542 1118 547
rect 1369 542 1566 547
rect 1633 547 1638 552
rect 4233 547 4238 552
rect 4313 552 4510 557
rect 4521 552 4590 557
rect 4625 552 4662 557
rect 4313 547 4318 552
rect 1633 542 1662 547
rect 2121 542 2166 547
rect 2273 542 2318 547
rect 2553 542 2846 547
rect 3073 542 3238 547
rect 3553 542 3590 547
rect 3673 542 3766 547
rect 3977 542 4046 547
rect 4089 542 4214 547
rect 4233 542 4318 547
rect 4385 542 4750 547
rect 1137 537 1254 542
rect 377 532 478 537
rect 745 532 870 537
rect 993 532 1142 537
rect 1249 532 1278 537
rect 1329 532 1446 537
rect 1649 532 1750 537
rect 2705 532 2734 537
rect 329 522 518 527
rect 649 522 702 527
rect 849 522 918 527
rect 1065 522 1142 527
rect 1185 522 1846 527
rect 1945 522 1966 527
rect 1841 517 1846 522
rect 2729 517 2734 532
rect 2857 532 2926 537
rect 3241 532 3326 537
rect 3681 532 3846 537
rect 3865 532 3942 537
rect 4617 532 4646 537
rect 2857 517 2862 532
rect 4641 527 4646 532
rect 2929 522 2958 527
rect 3577 522 3654 527
rect 3713 522 3862 527
rect 3889 522 4110 527
rect 4625 522 4646 527
rect 3577 517 3582 522
rect 241 512 422 517
rect 561 512 742 517
rect 777 512 838 517
rect 833 507 838 512
rect 897 512 926 517
rect 1153 512 1222 517
rect 1297 512 1718 517
rect 1729 512 1830 517
rect 1841 512 1974 517
rect 2729 512 2862 517
rect 3017 512 3254 517
rect 3505 512 3582 517
rect 897 507 902 512
rect 1729 507 1734 512
rect 3649 507 3654 522
rect 3809 512 3846 517
rect 4025 512 4094 517
rect 4577 512 4638 517
rect 4681 512 4742 517
rect 233 502 430 507
rect 473 502 502 507
rect 497 497 502 502
rect 577 502 702 507
rect 833 502 902 507
rect 937 502 1286 507
rect 577 497 582 502
rect 209 492 398 497
rect 497 492 582 497
rect 633 492 678 497
rect 697 487 702 502
rect 937 487 942 502
rect 1281 497 1286 502
rect 1353 502 1406 507
rect 1353 497 1358 502
rect 1281 492 1358 497
rect 1401 497 1406 502
rect 1481 502 1526 507
rect 1713 502 1734 507
rect 1793 502 1854 507
rect 3241 502 3366 507
rect 3593 502 3630 507
rect 3649 502 3870 507
rect 1481 497 1486 502
rect 1401 492 1486 497
rect 1521 497 1526 502
rect 1521 492 1702 497
rect 1777 492 1862 497
rect 3457 492 3494 497
rect 1697 487 1782 492
rect 3489 487 3494 492
rect 3881 492 4102 497
rect 3881 487 3886 492
rect 697 482 942 487
rect 1969 482 2118 487
rect 3489 482 3886 487
rect 393 472 462 477
rect 1049 472 1270 477
rect 1305 472 1550 477
rect 1545 467 1550 472
rect 1641 472 1670 477
rect 1681 472 1998 477
rect 4537 472 4622 477
rect 1641 467 1646 472
rect 1545 462 1646 467
rect 2017 462 2150 467
rect 4457 462 4502 467
rect 1889 457 2022 462
rect 2145 457 2150 462
rect 689 452 838 457
rect 409 442 598 447
rect 409 437 414 442
rect 385 432 414 437
rect 593 437 598 442
rect 689 437 694 452
rect 593 432 694 437
rect 833 437 838 452
rect 881 452 1030 457
rect 1865 452 1894 457
rect 2145 452 2174 457
rect 3457 452 4006 457
rect 881 447 886 452
rect 857 442 886 447
rect 1025 447 1030 452
rect 1025 442 1238 447
rect 1745 442 1814 447
rect 1857 442 2286 447
rect 3681 442 3710 447
rect 3969 442 3990 447
rect 4097 442 4206 447
rect 4281 442 4366 447
rect 1745 437 1750 442
rect 833 432 862 437
rect 937 432 990 437
rect 1721 432 1750 437
rect 1809 437 1814 442
rect 4097 437 4102 442
rect 1809 432 1910 437
rect 2001 432 2078 437
rect 4073 432 4102 437
rect 4201 437 4206 442
rect 4201 432 4270 437
rect 4265 427 4270 432
rect 4369 432 4430 437
rect 4369 427 4374 432
rect 129 422 174 427
rect 193 422 230 427
rect 273 422 334 427
rect 433 422 510 427
rect 433 417 438 422
rect 209 412 238 417
rect 369 412 398 417
rect 409 412 438 417
rect 505 417 510 422
rect 593 417 598 427
rect 705 422 750 427
rect 801 422 886 427
rect 977 422 1022 427
rect 1329 422 1454 427
rect 1601 422 1646 427
rect 1657 422 1702 427
rect 1897 422 1918 427
rect 1929 422 2014 427
rect 2065 422 2110 427
rect 2553 422 2582 427
rect 2705 422 2934 427
rect 2945 422 2998 427
rect 3065 422 3134 427
rect 3313 422 3430 427
rect 3665 422 3702 427
rect 3713 422 3734 427
rect 4153 422 4190 427
rect 4265 422 4374 427
rect 4393 422 4438 427
rect 505 412 598 417
rect 665 412 798 417
rect 913 412 958 417
rect 1145 412 1310 417
rect 1689 412 1798 417
rect 2561 412 2606 417
rect 3521 412 3574 417
rect 3649 412 3678 417
rect 233 407 374 412
rect 1145 407 1150 412
rect 417 402 598 407
rect 1121 402 1150 407
rect 1305 407 1310 412
rect 1529 407 1622 412
rect 1873 407 1950 412
rect 3745 407 3750 417
rect 3841 412 4062 417
rect 4105 412 4150 417
rect 1305 402 1398 407
rect 169 392 278 397
rect 273 387 278 392
rect 417 387 422 402
rect 1393 397 1398 402
rect 1465 402 1534 407
rect 1617 402 1646 407
rect 1665 402 1734 407
rect 1809 402 1878 407
rect 1945 402 1974 407
rect 2801 402 2846 407
rect 3505 402 3790 407
rect 4273 402 4318 407
rect 4497 402 4574 407
rect 1465 397 1470 402
rect 1729 397 1814 402
rect 4497 397 4502 402
rect 441 392 478 397
rect 697 392 726 397
rect 1137 392 1374 397
rect 1393 392 1470 397
rect 1545 392 1710 397
rect 1889 392 1966 397
rect 1985 392 2182 397
rect 2257 392 2438 397
rect 2465 392 2526 397
rect 2585 392 2622 397
rect 2657 392 3030 397
rect 3433 392 3470 397
rect 3529 392 3598 397
rect 3657 392 3894 397
rect 4065 392 4182 397
rect 4233 392 4502 397
rect 4569 397 4574 402
rect 4569 392 4702 397
rect 81 382 158 387
rect 153 377 158 382
rect 225 382 254 387
rect 273 382 422 387
rect 585 382 1086 387
rect 1129 382 1158 387
rect 225 377 230 382
rect 153 372 230 377
rect 1153 377 1158 382
rect 1225 382 1262 387
rect 1625 382 1654 387
rect 1225 377 1230 382
rect 1153 372 1230 377
rect 1649 377 1654 382
rect 1817 382 1886 387
rect 1969 382 1998 387
rect 1817 377 1822 382
rect 1649 372 1822 377
rect 1993 377 1998 382
rect 2193 382 2246 387
rect 2369 382 2414 387
rect 2193 377 2198 382
rect 1993 372 2198 377
rect 2409 377 2414 382
rect 2481 382 2510 387
rect 2481 377 2486 382
rect 4041 377 4302 382
rect 2409 372 2486 377
rect 3049 372 3150 377
rect 3593 372 4046 377
rect 4297 372 4638 377
rect 3049 367 3054 372
rect 873 362 1054 367
rect 1313 362 1342 367
rect 2361 362 2390 367
rect 2537 362 2630 367
rect 3025 362 3054 367
rect 3145 367 3150 372
rect 3145 362 3342 367
rect 4057 362 4294 367
rect 873 357 878 362
rect 553 352 878 357
rect 1049 357 1054 362
rect 2537 357 2542 362
rect 1049 352 1078 357
rect 1249 352 1438 357
rect 1945 352 2054 357
rect 2145 352 2190 357
rect 2441 352 2542 357
rect 2625 357 2630 362
rect 2625 352 2654 357
rect 3121 352 3198 357
rect 3417 352 3510 357
rect 4025 352 4150 357
rect 4161 352 4246 357
rect 329 342 550 347
rect 889 342 1062 347
rect 1321 342 1382 347
rect 1473 342 1614 347
rect 1633 342 1702 347
rect 1745 342 1774 347
rect 2041 342 2198 347
rect 2553 342 2582 347
rect 1633 337 1638 342
rect 201 332 374 337
rect 545 332 566 337
rect 1073 332 1110 337
rect 1145 332 1350 337
rect 1505 332 1638 337
rect 1697 337 1702 342
rect 2577 337 2582 342
rect 2665 342 2822 347
rect 2841 342 3006 347
rect 3049 342 3126 347
rect 3209 342 3310 347
rect 3657 342 3846 347
rect 3969 342 4078 347
rect 4105 342 4198 347
rect 4257 342 4462 347
rect 4617 342 4710 347
rect 2665 337 2670 342
rect 2841 337 2846 342
rect 1697 332 1726 337
rect 1793 332 1926 337
rect 2577 332 2670 337
rect 2793 332 2846 337
rect 3001 337 3006 342
rect 3121 337 3214 342
rect 4193 337 4262 342
rect 3001 332 3054 337
rect 3321 332 3414 337
rect 3497 332 3614 337
rect 3825 332 3878 337
rect 3889 332 4174 337
rect 4609 332 4638 337
rect 4721 332 4750 337
rect 873 327 1030 332
rect 1393 327 1486 332
rect 1793 327 1798 332
rect 849 322 878 327
rect 1025 322 1062 327
rect 1137 322 1166 327
rect 1369 322 1398 327
rect 1481 322 1518 327
rect 1673 322 1798 327
rect 1921 327 1926 332
rect 3049 327 3054 332
rect 3241 327 3326 332
rect 3641 327 3806 332
rect 3889 327 3894 332
rect 4633 327 4726 332
rect 1921 322 2110 327
rect 2129 322 2182 327
rect 3049 322 3246 327
rect 3417 322 3646 327
rect 3801 322 3894 327
rect 3929 322 4030 327
rect 4041 322 4102 327
rect 4193 322 4390 327
rect 1057 317 1142 322
rect 4193 317 4198 322
rect 137 312 182 317
rect 297 312 342 317
rect 385 312 494 317
rect 561 312 582 317
rect 681 312 726 317
rect 737 312 950 317
rect 969 312 1014 317
rect 1201 312 1262 317
rect 1361 312 1686 317
rect 1745 312 1910 317
rect 2033 312 2086 317
rect 2153 312 2198 317
rect 2233 312 2262 317
rect 2361 312 2406 317
rect 2817 312 3030 317
rect 3265 312 3446 317
rect 3481 312 3510 317
rect 3657 312 3838 317
rect 3953 312 4198 317
rect 4385 317 4390 322
rect 4385 312 4566 317
rect 4641 312 4774 317
rect 1905 307 2038 312
rect 2081 307 2086 312
rect 3505 307 3662 312
rect 3833 307 3958 312
rect 4217 307 4350 312
rect 177 302 206 307
rect 201 287 206 302
rect 465 302 574 307
rect 929 302 982 307
rect 1121 302 1694 307
rect 2081 302 2238 307
rect 2409 302 2678 307
rect 3417 302 3470 307
rect 3785 302 3814 307
rect 465 297 470 302
rect 3809 297 3814 302
rect 3977 302 4222 307
rect 4345 302 4374 307
rect 3977 297 3982 302
rect 345 292 470 297
rect 713 292 910 297
rect 945 292 1110 297
rect 1345 292 1502 297
rect 1625 292 1726 297
rect 345 287 350 292
rect 713 287 718 292
rect 201 282 350 287
rect 489 282 718 287
rect 905 287 910 292
rect 1105 287 1350 292
rect 1721 287 1726 292
rect 1817 292 2006 297
rect 2161 292 2214 297
rect 3057 292 3254 297
rect 1817 287 1822 292
rect 3249 287 3254 292
rect 3561 292 3646 297
rect 3809 292 3982 297
rect 4001 292 4030 297
rect 4145 292 4670 297
rect 3561 287 3566 292
rect 4025 287 4150 292
rect 905 282 974 287
rect 1721 282 1822 287
rect 2577 282 2606 287
rect 1369 277 1486 282
rect 2601 277 2606 282
rect 2689 282 3046 287
rect 3249 282 3566 287
rect 4169 282 4318 287
rect 2689 277 2694 282
rect 393 272 470 277
rect 729 272 894 277
rect 985 272 1142 277
rect 1249 272 1374 277
rect 1481 272 1702 277
rect 2601 272 2694 277
rect 3857 272 4206 277
rect 393 267 398 272
rect 369 262 398 267
rect 465 267 470 272
rect 889 267 990 272
rect 4201 267 4206 272
rect 4585 272 4614 277
rect 4585 267 4590 272
rect 465 262 742 267
rect 1193 262 1470 267
rect 1841 262 1974 267
rect 4201 262 4590 267
rect 561 252 742 257
rect 825 252 934 257
rect 1153 252 1374 257
rect 1721 252 1798 257
rect 1721 247 1726 252
rect 225 242 622 247
rect 969 242 1198 247
rect 1209 242 1254 247
rect 1465 242 1726 247
rect 1793 247 1798 252
rect 1841 247 1846 262
rect 1793 242 1846 247
rect 1969 247 1974 262
rect 3137 252 3486 257
rect 3137 247 3142 252
rect 1969 242 2070 247
rect 2737 242 2846 247
rect 3065 242 3142 247
rect 3481 247 3486 252
rect 3633 252 3838 257
rect 3633 247 3638 252
rect 3481 242 3534 247
rect 3553 242 3638 247
rect 3833 247 3838 252
rect 3833 242 3950 247
rect 4009 242 4046 247
rect 4121 242 4182 247
rect 2737 237 2742 242
rect 121 232 374 237
rect 521 232 678 237
rect 745 232 862 237
rect 1097 232 1158 237
rect 1201 232 1342 237
rect 1433 232 1494 237
rect 1777 232 1958 237
rect 2617 232 2702 237
rect 2713 232 2742 237
rect 2841 237 2846 242
rect 3553 237 3558 242
rect 2841 232 2870 237
rect 3153 232 3238 237
rect 3473 232 3558 237
rect 3945 237 3950 242
rect 3945 232 3974 237
rect 4297 232 4334 237
rect 1201 227 1206 232
rect 169 222 270 227
rect 297 222 334 227
rect 353 222 422 227
rect 457 222 510 227
rect 545 222 838 227
rect 921 222 966 227
rect 985 222 1078 227
rect 1129 222 1206 227
rect 1233 222 1366 227
rect 1401 222 1518 227
rect 1665 222 1758 227
rect 1921 222 2014 227
rect 2409 222 2518 227
rect 2681 222 2782 227
rect 2913 222 2942 227
rect 3193 222 3414 227
rect 3649 222 3694 227
rect 3753 222 3790 227
rect 3841 222 3878 227
rect 3953 222 3990 227
rect 4089 222 4166 227
rect 4249 222 4366 227
rect 4409 222 4446 227
rect 4465 222 4494 227
rect 4601 222 4774 227
rect 985 217 990 222
rect 161 212 182 217
rect 209 212 246 217
rect 321 212 382 217
rect 393 212 534 217
rect 665 212 710 217
rect 809 212 990 217
rect 1073 217 1078 222
rect 1073 212 1118 217
rect 1169 212 1246 217
rect 1353 212 1390 217
rect 1409 212 1430 217
rect 1505 212 1582 217
rect 1761 212 1830 217
rect 1945 207 1950 217
rect 2057 212 2078 217
rect 2833 212 2982 217
rect 3497 212 3526 217
rect 3569 212 3662 217
rect 3673 212 4174 217
rect 4201 212 4230 217
rect 4441 212 4470 217
rect 4593 212 4662 217
rect 4225 207 4446 212
rect 481 202 558 207
rect 625 202 926 207
rect 625 197 630 202
rect 921 197 926 202
rect 993 202 1022 207
rect 1081 202 1654 207
rect 1713 202 1774 207
rect 1801 202 1886 207
rect 1945 202 2054 207
rect 2273 202 2366 207
rect 2649 202 2774 207
rect 2793 202 2854 207
rect 3489 202 3518 207
rect 993 197 998 202
rect 3513 197 3518 202
rect 3601 202 3654 207
rect 4105 202 4166 207
rect 3601 197 3606 202
rect 377 192 526 197
rect 545 192 630 197
rect 641 192 758 197
rect 873 192 902 197
rect 921 192 998 197
rect 1153 192 1206 197
rect 1321 192 1382 197
rect 1497 192 1518 197
rect 1633 192 1686 197
rect 1745 192 1814 197
rect 2209 192 2494 197
rect 2761 192 2806 197
rect 2841 192 2886 197
rect 2921 192 3006 197
rect 3105 192 3286 197
rect 3305 192 3470 197
rect 3513 192 3606 197
rect 3625 192 4150 197
rect 4185 192 4246 197
rect 4321 192 4598 197
rect 4609 192 4702 197
rect 257 182 366 187
rect 361 177 366 182
rect 473 182 566 187
rect 817 182 838 187
rect 1233 182 1510 187
rect 1673 182 1870 187
rect 2065 182 2198 187
rect 473 177 478 182
rect 817 177 822 182
rect 2193 177 2198 182
rect 2273 182 2374 187
rect 2721 182 2910 187
rect 2977 182 3318 187
rect 4289 182 4366 187
rect 4465 182 4518 187
rect 4649 182 4678 187
rect 2273 177 2278 182
rect 4513 177 4654 182
rect 361 172 478 177
rect 513 172 822 177
rect 1137 172 1326 177
rect 1321 167 1326 172
rect 1385 172 1438 177
rect 1385 167 1390 172
rect 497 162 654 167
rect 809 162 886 167
rect 1241 162 1270 167
rect 1321 162 1390 167
rect 1433 167 1438 172
rect 1521 172 1662 177
rect 1521 167 1526 172
rect 1433 162 1526 167
rect 1657 167 1662 172
rect 1753 172 1782 177
rect 2193 172 2278 177
rect 2297 172 2334 177
rect 2721 172 2750 177
rect 1753 167 1758 172
rect 1657 162 1758 167
rect 2745 167 2750 172
rect 2873 172 3158 177
rect 2873 167 2878 172
rect 3153 167 3158 172
rect 3233 172 3630 177
rect 4001 172 4030 177
rect 4137 172 4206 177
rect 3233 167 3238 172
rect 4137 167 4142 172
rect 2745 162 2878 167
rect 2993 162 3110 167
rect 3153 162 3238 167
rect 3257 162 3302 167
rect 3649 162 4142 167
rect 4201 167 4206 172
rect 4201 162 4278 167
rect 1985 157 2054 162
rect 833 152 1014 157
rect 1073 152 1302 157
rect 1961 152 1990 157
rect 2049 152 2166 157
rect 2585 152 2622 157
rect 2897 152 2958 157
rect 3105 147 3110 162
rect 3257 147 3262 162
rect 4273 157 4278 162
rect 4377 162 4454 167
rect 4377 157 4382 162
rect 4153 152 4190 157
rect 4273 152 4382 157
rect 4449 157 4454 162
rect 4513 162 4726 167
rect 4513 157 4518 162
rect 4449 152 4518 157
rect 4577 152 4606 157
rect 81 142 182 147
rect 297 142 414 147
rect 529 142 694 147
rect 745 142 854 147
rect 1049 142 1110 147
rect 1481 142 1606 147
rect 1713 142 1870 147
rect 2009 142 2038 147
rect 2033 137 2038 142
rect 2105 142 2134 147
rect 2105 137 2110 142
rect 873 132 918 137
rect 2033 132 2110 137
rect 2225 127 2230 147
rect 2241 142 2278 147
rect 2289 142 2326 147
rect 2585 142 2638 147
rect 2697 142 2726 147
rect 2769 142 2830 147
rect 2897 142 2942 147
rect 2969 142 3006 147
rect 3105 142 3262 147
rect 3281 142 3422 147
rect 3569 142 3646 147
rect 4537 142 4574 147
rect 4641 142 4710 147
rect 2273 127 2278 142
rect 2833 132 2886 137
rect 2921 132 2950 137
rect 3017 132 3086 137
rect 2945 127 3022 132
rect 617 122 646 127
rect 641 117 646 122
rect 873 122 1142 127
rect 2225 122 2246 127
rect 2273 122 2294 127
rect 2865 122 2918 127
rect 3625 122 4390 127
rect 873 117 878 122
rect 641 112 878 117
rect 1057 112 1102 117
rect 1689 112 1734 117
rect 1841 112 1886 117
rect 2273 112 2318 117
rect 2393 112 2518 117
rect 2601 112 2654 117
rect 2873 112 2990 117
rect 3257 112 3446 117
rect 3817 112 3870 117
rect 4649 112 4774 117
rect 2889 102 2918 107
rect 2913 97 2918 102
rect 3001 102 3150 107
rect 3001 97 3006 102
rect 2089 92 2118 97
rect 2161 92 2262 97
rect 2257 87 2262 92
rect 2329 92 2422 97
rect 2913 92 3006 97
rect 3601 92 3646 97
rect 2329 87 2334 92
rect 2025 82 2094 87
rect 2257 82 2334 87
rect 4113 72 4142 77
rect 3713 62 3750 67
rect 2169 32 2230 37
rect 2465 12 2726 17
rect 3889 12 3918 17
rect 3961 12 4030 17
rect 4065 12 4102 17
rect 4209 12 4246 17
use M3_M2  M3_M2_0
timestamp 1677622389
transform 1 0 1684 0 1 4735
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1677622389
transform 1 0 3252 0 1 4735
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_0
timestamp 1677622389
transform 1 0 24 0 1 4717
box -10 -10 10 10
use M3_M2  M3_M2_2
timestamp 1677622389
transform 1 0 1940 0 1 4725
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1677622389
transform 1 0 2644 0 1 4725
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_1
timestamp 1677622389
transform 1 0 4843 0 1 4717
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_2
timestamp 1677622389
transform 1 0 48 0 1 4693
box -10 -10 10 10
use M3_M2  M3_M2_4
timestamp 1677622389
transform 1 0 1148 0 1 4685
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1677622389
transform 1 0 2836 0 1 4685
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_3
timestamp 1677622389
transform 1 0 4819 0 1 4693
box -10 -10 10 10
use top_level_VIA0  top_level_VIA0_0
timestamp 1677622389
transform 1 0 24 0 1 4670
box -10 -3 10 3
use M2_M1  M2_M1_3
timestamp 1677622389
transform 1 0 116 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1677622389
transform 1 0 172 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1677622389
transform 1 0 92 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_74
timestamp 1677622389
transform 1 0 92 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1677622389
transform 1 0 244 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1677622389
transform 1 0 284 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1677622389
transform 1 0 244 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1677622389
transform 1 0 284 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1677622389
transform 1 0 340 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1677622389
transform 1 0 236 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1677622389
transform 1 0 260 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1677622389
transform 1 0 260 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1677622389
transform 1 0 276 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1677622389
transform 1 0 388 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1677622389
transform 1 0 428 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_8
timestamp 1677622389
transform 1 0 388 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_34
timestamp 1677622389
transform 1 0 404 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1677622389
transform 1 0 428 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1677622389
transform 1 0 484 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1677622389
transform 1 0 380 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1677622389
transform 1 0 404 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1677622389
transform 1 0 380 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1677622389
transform 1 0 404 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1677622389
transform 1 0 532 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1677622389
transform 1 0 588 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1677622389
transform 1 0 508 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1677622389
transform 1 0 508 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1677622389
transform 1 0 660 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1677622389
transform 1 0 700 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1677622389
transform 1 0 660 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1677622389
transform 1 0 692 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1677622389
transform 1 0 700 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1677622389
transform 1 0 612 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1677622389
transform 1 0 700 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1677622389
transform 1 0 612 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1677622389
transform 1 0 716 0 1 4615
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1677622389
transform 1 0 812 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1677622389
transform 1 0 852 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1677622389
transform 1 0 812 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1677622389
transform 1 0 844 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1677622389
transform 1 0 852 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1677622389
transform 1 0 764 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1677622389
transform 1 0 852 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1677622389
transform 1 0 868 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_115
timestamp 1677622389
transform 1 0 844 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1677622389
transform 1 0 860 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1677622389
transform 1 0 940 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_81
timestamp 1677622389
transform 1 0 940 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_98
timestamp 1677622389
transform 1 0 964 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_82
timestamp 1677622389
transform 1 0 964 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_0
timestamp 1677622389
transform 1 0 980 0 1 4625
box -2 -2 2 2
use M3_M2  M3_M2_12
timestamp 1677622389
transform 1 0 1076 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1677622389
transform 1 0 1044 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1677622389
transform 1 0 1084 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1677622389
transform 1 0 1044 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1677622389
transform 1 0 1076 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1677622389
transform 1 0 1084 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1677622389
transform 1 0 996 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_83
timestamp 1677622389
transform 1 0 996 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1677622389
transform 1 0 1132 0 1 4645
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1677622389
transform 1 0 1108 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1677622389
transform 1 0 1132 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1677622389
transform 1 0 1092 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1677622389
transform 1 0 1116 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_36
timestamp 1677622389
transform 1 0 1124 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_25
timestamp 1677622389
transform 1 0 1132 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1677622389
transform 1 0 1092 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_100
timestamp 1677622389
transform 1 0 1100 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1677622389
transform 1 0 1108 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1677622389
transform 1 0 1124 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1677622389
transform 1 0 1132 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1677622389
transform 1 0 1140 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1677622389
transform 1 0 1156 0 1 4615
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1677622389
transform 1 0 1172 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1677622389
transform 1 0 1180 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1677622389
transform 1 0 1220 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_26
timestamp 1677622389
transform 1 0 1180 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1677622389
transform 1 0 1188 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1677622389
transform 1 0 1220 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1677622389
transform 1 0 1268 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1677622389
transform 1 0 1268 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1677622389
transform 1 0 1356 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1677622389
transform 1 0 1388 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1677622389
transform 1 0 1308 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1677622389
transform 1 0 1356 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1677622389
transform 1 0 1308 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1677622389
transform 1 0 1404 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_31
timestamp 1677622389
transform 1 0 1468 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1677622389
transform 1 0 1420 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1677622389
transform 1 0 1468 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1677622389
transform 1 0 1420 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1677622389
transform 1 0 1444 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1677622389
transform 1 0 1508 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_32
timestamp 1677622389
transform 1 0 1524 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1677622389
transform 1 0 1612 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1677622389
transform 1 0 1660 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1677622389
transform 1 0 1668 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1677622389
transform 1 0 1580 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1677622389
transform 1 0 1652 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1677622389
transform 1 0 1580 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1677622389
transform 1 0 1668 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1677622389
transform 1 0 1732 0 1 4645
box -3 -3 3 3
use M2_M1  M2_M1_108
timestamp 1677622389
transform 1 0 1732 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_10
timestamp 1677622389
transform 1 0 1796 0 1 4645
box -3 -3 3 3
use M2_M1  M2_M1_36
timestamp 1677622389
transform 1 0 1796 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_28
timestamp 1677622389
transform 1 0 1860 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1677622389
transform 1 0 1900 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1677622389
transform 1 0 1860 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1677622389
transform 1 0 1892 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1677622389
transform 1 0 1900 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1677622389
transform 1 0 1812 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1677622389
transform 1 0 1812 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_110
timestamp 1677622389
transform 1 0 1900 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_30
timestamp 1677622389
transform 1 0 1924 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1677622389
transform 1 0 2004 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1677622389
transform 1 0 2036 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1677622389
transform 1 0 2044 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1677622389
transform 1 0 1956 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1677622389
transform 1 0 2004 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1677622389
transform 1 0 1956 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1677622389
transform 1 0 1996 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1677622389
transform 1 0 2044 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_112
timestamp 1677622389
transform 1 0 2068 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1677622389
transform 1 0 2108 0 1 4665
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1677622389
transform 1 0 2188 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1677622389
transform 1 0 2220 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1677622389
transform 1 0 2228 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1677622389
transform 1 0 2140 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1677622389
transform 1 0 2188 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1677622389
transform 1 0 2140 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1677622389
transform 1 0 2172 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1677622389
transform 1 0 2228 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_114
timestamp 1677622389
transform 1 0 2236 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1677622389
transform 1 0 2300 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1677622389
transform 1 0 2316 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1677622389
transform 1 0 2324 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1677622389
transform 1 0 2316 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1677622389
transform 1 0 2380 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1677622389
transform 1 0 2380 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_116
timestamp 1677622389
transform 1 0 2428 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_118
timestamp 1677622389
transform 1 0 2396 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_117
timestamp 1677622389
transform 1 0 2532 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1677622389
transform 1 0 2564 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1677622389
transform 1 0 2564 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_50
timestamp 1677622389
transform 1 0 2604 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1677622389
transform 1 0 2660 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1677622389
transform 1 0 2580 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1677622389
transform 1 0 2604 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1677622389
transform 1 0 2580 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1677622389
transform 1 0 2660 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_119
timestamp 1677622389
transform 1 0 2684 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1677622389
transform 1 0 2708 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1677622389
transform 1 0 2708 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1677622389
transform 1 0 2748 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1677622389
transform 1 0 2804 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1677622389
transform 1 0 2724 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1677622389
transform 1 0 2748 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_121
timestamp 1677622389
transform 1 0 2812 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1677622389
transform 1 0 2724 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1677622389
transform 1 0 2804 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1677622389
transform 1 0 2812 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_55
timestamp 1677622389
transform 1 0 2836 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1677622389
transform 1 0 2852 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1677622389
transform 1 0 2860 0 1 4625
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1677622389
transform 1 0 2876 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1677622389
transform 1 0 2852 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_60
timestamp 1677622389
transform 1 0 2860 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_123
timestamp 1677622389
transform 1 0 2868 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1677622389
transform 1 0 2868 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1677622389
transform 1 0 2900 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_124
timestamp 1677622389
transform 1 0 2892 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1677622389
transform 1 0 2924 0 1 4625
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1677622389
transform 1 0 2932 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1677622389
transform 1 0 2924 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_58
timestamp 1677622389
transform 1 0 2956 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_98
timestamp 1677622389
transform 1 0 2940 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1677622389
transform 1 0 3036 0 1 4645
box -3 -3 3 3
use M2_M1  M2_M1_125
timestamp 1677622389
transform 1 0 3044 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1677622389
transform 1 0 3060 0 1 4615
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1677622389
transform 1 0 3148 0 1 4665
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1677622389
transform 1 0 3148 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_59
timestamp 1677622389
transform 1 0 3084 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1677622389
transform 1 0 3140 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1677622389
transform 1 0 3060 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1677622389
transform 1 0 3060 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1677622389
transform 1 0 3084 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1677622389
transform 1 0 3188 0 1 4615
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1677622389
transform 1 0 3204 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_61
timestamp 1677622389
transform 1 0 3228 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1677622389
transform 1 0 3204 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1677622389
transform 1 0 3284 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1677622389
transform 1 0 3204 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1677622389
transform 1 0 3228 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_62
timestamp 1677622389
transform 1 0 3316 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1677622389
transform 1 0 3332 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1677622389
transform 1 0 3348 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_63
timestamp 1677622389
transform 1 0 3372 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1677622389
transform 1 0 3428 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1677622389
transform 1 0 3348 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1677622389
transform 1 0 3372 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1677622389
transform 1 0 3428 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1677622389
transform 1 0 3444 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1677622389
transform 1 0 3500 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1677622389
transform 1 0 3532 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1677622389
transform 1 0 3532 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_67
timestamp 1677622389
transform 1 0 3604 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1677622389
transform 1 0 3580 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_106
timestamp 1677622389
transform 1 0 3580 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1677622389
transform 1 0 3596 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1677622389
transform 1 0 3572 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1677622389
transform 1 0 3604 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_68
timestamp 1677622389
transform 1 0 3676 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1677622389
transform 1 0 3772 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1677622389
transform 1 0 3724 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1677622389
transform 1 0 3772 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1677622389
transform 1 0 3796 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1677622389
transform 1 0 3724 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_70
timestamp 1677622389
transform 1 0 3820 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1677622389
transform 1 0 3884 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1677622389
transform 1 0 3860 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_109
timestamp 1677622389
transform 1 0 3860 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1677622389
transform 1 0 3956 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_33
timestamp 1677622389
transform 1 0 4044 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_73
timestamp 1677622389
transform 1 0 4020 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1677622389
transform 1 0 3972 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1677622389
transform 1 0 4060 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1677622389
transform 1 0 4124 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1677622389
transform 1 0 4172 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1677622389
transform 1 0 4076 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1677622389
transform 1 0 4124 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1677622389
transform 1 0 4164 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1677622389
transform 1 0 4076 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1677622389
transform 1 0 4260 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1677622389
transform 1 0 4300 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1677622389
transform 1 0 4220 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_111
timestamp 1677622389
transform 1 0 4220 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_79
timestamp 1677622389
transform 1 0 4388 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1677622389
transform 1 0 4340 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_68
timestamp 1677622389
transform 1 0 4388 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1677622389
transform 1 0 4420 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1677622389
transform 1 0 4340 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_80
timestamp 1677622389
transform 1 0 4444 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1677622389
transform 1 0 4452 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1677622389
transform 1 0 4484 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1677622389
transform 1 0 4500 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_70
timestamp 1677622389
transform 1 0 4484 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1677622389
transform 1 0 4492 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1677622389
transform 1 0 4524 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_123
timestamp 1677622389
transform 1 0 4524 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_83
timestamp 1677622389
transform 1 0 4604 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1677622389
transform 1 0 4652 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1677622389
transform 1 0 4572 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1677622389
transform 1 0 4596 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1677622389
transform 1 0 4572 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1677622389
transform 1 0 4620 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1677622389
transform 1 0 4684 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_85
timestamp 1677622389
transform 1 0 4724 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1677622389
transform 1 0 4780 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1677622389
transform 1 0 4700 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1677622389
transform 1 0 4724 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1677622389
transform 1 0 4700 0 1 4595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_1
timestamp 1677622389
transform 1 0 4843 0 1 4670
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_2
timestamp 1677622389
transform 1 0 48 0 1 4570
box -10 -3 10 3
use FILL  FILL_0
timestamp 1677622389
transform 1 0 72 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1677622389
transform 1 0 80 0 1 4570
box -8 -3 104 105
use FILL  FILL_2
timestamp 1677622389
transform 1 0 176 0 1 4570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1677622389
transform 1 0 184 0 1 4570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1677622389
transform 1 0 192 0 1 4570
box -8 -3 16 105
use FILL  FILL_11
timestamp 1677622389
transform 1 0 200 0 1 4570
box -8 -3 16 105
use FILL  FILL_12
timestamp 1677622389
transform 1 0 208 0 1 4570
box -8 -3 16 105
use FILL  FILL_13
timestamp 1677622389
transform 1 0 216 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_125
timestamp 1677622389
transform 1 0 236 0 1 4575
box -3 -3 3 3
use FILL  FILL_14
timestamp 1677622389
transform 1 0 224 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1677622389
transform 1 0 232 0 1 4570
box -9 -3 26 105
use M3_M2  M3_M2_126
timestamp 1677622389
transform 1 0 268 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_1
timestamp 1677622389
transform 1 0 248 0 1 4570
box -8 -3 104 105
use FILL  FILL_15
timestamp 1677622389
transform 1 0 344 0 1 4570
box -8 -3 16 105
use FILL  FILL_16
timestamp 1677622389
transform 1 0 352 0 1 4570
box -8 -3 16 105
use FILL  FILL_17
timestamp 1677622389
transform 1 0 360 0 1 4570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1677622389
transform 1 0 368 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1677622389
transform 1 0 376 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1677622389
transform 1 0 392 0 1 4570
box -8 -3 104 105
use FILL  FILL_19
timestamp 1677622389
transform 1 0 488 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1677622389
transform 1 0 496 0 1 4570
box -8 -3 104 105
use FILL  FILL_20
timestamp 1677622389
transform 1 0 592 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1677622389
transform 1 0 600 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_4
timestamp 1677622389
transform 1 0 696 0 1 4570
box -9 -3 26 105
use FILL  FILL_21
timestamp 1677622389
transform 1 0 712 0 1 4570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1677622389
transform 1 0 720 0 1 4570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1677622389
transform 1 0 728 0 1 4570
box -8 -3 16 105
use FILL  FILL_24
timestamp 1677622389
transform 1 0 736 0 1 4570
box -8 -3 16 105
use FILL  FILL_25
timestamp 1677622389
transform 1 0 744 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1677622389
transform 1 0 752 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_5
timestamp 1677622389
transform 1 0 848 0 1 4570
box -9 -3 26 105
use FILL  FILL_26
timestamp 1677622389
transform 1 0 864 0 1 4570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1677622389
transform 1 0 872 0 1 4570
box -8 -3 16 105
use FILL  FILL_57
timestamp 1677622389
transform 1 0 880 0 1 4570
box -8 -3 16 105
use FILL  FILL_59
timestamp 1677622389
transform 1 0 888 0 1 4570
box -8 -3 16 105
use FILL  FILL_61
timestamp 1677622389
transform 1 0 896 0 1 4570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1677622389
transform 1 0 904 0 1 4570
box -8 -3 16 105
use FILL  FILL_65
timestamp 1677622389
transform 1 0 912 0 1 4570
box -8 -3 16 105
use FILL  FILL_67
timestamp 1677622389
transform 1 0 920 0 1 4570
box -8 -3 16 105
use FILL  FILL_69
timestamp 1677622389
transform 1 0 928 0 1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1677622389
transform 1 0 936 0 1 4570
box -8 -3 34 105
use FILL  FILL_70
timestamp 1677622389
transform 1 0 968 0 1 4570
box -8 -3 16 105
use FILL  FILL_71
timestamp 1677622389
transform 1 0 976 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1677622389
transform 1 0 984 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_8
timestamp 1677622389
transform -1 0 1096 0 1 4570
box -9 -3 26 105
use AOI22X1  AOI22X1_8
timestamp 1677622389
transform -1 0 1136 0 1 4570
box -8 -3 46 105
use FILL  FILL_72
timestamp 1677622389
transform 1 0 1136 0 1 4570
box -8 -3 16 105
use FILL  FILL_73
timestamp 1677622389
transform 1 0 1144 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1677622389
transform 1 0 1152 0 1 4570
box -9 -3 26 105
use FILL  FILL_78
timestamp 1677622389
transform 1 0 1168 0 1 4570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1677622389
transform 1 0 1176 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1677622389
transform -1 0 1280 0 1 4570
box -8 -3 104 105
use FILL  FILL_83
timestamp 1677622389
transform 1 0 1280 0 1 4570
box -8 -3 16 105
use FILL  FILL_84
timestamp 1677622389
transform 1 0 1288 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1677622389
transform 1 0 1296 0 1 4570
box -8 -3 104 105
use FILL  FILL_85
timestamp 1677622389
transform 1 0 1392 0 1 4570
box -8 -3 16 105
use FILL  FILL_86
timestamp 1677622389
transform 1 0 1400 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1677622389
transform 1 0 1408 0 1 4570
box -8 -3 104 105
use FILL  FILL_87
timestamp 1677622389
transform 1 0 1504 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_10
timestamp 1677622389
transform 1 0 1512 0 1 4570
box -9 -3 26 105
use FILL  FILL_88
timestamp 1677622389
transform 1 0 1528 0 1 4570
box -8 -3 16 105
use FILL  FILL_106
timestamp 1677622389
transform 1 0 1536 0 1 4570
box -8 -3 16 105
use FILL  FILL_108
timestamp 1677622389
transform 1 0 1544 0 1 4570
box -8 -3 16 105
use FILL  FILL_110
timestamp 1677622389
transform 1 0 1552 0 1 4570
box -8 -3 16 105
use FILL  FILL_112
timestamp 1677622389
transform 1 0 1560 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1677622389
transform 1 0 1568 0 1 4570
box -8 -3 104 105
use FILL  FILL_114
timestamp 1677622389
transform 1 0 1664 0 1 4570
box -8 -3 16 105
use FILL  FILL_115
timestamp 1677622389
transform 1 0 1672 0 1 4570
box -8 -3 16 105
use FILL  FILL_116
timestamp 1677622389
transform 1 0 1680 0 1 4570
box -8 -3 16 105
use FILL  FILL_125
timestamp 1677622389
transform 1 0 1688 0 1 4570
box -8 -3 16 105
use FILL  FILL_127
timestamp 1677622389
transform 1 0 1696 0 1 4570
box -8 -3 16 105
use FILL  FILL_129
timestamp 1677622389
transform 1 0 1704 0 1 4570
box -8 -3 16 105
use FILL  FILL_131
timestamp 1677622389
transform 1 0 1712 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_13
timestamp 1677622389
transform -1 0 1736 0 1 4570
box -9 -3 26 105
use FILL  FILL_132
timestamp 1677622389
transform 1 0 1736 0 1 4570
box -8 -3 16 105
use FILL  FILL_135
timestamp 1677622389
transform 1 0 1744 0 1 4570
box -8 -3 16 105
use FILL  FILL_137
timestamp 1677622389
transform 1 0 1752 0 1 4570
box -8 -3 16 105
use FILL  FILL_138
timestamp 1677622389
transform 1 0 1760 0 1 4570
box -8 -3 16 105
use FILL  FILL_139
timestamp 1677622389
transform 1 0 1768 0 1 4570
box -8 -3 16 105
use FILL  FILL_140
timestamp 1677622389
transform 1 0 1776 0 1 4570
box -8 -3 16 105
use FILL  FILL_141
timestamp 1677622389
transform 1 0 1784 0 1 4570
box -8 -3 16 105
use FILL  FILL_142
timestamp 1677622389
transform 1 0 1792 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_127
timestamp 1677622389
transform 1 0 1892 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_13
timestamp 1677622389
transform 1 0 1800 0 1 4570
box -8 -3 104 105
use M3_M2  M3_M2_128
timestamp 1677622389
transform 1 0 1908 0 1 4575
box -3 -3 3 3
use FILL  FILL_143
timestamp 1677622389
transform 1 0 1896 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1677622389
transform 1 0 1904 0 1 4570
box -9 -3 26 105
use FILL  FILL_144
timestamp 1677622389
transform 1 0 1920 0 1 4570
box -8 -3 16 105
use FILL  FILL_145
timestamp 1677622389
transform 1 0 1928 0 1 4570
box -8 -3 16 105
use FILL  FILL_150
timestamp 1677622389
transform 1 0 1936 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1677622389
transform 1 0 1944 0 1 4570
box -8 -3 104 105
use FILL  FILL_152
timestamp 1677622389
transform 1 0 2040 0 1 4570
box -8 -3 16 105
use FILL  FILL_153
timestamp 1677622389
transform 1 0 2048 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_17
timestamp 1677622389
transform -1 0 2072 0 1 4570
box -9 -3 26 105
use FILL  FILL_154
timestamp 1677622389
transform 1 0 2072 0 1 4570
box -8 -3 16 105
use FILL  FILL_155
timestamp 1677622389
transform 1 0 2080 0 1 4570
box -8 -3 16 105
use FILL  FILL_156
timestamp 1677622389
transform 1 0 2088 0 1 4570
box -8 -3 16 105
use FILL  FILL_166
timestamp 1677622389
transform 1 0 2096 0 1 4570
box -8 -3 16 105
use FILL  FILL_168
timestamp 1677622389
transform 1 0 2104 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_129
timestamp 1677622389
transform 1 0 2124 0 1 4575
box -3 -3 3 3
use FILL  FILL_170
timestamp 1677622389
transform 1 0 2112 0 1 4570
box -8 -3 16 105
use FILL  FILL_172
timestamp 1677622389
transform 1 0 2120 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1677622389
transform 1 0 2128 0 1 4570
box -8 -3 104 105
use FILL  FILL_174
timestamp 1677622389
transform 1 0 2224 0 1 4570
box -8 -3 16 105
use FILL  FILL_175
timestamp 1677622389
transform 1 0 2232 0 1 4570
box -8 -3 16 105
use FILL  FILL_176
timestamp 1677622389
transform 1 0 2240 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_18
timestamp 1677622389
transform 1 0 2248 0 1 4570
box -9 -3 26 105
use FILL  FILL_177
timestamp 1677622389
transform 1 0 2264 0 1 4570
box -8 -3 16 105
use FILL  FILL_186
timestamp 1677622389
transform 1 0 2272 0 1 4570
box -8 -3 16 105
use FILL  FILL_188
timestamp 1677622389
transform 1 0 2280 0 1 4570
box -8 -3 16 105
use FILL  FILL_189
timestamp 1677622389
transform 1 0 2288 0 1 4570
box -8 -3 16 105
use FILL  FILL_190
timestamp 1677622389
transform 1 0 2296 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_19
timestamp 1677622389
transform 1 0 2304 0 1 4570
box -9 -3 26 105
use FILL  FILL_191
timestamp 1677622389
transform 1 0 2320 0 1 4570
box -8 -3 16 105
use FILL  FILL_193
timestamp 1677622389
transform 1 0 2328 0 1 4570
box -8 -3 16 105
use FILL  FILL_195
timestamp 1677622389
transform 1 0 2336 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1677622389
transform -1 0 2440 0 1 4570
box -8 -3 104 105
use FILL  FILL_196
timestamp 1677622389
transform 1 0 2440 0 1 4570
box -8 -3 16 105
use FILL  FILL_197
timestamp 1677622389
transform 1 0 2448 0 1 4570
box -8 -3 16 105
use FILL  FILL_198
timestamp 1677622389
transform 1 0 2456 0 1 4570
box -8 -3 16 105
use FILL  FILL_199
timestamp 1677622389
transform 1 0 2464 0 1 4570
box -8 -3 16 105
use FILL  FILL_200
timestamp 1677622389
transform 1 0 2472 0 1 4570
box -8 -3 16 105
use FILL  FILL_201
timestamp 1677622389
transform 1 0 2480 0 1 4570
box -8 -3 16 105
use FILL  FILL_211
timestamp 1677622389
transform 1 0 2488 0 1 4570
box -8 -3 16 105
use FILL  FILL_213
timestamp 1677622389
transform 1 0 2496 0 1 4570
box -8 -3 16 105
use FILL  FILL_215
timestamp 1677622389
transform 1 0 2504 0 1 4570
box -8 -3 16 105
use FILL  FILL_217
timestamp 1677622389
transform 1 0 2512 0 1 4570
box -8 -3 16 105
use FILL  FILL_219
timestamp 1677622389
transform 1 0 2520 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1677622389
transform 1 0 2528 0 1 4570
box -9 -3 26 105
use FILL  FILL_220
timestamp 1677622389
transform 1 0 2544 0 1 4570
box -8 -3 16 105
use FILL  FILL_221
timestamp 1677622389
transform 1 0 2552 0 1 4570
box -8 -3 16 105
use FILL  FILL_222
timestamp 1677622389
transform 1 0 2560 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1677622389
transform 1 0 2568 0 1 4570
box -8 -3 104 105
use FILL  FILL_224
timestamp 1677622389
transform 1 0 2664 0 1 4570
box -8 -3 16 105
use FILL  FILL_238
timestamp 1677622389
transform 1 0 2672 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_21
timestamp 1677622389
transform 1 0 2680 0 1 4570
box -9 -3 26 105
use FILL  FILL_239
timestamp 1677622389
transform 1 0 2696 0 1 4570
box -8 -3 16 105
use FILL  FILL_240
timestamp 1677622389
transform 1 0 2704 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1677622389
transform 1 0 2712 0 1 4570
box -8 -3 104 105
use FILL  FILL_241
timestamp 1677622389
transform 1 0 2808 0 1 4570
box -8 -3 16 105
use FILL  FILL_252
timestamp 1677622389
transform 1 0 2816 0 1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1677622389
transform 1 0 2824 0 1 4570
box -8 -3 34 105
use FILL  FILL_254
timestamp 1677622389
transform 1 0 2856 0 1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_7
timestamp 1677622389
transform 1 0 2864 0 1 4570
box -8 -3 34 105
use FILL  FILL_257
timestamp 1677622389
transform 1 0 2896 0 1 4570
box -8 -3 16 105
use FILL  FILL_258
timestamp 1677622389
transform 1 0 2904 0 1 4570
box -8 -3 16 105
use FILL  FILL_259
timestamp 1677622389
transform 1 0 2912 0 1 4570
box -8 -3 16 105
use FILL  FILL_260
timestamp 1677622389
transform 1 0 2920 0 1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1677622389
transform -1 0 2960 0 1 4570
box -8 -3 34 105
use FILL  FILL_261
timestamp 1677622389
transform 1 0 2960 0 1 4570
box -8 -3 16 105
use FILL  FILL_262
timestamp 1677622389
transform 1 0 2968 0 1 4570
box -8 -3 16 105
use FILL  FILL_263
timestamp 1677622389
transform 1 0 2976 0 1 4570
box -8 -3 16 105
use FILL  FILL_264
timestamp 1677622389
transform 1 0 2984 0 1 4570
box -8 -3 16 105
use FILL  FILL_265
timestamp 1677622389
transform 1 0 2992 0 1 4570
box -8 -3 16 105
use FILL  FILL_266
timestamp 1677622389
transform 1 0 3000 0 1 4570
box -8 -3 16 105
use FILL  FILL_267
timestamp 1677622389
transform 1 0 3008 0 1 4570
box -8 -3 16 105
use FILL  FILL_275
timestamp 1677622389
transform 1 0 3016 0 1 4570
box -8 -3 16 105
use FILL  FILL_276
timestamp 1677622389
transform 1 0 3024 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_130
timestamp 1677622389
transform 1 0 3044 0 1 4575
box -3 -3 3 3
use FILL  FILL_277
timestamp 1677622389
transform 1 0 3032 0 1 4570
box -8 -3 16 105
use FILL  FILL_278
timestamp 1677622389
transform 1 0 3040 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1677622389
transform 1 0 3048 0 1 4570
box -8 -3 104 105
use FILL  FILL_279
timestamp 1677622389
transform 1 0 3144 0 1 4570
box -8 -3 16 105
use FILL  FILL_288
timestamp 1677622389
transform 1 0 3152 0 1 4570
box -8 -3 16 105
use FILL  FILL_290
timestamp 1677622389
transform 1 0 3160 0 1 4570
box -8 -3 16 105
use FILL  FILL_292
timestamp 1677622389
transform 1 0 3168 0 1 4570
box -8 -3 16 105
use FILL  FILL_294
timestamp 1677622389
transform 1 0 3176 0 1 4570
box -8 -3 16 105
use FILL  FILL_296
timestamp 1677622389
transform 1 0 3184 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_131
timestamp 1677622389
transform 1 0 3212 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_21
timestamp 1677622389
transform 1 0 3192 0 1 4570
box -8 -3 104 105
use FILL  FILL_297
timestamp 1677622389
transform 1 0 3288 0 1 4570
box -8 -3 16 105
use FILL  FILL_298
timestamp 1677622389
transform 1 0 3296 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_132
timestamp 1677622389
transform 1 0 3316 0 1 4575
box -3 -3 3 3
use INVX2  INVX2_24
timestamp 1677622389
transform 1 0 3304 0 1 4570
box -9 -3 26 105
use FILL  FILL_299
timestamp 1677622389
transform 1 0 3320 0 1 4570
box -8 -3 16 105
use FILL  FILL_300
timestamp 1677622389
transform 1 0 3328 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1677622389
transform 1 0 3336 0 1 4570
box -8 -3 104 105
use FILL  FILL_301
timestamp 1677622389
transform 1 0 3432 0 1 4570
box -8 -3 16 105
use FILL  FILL_314
timestamp 1677622389
transform 1 0 3440 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1677622389
transform -1 0 3544 0 1 4570
box -8 -3 104 105
use FILL  FILL_315
timestamp 1677622389
transform 1 0 3544 0 1 4570
box -8 -3 16 105
use FILL  FILL_323
timestamp 1677622389
transform 1 0 3552 0 1 4570
box -8 -3 16 105
use FILL  FILL_324
timestamp 1677622389
transform 1 0 3560 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_133
timestamp 1677622389
transform 1 0 3604 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_24
timestamp 1677622389
transform 1 0 3568 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_27
timestamp 1677622389
transform 1 0 3664 0 1 4570
box -9 -3 26 105
use FILL  FILL_325
timestamp 1677622389
transform 1 0 3680 0 1 4570
box -8 -3 16 105
use FILL  FILL_333
timestamp 1677622389
transform 1 0 3688 0 1 4570
box -8 -3 16 105
use FILL  FILL_334
timestamp 1677622389
transform 1 0 3696 0 1 4570
box -8 -3 16 105
use FILL  FILL_335
timestamp 1677622389
transform 1 0 3704 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1677622389
transform 1 0 3712 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_28
timestamp 1677622389
transform 1 0 3808 0 1 4570
box -9 -3 26 105
use FILL  FILL_336
timestamp 1677622389
transform 1 0 3824 0 1 4570
box -8 -3 16 105
use FILL  FILL_345
timestamp 1677622389
transform 1 0 3832 0 1 4570
box -8 -3 16 105
use FILL  FILL_347
timestamp 1677622389
transform 1 0 3840 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1677622389
transform 1 0 3848 0 1 4570
box -8 -3 104 105
use FILL  FILL_348
timestamp 1677622389
transform 1 0 3944 0 1 4570
box -8 -3 16 105
use FILL  FILL_353
timestamp 1677622389
transform 1 0 3952 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_134
timestamp 1677622389
transform 1 0 3972 0 1 4575
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1677622389
transform 1 0 4052 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_27
timestamp 1677622389
transform 1 0 3960 0 1 4570
box -8 -3 104 105
use FILL  FILL_354
timestamp 1677622389
transform 1 0 4056 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1677622389
transform 1 0 4064 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_29
timestamp 1677622389
transform 1 0 4160 0 1 4570
box -9 -3 26 105
use FILL  FILL_355
timestamp 1677622389
transform 1 0 4176 0 1 4570
box -8 -3 16 105
use FILL  FILL_356
timestamp 1677622389
transform 1 0 4184 0 1 4570
box -8 -3 16 105
use FILL  FILL_371
timestamp 1677622389
transform 1 0 4192 0 1 4570
box -8 -3 16 105
use FILL  FILL_373
timestamp 1677622389
transform 1 0 4200 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1677622389
transform 1 0 4208 0 1 4570
box -8 -3 104 105
use FILL  FILL_375
timestamp 1677622389
transform 1 0 4304 0 1 4570
box -8 -3 16 105
use FILL  FILL_382
timestamp 1677622389
transform 1 0 4312 0 1 4570
box -8 -3 16 105
use FILL  FILL_384
timestamp 1677622389
transform 1 0 4320 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1677622389
transform 1 0 4328 0 1 4570
box -8 -3 104 105
use FILL  FILL_385
timestamp 1677622389
transform 1 0 4424 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_34
timestamp 1677622389
transform 1 0 4432 0 1 4570
box -9 -3 26 105
use FILL  FILL_386
timestamp 1677622389
transform 1 0 4448 0 1 4570
box -8 -3 16 105
use FILL  FILL_394
timestamp 1677622389
transform 1 0 4456 0 1 4570
box -8 -3 16 105
use FILL  FILL_396
timestamp 1677622389
transform 1 0 4464 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_136
timestamp 1677622389
transform 1 0 4500 0 1 4575
box -3 -3 3 3
use OAI22X1  OAI22X1_18
timestamp 1677622389
transform 1 0 4472 0 1 4570
box -8 -3 46 105
use FILL  FILL_398
timestamp 1677622389
transform 1 0 4512 0 1 4570
box -8 -3 16 105
use FILL  FILL_399
timestamp 1677622389
transform 1 0 4520 0 1 4570
box -8 -3 16 105
use FILL  FILL_400
timestamp 1677622389
transform 1 0 4528 0 1 4570
box -8 -3 16 105
use FILL  FILL_401
timestamp 1677622389
transform 1 0 4536 0 1 4570
box -8 -3 16 105
use FILL  FILL_402
timestamp 1677622389
transform 1 0 4544 0 1 4570
box -8 -3 16 105
use FILL  FILL_403
timestamp 1677622389
transform 1 0 4552 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_137
timestamp 1677622389
transform 1 0 4580 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_31
timestamp 1677622389
transform 1 0 4560 0 1 4570
box -8 -3 104 105
use FILL  FILL_404
timestamp 1677622389
transform 1 0 4656 0 1 4570
box -8 -3 16 105
use FILL  FILL_405
timestamp 1677622389
transform 1 0 4664 0 1 4570
box -8 -3 16 105
use FILL  FILL_406
timestamp 1677622389
transform 1 0 4672 0 1 4570
box -8 -3 16 105
use FILL  FILL_407
timestamp 1677622389
transform 1 0 4680 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1677622389
transform 1 0 4688 0 1 4570
box -8 -3 104 105
use FILL  FILL_408
timestamp 1677622389
transform 1 0 4784 0 1 4570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_3
timestamp 1677622389
transform 1 0 4819 0 1 4570
box -10 -3 10 3
use M2_M1  M2_M1_145
timestamp 1677622389
transform 1 0 92 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1677622389
transform 1 0 92 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1677622389
transform 1 0 108 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1677622389
transform 1 0 116 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_283
timestamp 1677622389
transform 1 0 100 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1677622389
transform 1 0 116 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_175
timestamp 1677622389
transform 1 0 140 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1677622389
transform 1 0 140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1677622389
transform 1 0 132 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1677622389
transform 1 0 148 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_260
timestamp 1677622389
transform 1 0 148 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1677622389
transform 1 0 132 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1677622389
transform 1 0 172 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1677622389
transform 1 0 196 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_148
timestamp 1677622389
transform 1 0 196 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1677622389
transform 1 0 236 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1677622389
transform 1 0 212 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_218
timestamp 1677622389
transform 1 0 220 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1677622389
transform 1 0 228 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1677622389
transform 1 0 236 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1677622389
transform 1 0 204 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1677622389
transform 1 0 212 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_288
timestamp 1677622389
transform 1 0 220 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_346
timestamp 1677622389
transform 1 0 204 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_289
timestamp 1677622389
transform 1 0 244 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1677622389
transform 1 0 252 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1677622389
transform 1 0 260 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_291
timestamp 1677622389
transform 1 0 268 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1677622389
transform 1 0 284 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1677622389
transform 1 0 252 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1677622389
transform 1 0 284 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1677622389
transform 1 0 308 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1677622389
transform 1 0 308 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1677622389
transform 1 0 308 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1677622389
transform 1 0 324 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1677622389
transform 1 0 324 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1677622389
transform 1 0 340 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1677622389
transform 1 0 380 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1677622389
transform 1 0 372 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1677622389
transform 1 0 348 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1677622389
transform 1 0 356 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1677622389
transform 1 0 372 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1677622389
transform 1 0 364 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1677622389
transform 1 0 380 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1677622389
transform 1 0 388 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1677622389
transform 1 0 404 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1677622389
transform 1 0 420 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_302
timestamp 1677622389
transform 1 0 420 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1677622389
transform 1 0 436 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1677622389
transform 1 0 484 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1677622389
transform 1 0 484 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1677622389
transform 1 0 492 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1677622389
transform 1 0 492 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1677622389
transform 1 0 532 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1677622389
transform 1 0 516 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1677622389
transform 1 0 524 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1677622389
transform 1 0 540 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1677622389
transform 1 0 516 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1677622389
transform 1 0 540 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1677622389
transform 1 0 532 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1677622389
transform 1 0 540 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1677622389
transform 1 0 572 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1677622389
transform 1 0 564 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1677622389
transform 1 0 588 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1677622389
transform 1 0 604 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1677622389
transform 1 0 564 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1677622389
transform 1 0 572 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1677622389
transform 1 0 588 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1677622389
transform 1 0 604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1677622389
transform 1 0 564 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1677622389
transform 1 0 580 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1677622389
transform 1 0 588 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_305
timestamp 1677622389
transform 1 0 596 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1677622389
transform 1 0 564 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1677622389
transform 1 0 596 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1677622389
transform 1 0 612 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_306
timestamp 1677622389
transform 1 0 620 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_264
timestamp 1677622389
transform 1 0 620 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1677622389
transform 1 0 644 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1677622389
transform 1 0 716 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_163
timestamp 1677622389
transform 1 0 692 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1677622389
transform 1 0 708 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_184
timestamp 1677622389
transform 1 0 732 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1677622389
transform 1 0 764 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1677622389
transform 1 0 812 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1677622389
transform 1 0 732 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1677622389
transform 1 0 820 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1677622389
transform 1 0 700 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1677622389
transform 1 0 716 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1677622389
transform 1 0 756 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1677622389
transform 1 0 812 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1677622389
transform 1 0 708 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1677622389
transform 1 0 764 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1677622389
transform 1 0 772 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_142
timestamp 1677622389
transform 1 0 868 0 1 4545
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1677622389
transform 1 0 860 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1677622389
transform 1 0 828 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1677622389
transform 1 0 844 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1677622389
transform 1 0 860 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_307
timestamp 1677622389
transform 1 0 820 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1677622389
transform 1 0 836 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1677622389
transform 1 0 868 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1677622389
transform 1 0 900 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1677622389
transform 1 0 956 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1677622389
transform 1 0 956 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1677622389
transform 1 0 980 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_314
timestamp 1677622389
transform 1 0 948 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1677622389
transform 1 0 964 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_267
timestamp 1677622389
transform 1 0 964 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1677622389
transform 1 0 988 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1677622389
transform 1 0 1004 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_424
timestamp 1677622389
transform 1 0 1004 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_308
timestamp 1677622389
transform 1 0 996 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1677622389
transform 1 0 1108 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1677622389
transform 1 0 1020 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1677622389
transform 1 0 1108 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1677622389
transform 1 0 1052 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1677622389
transform 1 0 1100 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1677622389
transform 1 0 1108 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1677622389
transform 1 0 1124 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1677622389
transform 1 0 1140 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1677622389
transform 1 0 1148 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_309
timestamp 1677622389
transform 1 0 1020 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1677622389
transform 1 0 1092 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1677622389
transform 1 0 1108 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1677622389
transform 1 0 1156 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1677622389
transform 1 0 1148 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1677622389
transform 1 0 1164 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_173
timestamp 1677622389
transform 1 0 1164 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1677622389
transform 1 0 1172 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1677622389
transform 1 0 1188 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1677622389
transform 1 0 1204 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1677622389
transform 1 0 1212 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1677622389
transform 1 0 1212 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1677622389
transform 1 0 1228 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1677622389
transform 1 0 1228 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_142
timestamp 1677622389
transform 1 0 1276 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1677622389
transform 1 0 1268 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1677622389
transform 1 0 1268 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1677622389
transform 1 0 1252 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1677622389
transform 1 0 1236 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_269
timestamp 1677622389
transform 1 0 1252 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_427
timestamp 1677622389
transform 1 0 1268 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1677622389
transform 1 0 1236 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1677622389
transform 1 0 1276 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_311
timestamp 1677622389
transform 1 0 1268 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1677622389
transform 1 0 1308 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1677622389
transform 1 0 1308 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1677622389
transform 1 0 1292 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_270
timestamp 1677622389
transform 1 0 1292 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_428
timestamp 1677622389
transform 1 0 1308 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1677622389
transform 1 0 1316 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1677622389
transform 1 0 1316 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1677622389
transform 1 0 1332 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1677622389
transform 1 0 1308 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1677622389
transform 1 0 1332 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1677622389
transform 1 0 1348 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_325
timestamp 1677622389
transform 1 0 1348 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1677622389
transform 1 0 1356 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1677622389
transform 1 0 1356 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1677622389
transform 1 0 1396 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_182
timestamp 1677622389
transform 1 0 1380 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1677622389
transform 1 0 1388 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1677622389
transform 1 0 1404 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1677622389
transform 1 0 1388 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_326
timestamp 1677622389
transform 1 0 1396 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1677622389
transform 1 0 1428 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1677622389
transform 1 0 1436 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1677622389
transform 1 0 1436 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1677622389
transform 1 0 1428 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_327
timestamp 1677622389
transform 1 0 1460 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1677622389
transform 1 0 1476 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1677622389
transform 1 0 1476 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1677622389
transform 1 0 1500 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1677622389
transform 1 0 1524 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1677622389
transform 1 0 1508 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1677622389
transform 1 0 1500 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1677622389
transform 1 0 1516 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1677622389
transform 1 0 1516 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1677622389
transform 1 0 1508 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1677622389
transform 1 0 1588 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1677622389
transform 1 0 1588 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1677622389
transform 1 0 1596 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1677622389
transform 1 0 1612 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1677622389
transform 1 0 1596 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_330
timestamp 1677622389
transform 1 0 1604 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1677622389
transform 1 0 1620 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1677622389
transform 1 0 1628 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_273
timestamp 1677622389
transform 1 0 1604 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1677622389
transform 1 0 1628 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1677622389
transform 1 0 1620 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_192
timestamp 1677622389
transform 1 0 1652 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1677622389
transform 1 0 1660 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1677622389
transform 1 0 1684 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_333
timestamp 1677622389
transform 1 0 1684 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_348
timestamp 1677622389
transform 1 0 1684 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_194
timestamp 1677622389
transform 1 0 1692 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_157
timestamp 1677622389
transform 1 0 1732 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_195
timestamp 1677622389
transform 1 0 1724 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_220
timestamp 1677622389
transform 1 0 1732 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1677622389
transform 1 0 1764 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1677622389
transform 1 0 1812 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1677622389
transform 1 0 1764 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1677622389
transform 1 0 1812 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_275
timestamp 1677622389
transform 1 0 1812 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_197
timestamp 1677622389
transform 1 0 1852 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1677622389
transform 1 0 1852 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1677622389
transform 1 0 1876 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1677622389
transform 1 0 1868 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_198
timestamp 1677622389
transform 1 0 1908 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1677622389
transform 1 0 1868 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1677622389
transform 1 0 1876 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1677622389
transform 1 0 1892 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1677622389
transform 1 0 1908 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1677622389
transform 1 0 1916 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_276
timestamp 1677622389
transform 1 0 1916 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1677622389
transform 1 0 1908 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1677622389
transform 1 0 1932 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_340
timestamp 1677622389
transform 1 0 1932 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_198
timestamp 1677622389
transform 1 0 1996 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_199
timestamp 1677622389
transform 1 0 1972 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1677622389
transform 1 0 1980 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1677622389
transform 1 0 1996 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1677622389
transform 1 0 1972 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1677622389
transform 1 0 1980 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_342
timestamp 1677622389
transform 1 0 1988 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1677622389
transform 1 0 2004 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1677622389
transform 1 0 1972 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1677622389
transform 1 0 2004 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1677622389
transform 1 0 2036 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1677622389
transform 1 0 2036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1677622389
transform 1 0 2076 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1677622389
transform 1 0 2068 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1677622389
transform 1 0 2076 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_345
timestamp 1677622389
transform 1 0 2084 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_315
timestamp 1677622389
transform 1 0 2108 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1677622389
transform 1 0 2124 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_199
timestamp 1677622389
transform 1 0 2148 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1677622389
transform 1 0 2148 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1677622389
transform 1 0 2140 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1677622389
transform 1 0 2156 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1677622389
transform 1 0 2140 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1677622389
transform 1 0 2156 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_348
timestamp 1677622389
transform 1 0 2180 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1677622389
transform 1 0 2244 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_206
timestamp 1677622389
transform 1 0 2220 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1677622389
transform 1 0 2228 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1677622389
transform 1 0 2244 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_278
timestamp 1677622389
transform 1 0 2236 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1677622389
transform 1 0 2244 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_351
timestamp 1677622389
transform 1 0 2276 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1677622389
transform 1 0 2292 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_144
timestamp 1677622389
transform 1 0 2332 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1677622389
transform 1 0 2324 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1677622389
transform 1 0 2324 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1677622389
transform 1 0 2300 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1677622389
transform 1 0 2316 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1677622389
transform 1 0 2324 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_350
timestamp 1677622389
transform 1 0 2284 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_209
timestamp 1677622389
transform 1 0 2332 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_279
timestamp 1677622389
transform 1 0 2324 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1677622389
transform 1 0 2388 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_210
timestamp 1677622389
transform 1 0 2372 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1677622389
transform 1 0 2380 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1677622389
transform 1 0 2388 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1677622389
transform 1 0 2396 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1677622389
transform 1 0 2380 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1677622389
transform 1 0 2380 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_356
timestamp 1677622389
transform 1 0 2396 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_280
timestamp 1677622389
transform 1 0 2396 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_213
timestamp 1677622389
transform 1 0 2460 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1677622389
transform 1 0 2476 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1677622389
transform 1 0 2468 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1677622389
transform 1 0 2468 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_358
timestamp 1677622389
transform 1 0 2484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_317
timestamp 1677622389
transform 1 0 2484 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_215
timestamp 1677622389
transform 1 0 2524 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1677622389
transform 1 0 2540 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1677622389
transform 1 0 2556 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1677622389
transform 1 0 2572 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1677622389
transform 1 0 2660 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1677622389
transform 1 0 2684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1677622389
transform 1 0 2692 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1677622389
transform 1 0 2716 0 1 4545
box -2 -2 2 2
use M3_M2  M3_M2_223
timestamp 1677622389
transform 1 0 2716 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_363
timestamp 1677622389
transform 1 0 2740 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_162
timestamp 1677622389
transform 1 0 2780 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1677622389
transform 1 0 2780 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_163
timestamp 1677622389
transform 1 0 2804 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1677622389
transform 1 0 2796 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1677622389
transform 1 0 2804 0 1 4545
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1677622389
transform 1 0 2828 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1677622389
transform 1 0 2836 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1677622389
transform 1 0 2844 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1677622389
transform 1 0 2836 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1677622389
transform 1 0 2860 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1677622389
transform 1 0 2852 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_351
timestamp 1677622389
transform 1 0 2844 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_366
timestamp 1677622389
transform 1 0 2876 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1677622389
transform 1 0 2892 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_222
timestamp 1677622389
transform 1 0 2924 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1677622389
transform 1 0 2932 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1677622389
transform 1 0 2908 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1677622389
transform 1 0 2932 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1677622389
transform 1 0 2964 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_224
timestamp 1677622389
transform 1 0 2964 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1677622389
transform 1 0 2972 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1677622389
transform 1 0 2956 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1677622389
transform 1 0 2932 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1677622389
transform 1 0 2940 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_318
timestamp 1677622389
transform 1 0 2940 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1677622389
transform 1 0 2972 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_369
timestamp 1677622389
transform 1 0 2980 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1677622389
transform 1 0 2996 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1677622389
transform 1 0 2972 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1677622389
transform 1 0 2980 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_319
timestamp 1677622389
transform 1 0 2980 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1677622389
transform 1 0 3068 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1677622389
transform 1 0 3044 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1677622389
transform 1 0 3020 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_226
timestamp 1677622389
transform 1 0 3028 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_227
timestamp 1677622389
transform 1 0 3036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1677622389
transform 1 0 3044 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1677622389
transform 1 0 3060 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1677622389
transform 1 0 3028 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1677622389
transform 1 0 3044 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1677622389
transform 1 0 3068 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1677622389
transform 1 0 3068 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1677622389
transform 1 0 3044 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1677622389
transform 1 0 3092 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1677622389
transform 1 0 3084 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_321
timestamp 1677622389
transform 1 0 3092 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_231
timestamp 1677622389
transform 1 0 3140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1677622389
transform 1 0 3148 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1677622389
transform 1 0 3148 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1677622389
transform 1 0 3148 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1677622389
transform 1 0 3204 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1677622389
transform 1 0 3220 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1677622389
transform 1 0 3212 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1677622389
transform 1 0 3220 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1677622389
transform 1 0 3252 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1677622389
transform 1 0 3276 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_235
timestamp 1677622389
transform 1 0 3284 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1677622389
transform 1 0 3276 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1677622389
transform 1 0 3292 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_343
timestamp 1677622389
transform 1 0 3292 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1677622389
transform 1 0 3308 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_236
timestamp 1677622389
transform 1 0 3308 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1677622389
transform 1 0 3316 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_379
timestamp 1677622389
transform 1 0 3316 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1677622389
transform 1 0 3332 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1677622389
transform 1 0 3356 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1677622389
transform 1 0 3340 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1677622389
transform 1 0 3348 0 1 4505
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1677622389
transform 1 0 3396 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1677622389
transform 1 0 3396 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1677622389
transform 1 0 3372 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1677622389
transform 1 0 3380 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1677622389
transform 1 0 3372 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_438
timestamp 1677622389
transform 1 0 3396 0 1 4505
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1677622389
transform 1 0 3396 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1677622389
transform 1 0 3444 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1677622389
transform 1 0 3436 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_436
timestamp 1677622389
transform 1 0 3436 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1677622389
transform 1 0 3460 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1677622389
transform 1 0 3460 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_239
timestamp 1677622389
transform 1 0 3460 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1677622389
transform 1 0 3500 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1677622389
transform 1 0 3484 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1677622389
transform 1 0 3492 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1677622389
transform 1 0 3508 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1677622389
transform 1 0 3484 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1677622389
transform 1 0 3508 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_385
timestamp 1677622389
transform 1 0 3524 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_166
timestamp 1677622389
transform 1 0 3540 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1677622389
transform 1 0 3548 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_241
timestamp 1677622389
transform 1 0 3540 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1677622389
transform 1 0 3548 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1677622389
transform 1 0 3548 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1677622389
transform 1 0 3588 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1677622389
transform 1 0 3580 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_243
timestamp 1677622389
transform 1 0 3572 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1677622389
transform 1 0 3588 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1677622389
transform 1 0 3564 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1677622389
transform 1 0 3580 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1677622389
transform 1 0 3620 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_168
timestamp 1677622389
transform 1 0 3652 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1677622389
transform 1 0 3660 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_246
timestamp 1677622389
transform 1 0 3652 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1677622389
transform 1 0 3660 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1677622389
transform 1 0 3628 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1677622389
transform 1 0 3644 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_283
timestamp 1677622389
transform 1 0 3620 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1677622389
transform 1 0 3644 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1677622389
transform 1 0 3628 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_248
timestamp 1677622389
transform 1 0 3676 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_354
timestamp 1677622389
transform 1 0 3668 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_390
timestamp 1677622389
transform 1 0 3692 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1677622389
transform 1 0 3700 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_284
timestamp 1677622389
transform 1 0 3692 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1677622389
transform 1 0 3708 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_392
timestamp 1677622389
transform 1 0 3716 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1677622389
transform 1 0 3732 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_345
timestamp 1677622389
transform 1 0 3700 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1677622389
transform 1 0 3732 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1677622389
transform 1 0 3780 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1677622389
transform 1 0 3804 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_249
timestamp 1677622389
transform 1 0 3772 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1677622389
transform 1 0 3780 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1677622389
transform 1 0 3796 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1677622389
transform 1 0 3756 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1677622389
transform 1 0 3764 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1677622389
transform 1 0 3772 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_395
timestamp 1677622389
transform 1 0 3788 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1677622389
transform 1 0 3804 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_325
timestamp 1677622389
transform 1 0 3788 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1677622389
transform 1 0 3820 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_252
timestamp 1677622389
transform 1 0 3820 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1677622389
transform 1 0 3900 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1677622389
transform 1 0 3868 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1677622389
transform 1 0 3884 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1677622389
transform 1 0 3900 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1677622389
transform 1 0 3860 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1677622389
transform 1 0 3876 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1677622389
transform 1 0 3892 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1677622389
transform 1 0 3860 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1677622389
transform 1 0 3876 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1677622389
transform 1 0 3900 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_400
timestamp 1677622389
transform 1 0 3908 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1677622389
transform 1 0 3924 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1677622389
transform 1 0 3932 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1677622389
transform 1 0 3884 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1677622389
transform 1 0 3932 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_256
timestamp 1677622389
transform 1 0 3948 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_289
timestamp 1677622389
transform 1 0 3948 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1677622389
transform 1 0 3972 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1677622389
transform 1 0 4044 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_258
timestamp 1677622389
transform 1 0 4012 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1677622389
transform 1 0 4028 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1677622389
transform 1 0 4044 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1677622389
transform 1 0 4020 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1677622389
transform 1 0 4036 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1677622389
transform 1 0 4044 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1677622389
transform 1 0 4020 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1677622389
transform 1 0 4044 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1677622389
transform 1 0 4060 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_292
timestamp 1677622389
transform 1 0 4076 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_406
timestamp 1677622389
transform 1 0 4084 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_172
timestamp 1677622389
transform 1 0 4148 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1677622389
transform 1 0 4172 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_262
timestamp 1677622389
transform 1 0 4140 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1677622389
transform 1 0 4148 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1677622389
transform 1 0 4164 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1677622389
transform 1 0 4156 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1677622389
transform 1 0 4172 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1677622389
transform 1 0 4172 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1677622389
transform 1 0 4196 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1677622389
transform 1 0 4204 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1677622389
transform 1 0 4204 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1677622389
transform 1 0 4244 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1677622389
transform 1 0 4276 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_267
timestamp 1677622389
transform 1 0 4244 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1677622389
transform 1 0 4260 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1677622389
transform 1 0 4276 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1677622389
transform 1 0 4252 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1677622389
transform 1 0 4260 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_410
timestamp 1677622389
transform 1 0 4268 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1677622389
transform 1 0 4284 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1677622389
transform 1 0 4300 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_256
timestamp 1677622389
transform 1 0 4324 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1677622389
transform 1 0 4364 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1677622389
transform 1 0 4348 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_412
timestamp 1677622389
transform 1 0 4332 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1677622389
transform 1 0 4348 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_327
timestamp 1677622389
transform 1 0 4332 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_271
timestamp 1677622389
transform 1 0 4380 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1677622389
transform 1 0 4380 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1677622389
transform 1 0 4396 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1677622389
transform 1 0 4396 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1677622389
transform 1 0 4396 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1677622389
transform 1 0 4436 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_273
timestamp 1677622389
transform 1 0 4420 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1677622389
transform 1 0 4436 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1677622389
transform 1 0 4412 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_257
timestamp 1677622389
transform 1 0 4420 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_416
timestamp 1677622389
transform 1 0 4428 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1677622389
transform 1 0 4412 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1677622389
transform 1 0 4452 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1677622389
transform 1 0 4460 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1677622389
transform 1 0 4588 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1677622389
transform 1 0 4484 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1677622389
transform 1 0 4572 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1677622389
transform 1 0 4484 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1677622389
transform 1 0 4508 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1677622389
transform 1 0 4620 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_276
timestamp 1677622389
transform 1 0 4588 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1677622389
transform 1 0 4596 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1677622389
transform 1 0 4604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1677622389
transform 1 0 4620 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1677622389
transform 1 0 4580 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1677622389
transform 1 0 4596 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1677622389
transform 1 0 4612 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_295
timestamp 1677622389
transform 1 0 4612 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_421
timestamp 1677622389
transform 1 0 4628 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_296
timestamp 1677622389
transform 1 0 4628 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1677622389
transform 1 0 4644 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1677622389
transform 1 0 4700 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_279
timestamp 1677622389
transform 1 0 4652 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1677622389
transform 1 0 4668 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1677622389
transform 1 0 4676 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_281
timestamp 1677622389
transform 1 0 4684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1677622389
transform 1 0 4700 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1677622389
transform 1 0 4676 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1677622389
transform 1 0 4692 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_297
timestamp 1677622389
transform 1 0 4692 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1677622389
transform 1 0 4788 0 1 4515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_4
timestamp 1677622389
transform 1 0 24 0 1 4470
box -10 -3 10 3
use FILL  FILL_1
timestamp 1677622389
transform 1 0 72 0 -1 4570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1677622389
transform 1 0 80 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1677622389
transform 1 0 88 0 -1 4570
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1677622389
transform 1 0 104 0 -1 4570
box -9 -3 26 105
use FILL  FILL_4
timestamp 1677622389
transform 1 0 120 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1677622389
transform -1 0 168 0 -1 4570
box -8 -3 46 105
use FILL  FILL_5
timestamp 1677622389
transform 1 0 168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1677622389
transform 1 0 176 0 -1 4570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1677622389
transform 1 0 184 0 -1 4570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1677622389
transform 1 0 192 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1677622389
transform 1 0 200 0 -1 4570
box -8 -3 46 105
use FILL  FILL_27
timestamp 1677622389
transform 1 0 240 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1677622389
transform 1 0 248 0 -1 4570
box -8 -3 46 105
use FILL  FILL_28
timestamp 1677622389
transform 1 0 288 0 -1 4570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1677622389
transform 1 0 296 0 -1 4570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1677622389
transform 1 0 304 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1677622389
transform -1 0 328 0 -1 4570
box -9 -3 26 105
use FILL  FILL_31
timestamp 1677622389
transform 1 0 328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1677622389
transform 1 0 336 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_357
timestamp 1677622389
transform 1 0 388 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_3
timestamp 1677622389
transform -1 0 384 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1677622389
transform 1 0 384 0 -1 4570
box -8 -3 46 105
use FILL  FILL_33
timestamp 1677622389
transform 1 0 424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1677622389
transform 1 0 432 0 -1 4570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1677622389
transform 1 0 440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1677622389
transform 1 0 448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1677622389
transform 1 0 456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_38
timestamp 1677622389
transform 1 0 464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_39
timestamp 1677622389
transform 1 0 472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1677622389
transform 1 0 480 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1677622389
transform 1 0 488 0 -1 4570
box -9 -3 26 105
use FILL  FILL_41
timestamp 1677622389
transform 1 0 504 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_358
timestamp 1677622389
transform 1 0 524 0 1 4475
box -3 -3 3 3
use FILL  FILL_42
timestamp 1677622389
transform 1 0 512 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1677622389
transform 1 0 520 0 -1 4570
box -8 -3 46 105
use FILL  FILL_43
timestamp 1677622389
transform 1 0 560 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_0
timestamp 1677622389
transform 1 0 568 0 -1 4570
box -8 -3 46 105
use FILL  FILL_44
timestamp 1677622389
transform 1 0 608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_45
timestamp 1677622389
transform 1 0 616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_46
timestamp 1677622389
transform 1 0 624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_47
timestamp 1677622389
transform 1 0 632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1677622389
transform 1 0 640 0 -1 4570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1677622389
transform 1 0 648 0 -1 4570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1677622389
transform 1 0 656 0 -1 4570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1677622389
transform 1 0 664 0 -1 4570
box -8 -3 16 105
use FILL  FILL_52
timestamp 1677622389
transform 1 0 672 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1677622389
transform -1 0 720 0 -1 4570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1677622389
transform 1 0 720 0 -1 4570
box -8 -3 104 105
use M3_M2  M3_M2_359
timestamp 1677622389
transform 1 0 828 0 1 4475
box -3 -3 3 3
use FILL  FILL_53
timestamp 1677622389
transform 1 0 816 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_7
timestamp 1677622389
transform 1 0 824 0 -1 4570
box -8 -3 46 105
use FILL  FILL_54
timestamp 1677622389
transform 1 0 864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1677622389
transform 1 0 872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1677622389
transform 1 0 880 0 -1 4570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1677622389
transform 1 0 888 0 -1 4570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1677622389
transform 1 0 896 0 -1 4570
box -8 -3 16 105
use FILL  FILL_64
timestamp 1677622389
transform 1 0 904 0 -1 4570
box -8 -3 16 105
use FILL  FILL_66
timestamp 1677622389
transform 1 0 912 0 -1 4570
box -8 -3 16 105
use FILL  FILL_68
timestamp 1677622389
transform 1 0 920 0 -1 4570
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1677622389
transform 1 0 928 0 -1 4570
box -8 -3 32 105
use OAI21X1  OAI21X1_1
timestamp 1677622389
transform 1 0 952 0 -1 4570
box -8 -3 34 105
use FILL  FILL_74
timestamp 1677622389
transform 1 0 984 0 -1 4570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1677622389
transform 1 0 992 0 -1 4570
box -8 -3 16 105
use FILL  FILL_76
timestamp 1677622389
transform 1 0 1000 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1677622389
transform 1 0 1008 0 -1 4570
box -8 -3 104 105
use AOI22X1  AOI22X1_9
timestamp 1677622389
transform 1 0 1104 0 -1 4570
box -8 -3 46 105
use FILL  FILL_77
timestamp 1677622389
transform 1 0 1144 0 -1 4570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1677622389
transform 1 0 1152 0 -1 4570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1677622389
transform 1 0 1160 0 -1 4570
box -8 -3 16 105
use FILL  FILL_81
timestamp 1677622389
transform 1 0 1168 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1677622389
transform 1 0 1176 0 -1 4570
box -8 -3 34 105
use FILL  FILL_89
timestamp 1677622389
transform 1 0 1208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_90
timestamp 1677622389
transform 1 0 1216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_91
timestamp 1677622389
transform 1 0 1224 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1677622389
transform -1 0 1264 0 -1 4570
box -8 -3 34 105
use FILL  FILL_92
timestamp 1677622389
transform 1 0 1264 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1677622389
transform -1 0 1304 0 -1 4570
box -8 -3 34 105
use FILL  FILL_93
timestamp 1677622389
transform 1 0 1304 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1677622389
transform -1 0 1344 0 -1 4570
box -8 -3 34 105
use FILL  FILL_94
timestamp 1677622389
transform 1 0 1344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_95
timestamp 1677622389
transform 1 0 1352 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1677622389
transform -1 0 1376 0 -1 4570
box -9 -3 26 105
use FILL  FILL_96
timestamp 1677622389
transform 1 0 1376 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_1
timestamp 1677622389
transform -1 0 1424 0 -1 4570
box -8 -3 46 105
use FILL  FILL_97
timestamp 1677622389
transform 1 0 1424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_98
timestamp 1677622389
transform 1 0 1432 0 -1 4570
box -8 -3 16 105
use FILL  FILL_99
timestamp 1677622389
transform 1 0 1440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_100
timestamp 1677622389
transform 1 0 1448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_101
timestamp 1677622389
transform 1 0 1456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_102
timestamp 1677622389
transform 1 0 1464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_103
timestamp 1677622389
transform 1 0 1472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_104
timestamp 1677622389
transform 1 0 1480 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_360
timestamp 1677622389
transform 1 0 1524 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_2
timestamp 1677622389
transform -1 0 1528 0 -1 4570
box -8 -3 46 105
use FILL  FILL_105
timestamp 1677622389
transform 1 0 1528 0 -1 4570
box -8 -3 16 105
use FILL  FILL_107
timestamp 1677622389
transform 1 0 1536 0 -1 4570
box -8 -3 16 105
use FILL  FILL_109
timestamp 1677622389
transform 1 0 1544 0 -1 4570
box -8 -3 16 105
use FILL  FILL_111
timestamp 1677622389
transform 1 0 1552 0 -1 4570
box -8 -3 16 105
use FILL  FILL_113
timestamp 1677622389
transform 1 0 1560 0 -1 4570
box -8 -3 16 105
use FILL  FILL_117
timestamp 1677622389
transform 1 0 1568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_118
timestamp 1677622389
transform 1 0 1576 0 -1 4570
box -8 -3 16 105
use FILL  FILL_119
timestamp 1677622389
transform 1 0 1584 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_3
timestamp 1677622389
transform -1 0 1632 0 -1 4570
box -8 -3 46 105
use FILL  FILL_120
timestamp 1677622389
transform 1 0 1632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_121
timestamp 1677622389
transform 1 0 1640 0 -1 4570
box -8 -3 16 105
use FILL  FILL_122
timestamp 1677622389
transform 1 0 1648 0 -1 4570
box -8 -3 16 105
use FILL  FILL_123
timestamp 1677622389
transform 1 0 1656 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1677622389
transform 1 0 1664 0 -1 4570
box -9 -3 26 105
use FILL  FILL_124
timestamp 1677622389
transform 1 0 1680 0 -1 4570
box -8 -3 16 105
use FILL  FILL_126
timestamp 1677622389
transform 1 0 1688 0 -1 4570
box -8 -3 16 105
use FILL  FILL_128
timestamp 1677622389
transform 1 0 1696 0 -1 4570
box -8 -3 16 105
use FILL  FILL_130
timestamp 1677622389
transform 1 0 1704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_133
timestamp 1677622389
transform 1 0 1712 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1677622389
transform 1 0 1720 0 -1 4570
box -9 -3 26 105
use FILL  FILL_134
timestamp 1677622389
transform 1 0 1736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_136
timestamp 1677622389
transform 1 0 1744 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1677622389
transform 1 0 1752 0 -1 4570
box -8 -3 104 105
use FILL  FILL_146
timestamp 1677622389
transform 1 0 1848 0 -1 4570
box -8 -3 16 105
use FILL  FILL_147
timestamp 1677622389
transform 1 0 1856 0 -1 4570
box -8 -3 16 105
use FILL  FILL_148
timestamp 1677622389
transform 1 0 1864 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1677622389
transform 1 0 1872 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_16
timestamp 1677622389
transform -1 0 1928 0 -1 4570
box -9 -3 26 105
use FILL  FILL_149
timestamp 1677622389
transform 1 0 1928 0 -1 4570
box -8 -3 16 105
use FILL  FILL_151
timestamp 1677622389
transform 1 0 1936 0 -1 4570
box -8 -3 16 105
use FILL  FILL_157
timestamp 1677622389
transform 1 0 1944 0 -1 4570
box -8 -3 16 105
use FILL  FILL_158
timestamp 1677622389
transform 1 0 1952 0 -1 4570
box -8 -3 16 105
use FILL  FILL_159
timestamp 1677622389
transform 1 0 1960 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_11
timestamp 1677622389
transform 1 0 1968 0 -1 4570
box -8 -3 46 105
use FILL  FILL_160
timestamp 1677622389
transform 1 0 2008 0 -1 4570
box -8 -3 16 105
use FILL  FILL_161
timestamp 1677622389
transform 1 0 2016 0 -1 4570
box -8 -3 16 105
use FILL  FILL_162
timestamp 1677622389
transform 1 0 2024 0 -1 4570
box -8 -3 16 105
use FILL  FILL_163
timestamp 1677622389
transform 1 0 2032 0 -1 4570
box -8 -3 16 105
use FILL  FILL_164
timestamp 1677622389
transform 1 0 2040 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_361
timestamp 1677622389
transform 1 0 2084 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_12
timestamp 1677622389
transform -1 0 2088 0 -1 4570
box -8 -3 46 105
use FILL  FILL_165
timestamp 1677622389
transform 1 0 2088 0 -1 4570
box -8 -3 16 105
use FILL  FILL_167
timestamp 1677622389
transform 1 0 2096 0 -1 4570
box -8 -3 16 105
use FILL  FILL_169
timestamp 1677622389
transform 1 0 2104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_171
timestamp 1677622389
transform 1 0 2112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_173
timestamp 1677622389
transform 1 0 2120 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_4
timestamp 1677622389
transform 1 0 2128 0 -1 4570
box -8 -3 46 105
use FILL  FILL_178
timestamp 1677622389
transform 1 0 2168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_179
timestamp 1677622389
transform 1 0 2176 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_362
timestamp 1677622389
transform 1 0 2196 0 1 4475
box -3 -3 3 3
use FILL  FILL_180
timestamp 1677622389
transform 1 0 2184 0 -1 4570
box -8 -3 16 105
use FILL  FILL_181
timestamp 1677622389
transform 1 0 2192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_182
timestamp 1677622389
transform 1 0 2200 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_13
timestamp 1677622389
transform -1 0 2248 0 -1 4570
box -8 -3 46 105
use FILL  FILL_183
timestamp 1677622389
transform 1 0 2248 0 -1 4570
box -8 -3 16 105
use FILL  FILL_184
timestamp 1677622389
transform 1 0 2256 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_363
timestamp 1677622389
transform 1 0 2276 0 1 4475
box -3 -3 3 3
use FILL  FILL_185
timestamp 1677622389
transform 1 0 2264 0 -1 4570
box -8 -3 16 105
use FILL  FILL_187
timestamp 1677622389
transform 1 0 2272 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_14
timestamp 1677622389
transform 1 0 2280 0 -1 4570
box -8 -3 46 105
use FILL  FILL_192
timestamp 1677622389
transform 1 0 2320 0 -1 4570
box -8 -3 16 105
use FILL  FILL_194
timestamp 1677622389
transform 1 0 2328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_202
timestamp 1677622389
transform 1 0 2336 0 -1 4570
box -8 -3 16 105
use FILL  FILL_203
timestamp 1677622389
transform 1 0 2344 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1677622389
transform 1 0 2352 0 -1 4570
box -8 -3 46 105
use FILL  FILL_204
timestamp 1677622389
transform 1 0 2392 0 -1 4570
box -8 -3 16 105
use FILL  FILL_205
timestamp 1677622389
transform 1 0 2400 0 -1 4570
box -8 -3 16 105
use FILL  FILL_206
timestamp 1677622389
transform 1 0 2408 0 -1 4570
box -8 -3 16 105
use FILL  FILL_207
timestamp 1677622389
transform 1 0 2416 0 -1 4570
box -8 -3 16 105
use FILL  FILL_208
timestamp 1677622389
transform 1 0 2424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_209
timestamp 1677622389
transform 1 0 2432 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_6
timestamp 1677622389
transform 1 0 2440 0 -1 4570
box -8 -3 46 105
use FILL  FILL_210
timestamp 1677622389
transform 1 0 2480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_212
timestamp 1677622389
transform 1 0 2488 0 -1 4570
box -8 -3 16 105
use FILL  FILL_214
timestamp 1677622389
transform 1 0 2496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_216
timestamp 1677622389
transform 1 0 2504 0 -1 4570
box -8 -3 16 105
use FILL  FILL_218
timestamp 1677622389
transform 1 0 2512 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_15
timestamp 1677622389
transform 1 0 2520 0 -1 4570
box -8 -3 46 105
use M3_M2  M3_M2_364
timestamp 1677622389
transform 1 0 2572 0 1 4475
box -3 -3 3 3
use FILL  FILL_223
timestamp 1677622389
transform 1 0 2560 0 -1 4570
box -8 -3 16 105
use FILL  FILL_225
timestamp 1677622389
transform 1 0 2568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_226
timestamp 1677622389
transform 1 0 2576 0 -1 4570
box -8 -3 16 105
use FILL  FILL_227
timestamp 1677622389
transform 1 0 2584 0 -1 4570
box -8 -3 16 105
use FILL  FILL_228
timestamp 1677622389
transform 1 0 2592 0 -1 4570
box -8 -3 16 105
use FILL  FILL_229
timestamp 1677622389
transform 1 0 2600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_230
timestamp 1677622389
transform 1 0 2608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_231
timestamp 1677622389
transform 1 0 2616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_232
timestamp 1677622389
transform 1 0 2624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_233
timestamp 1677622389
transform 1 0 2632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_234
timestamp 1677622389
transform 1 0 2640 0 -1 4570
box -8 -3 16 105
use FILL  FILL_235
timestamp 1677622389
transform 1 0 2648 0 -1 4570
box -8 -3 16 105
use FILL  FILL_236
timestamp 1677622389
transform 1 0 2656 0 -1 4570
box -8 -3 16 105
use FILL  FILL_237
timestamp 1677622389
transform 1 0 2664 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_16
timestamp 1677622389
transform 1 0 2672 0 -1 4570
box -8 -3 46 105
use FILL  FILL_242
timestamp 1677622389
transform 1 0 2712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_243
timestamp 1677622389
transform 1 0 2720 0 -1 4570
box -8 -3 16 105
use FILL  FILL_244
timestamp 1677622389
transform 1 0 2728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_245
timestamp 1677622389
transform 1 0 2736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_246
timestamp 1677622389
transform 1 0 2744 0 -1 4570
box -8 -3 16 105
use FILL  FILL_247
timestamp 1677622389
transform 1 0 2752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_248
timestamp 1677622389
transform 1 0 2760 0 -1 4570
box -8 -3 16 105
use FILL  FILL_249
timestamp 1677622389
transform 1 0 2768 0 -1 4570
box -8 -3 16 105
use FILL  FILL_250
timestamp 1677622389
transform 1 0 2776 0 -1 4570
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1677622389
transform 1 0 2784 0 -1 4570
box -8 -3 32 105
use FILL  FILL_251
timestamp 1677622389
transform 1 0 2808 0 -1 4570
box -8 -3 16 105
use FILL  FILL_253
timestamp 1677622389
transform 1 0 2816 0 -1 4570
box -8 -3 16 105
use FILL  FILL_255
timestamp 1677622389
transform 1 0 2824 0 -1 4570
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1677622389
transform 1 0 2832 0 -1 4570
box -8 -3 32 105
use FILL  FILL_256
timestamp 1677622389
transform 1 0 2856 0 -1 4570
box -8 -3 16 105
use FILL  FILL_268
timestamp 1677622389
transform 1 0 2864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_269
timestamp 1677622389
transform 1 0 2872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_270
timestamp 1677622389
transform 1 0 2880 0 -1 4570
box -8 -3 16 105
use FILL  FILL_271
timestamp 1677622389
transform 1 0 2888 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1677622389
transform 1 0 2896 0 -1 4570
box -8 -3 34 105
use FILL  FILL_272
timestamp 1677622389
transform 1 0 2928 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_10
timestamp 1677622389
transform -1 0 2968 0 -1 4570
box -8 -3 34 105
use FILL  FILL_273
timestamp 1677622389
transform 1 0 2968 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1677622389
transform -1 0 3008 0 -1 4570
box -8 -3 34 105
use FILL  FILL_274
timestamp 1677622389
transform 1 0 3008 0 -1 4570
box -8 -3 16 105
use FILL  FILL_280
timestamp 1677622389
transform 1 0 3016 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_22
timestamp 1677622389
transform -1 0 3040 0 -1 4570
box -9 -3 26 105
use OAI22X1  OAI22X1_7
timestamp 1677622389
transform 1 0 3040 0 -1 4570
box -8 -3 46 105
use FILL  FILL_281
timestamp 1677622389
transform 1 0 3080 0 -1 4570
box -8 -3 16 105
use FILL  FILL_282
timestamp 1677622389
transform 1 0 3088 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_23
timestamp 1677622389
transform -1 0 3112 0 -1 4570
box -9 -3 26 105
use FILL  FILL_283
timestamp 1677622389
transform 1 0 3112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_284
timestamp 1677622389
transform 1 0 3120 0 -1 4570
box -8 -3 16 105
use FILL  FILL_285
timestamp 1677622389
transform 1 0 3128 0 -1 4570
box -8 -3 16 105
use FILL  FILL_286
timestamp 1677622389
transform 1 0 3136 0 -1 4570
box -8 -3 16 105
use FILL  FILL_287
timestamp 1677622389
transform 1 0 3144 0 -1 4570
box -8 -3 16 105
use FILL  FILL_289
timestamp 1677622389
transform 1 0 3152 0 -1 4570
box -8 -3 16 105
use FILL  FILL_291
timestamp 1677622389
transform 1 0 3160 0 -1 4570
box -8 -3 16 105
use FILL  FILL_293
timestamp 1677622389
transform 1 0 3168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_295
timestamp 1677622389
transform 1 0 3176 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_8
timestamp 1677622389
transform 1 0 3184 0 -1 4570
box -8 -3 46 105
use FILL  FILL_302
timestamp 1677622389
transform 1 0 3224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_303
timestamp 1677622389
transform 1 0 3232 0 -1 4570
box -8 -3 16 105
use FILL  FILL_304
timestamp 1677622389
transform 1 0 3240 0 -1 4570
box -8 -3 16 105
use FILL  FILL_305
timestamp 1677622389
transform 1 0 3248 0 -1 4570
box -8 -3 16 105
use FILL  FILL_306
timestamp 1677622389
transform 1 0 3256 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1677622389
transform -1 0 3304 0 -1 4570
box -8 -3 46 105
use FILL  FILL_307
timestamp 1677622389
transform 1 0 3304 0 -1 4570
box -8 -3 16 105
use FILL  FILL_308
timestamp 1677622389
transform 1 0 3312 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_25
timestamp 1677622389
transform -1 0 3336 0 -1 4570
box -9 -3 26 105
use NAND3X1  NAND3X1_0
timestamp 1677622389
transform -1 0 3368 0 -1 4570
box -8 -3 40 105
use FILL  FILL_309
timestamp 1677622389
transform 1 0 3368 0 -1 4570
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1677622389
transform -1 0 3408 0 -1 4570
box -8 -3 40 105
use FILL  FILL_310
timestamp 1677622389
transform 1 0 3408 0 -1 4570
box -8 -3 16 105
use FILL  FILL_311
timestamp 1677622389
transform 1 0 3416 0 -1 4570
box -8 -3 16 105
use FILL  FILL_312
timestamp 1677622389
transform 1 0 3424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_313
timestamp 1677622389
transform 1 0 3432 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_26
timestamp 1677622389
transform 1 0 3440 0 -1 4570
box -9 -3 26 105
use FILL  FILL_316
timestamp 1677622389
transform 1 0 3456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_317
timestamp 1677622389
transform 1 0 3464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_318
timestamp 1677622389
transform 1 0 3472 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_10
timestamp 1677622389
transform 1 0 3480 0 -1 4570
box -8 -3 46 105
use FILL  FILL_319
timestamp 1677622389
transform 1 0 3520 0 -1 4570
box -8 -3 16 105
use FILL  FILL_320
timestamp 1677622389
transform 1 0 3528 0 -1 4570
box -8 -3 16 105
use FILL  FILL_321
timestamp 1677622389
transform 1 0 3536 0 -1 4570
box -8 -3 16 105
use FILL  FILL_322
timestamp 1677622389
transform 1 0 3544 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_365
timestamp 1677622389
transform 1 0 3588 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_11
timestamp 1677622389
transform 1 0 3552 0 -1 4570
box -8 -3 46 105
use FILL  FILL_326
timestamp 1677622389
transform 1 0 3592 0 -1 4570
box -8 -3 16 105
use FILL  FILL_327
timestamp 1677622389
transform 1 0 3600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_328
timestamp 1677622389
transform 1 0 3608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_329
timestamp 1677622389
transform 1 0 3616 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_366
timestamp 1677622389
transform 1 0 3636 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_17
timestamp 1677622389
transform -1 0 3664 0 -1 4570
box -8 -3 46 105
use FILL  FILL_330
timestamp 1677622389
transform 1 0 3664 0 -1 4570
box -8 -3 16 105
use FILL  FILL_331
timestamp 1677622389
transform 1 0 3672 0 -1 4570
box -8 -3 16 105
use FILL  FILL_332
timestamp 1677622389
transform 1 0 3680 0 -1 4570
box -8 -3 16 105
use FILL  FILL_337
timestamp 1677622389
transform 1 0 3688 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_18
timestamp 1677622389
transform -1 0 3736 0 -1 4570
box -8 -3 46 105
use FILL  FILL_338
timestamp 1677622389
transform 1 0 3736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_339
timestamp 1677622389
transform 1 0 3744 0 -1 4570
box -8 -3 16 105
use FILL  FILL_340
timestamp 1677622389
transform 1 0 3752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_341
timestamp 1677622389
transform 1 0 3760 0 -1 4570
box -8 -3 16 105
use FILL  FILL_342
timestamp 1677622389
transform 1 0 3768 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_12
timestamp 1677622389
transform 1 0 3776 0 -1 4570
box -8 -3 46 105
use FILL  FILL_343
timestamp 1677622389
transform 1 0 3816 0 -1 4570
box -8 -3 16 105
use FILL  FILL_344
timestamp 1677622389
transform 1 0 3824 0 -1 4570
box -8 -3 16 105
use FILL  FILL_346
timestamp 1677622389
transform 1 0 3832 0 -1 4570
box -8 -3 16 105
use FILL  FILL_349
timestamp 1677622389
transform 1 0 3840 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_13
timestamp 1677622389
transform -1 0 3888 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1677622389
transform 1 0 3888 0 -1 4570
box -8 -3 46 105
use FILL  FILL_350
timestamp 1677622389
transform 1 0 3928 0 -1 4570
box -8 -3 16 105
use FILL  FILL_351
timestamp 1677622389
transform 1 0 3936 0 -1 4570
box -8 -3 16 105
use FILL  FILL_352
timestamp 1677622389
transform 1 0 3944 0 -1 4570
box -8 -3 16 105
use FILL  FILL_357
timestamp 1677622389
transform 1 0 3952 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_30
timestamp 1677622389
transform -1 0 3976 0 -1 4570
box -9 -3 26 105
use FILL  FILL_358
timestamp 1677622389
transform 1 0 3976 0 -1 4570
box -8 -3 16 105
use FILL  FILL_359
timestamp 1677622389
transform 1 0 3984 0 -1 4570
box -8 -3 16 105
use FILL  FILL_360
timestamp 1677622389
transform 1 0 3992 0 -1 4570
box -8 -3 16 105
use FILL  FILL_361
timestamp 1677622389
transform 1 0 4000 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_14
timestamp 1677622389
transform -1 0 4048 0 -1 4570
box -8 -3 46 105
use FILL  FILL_362
timestamp 1677622389
transform 1 0 4048 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1677622389
transform 1 0 4056 0 -1 4570
box -9 -3 26 105
use FILL  FILL_363
timestamp 1677622389
transform 1 0 4072 0 -1 4570
box -8 -3 16 105
use FILL  FILL_364
timestamp 1677622389
transform 1 0 4080 0 -1 4570
box -8 -3 16 105
use FILL  FILL_365
timestamp 1677622389
transform 1 0 4088 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_32
timestamp 1677622389
transform -1 0 4112 0 -1 4570
box -9 -3 26 105
use FILL  FILL_366
timestamp 1677622389
transform 1 0 4112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_367
timestamp 1677622389
transform 1 0 4120 0 -1 4570
box -8 -3 16 105
use FILL  FILL_368
timestamp 1677622389
transform 1 0 4128 0 -1 4570
box -8 -3 16 105
use FILL  FILL_369
timestamp 1677622389
transform 1 0 4136 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_15
timestamp 1677622389
transform 1 0 4144 0 -1 4570
box -8 -3 46 105
use FILL  FILL_370
timestamp 1677622389
transform 1 0 4184 0 -1 4570
box -8 -3 16 105
use FILL  FILL_372
timestamp 1677622389
transform 1 0 4192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_374
timestamp 1677622389
transform 1 0 4200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_376
timestamp 1677622389
transform 1 0 4208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_377
timestamp 1677622389
transform 1 0 4216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_378
timestamp 1677622389
transform 1 0 4224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_379
timestamp 1677622389
transform 1 0 4232 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_16
timestamp 1677622389
transform 1 0 4240 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_33
timestamp 1677622389
transform -1 0 4296 0 -1 4570
box -9 -3 26 105
use FILL  FILL_380
timestamp 1677622389
transform 1 0 4296 0 -1 4570
box -8 -3 16 105
use FILL  FILL_381
timestamp 1677622389
transform 1 0 4304 0 -1 4570
box -8 -3 16 105
use FILL  FILL_383
timestamp 1677622389
transform 1 0 4312 0 -1 4570
box -8 -3 16 105
use FILL  FILL_387
timestamp 1677622389
transform 1 0 4320 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_20
timestamp 1677622389
transform -1 0 4368 0 -1 4570
box -8 -3 46 105
use FILL  FILL_388
timestamp 1677622389
transform 1 0 4368 0 -1 4570
box -8 -3 16 105
use FILL  FILL_389
timestamp 1677622389
transform 1 0 4376 0 -1 4570
box -8 -3 16 105
use FILL  FILL_390
timestamp 1677622389
transform 1 0 4384 0 -1 4570
box -8 -3 16 105
use FILL  FILL_391
timestamp 1677622389
transform 1 0 4392 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_17
timestamp 1677622389
transform 1 0 4400 0 -1 4570
box -8 -3 46 105
use FILL  FILL_392
timestamp 1677622389
transform 1 0 4440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_393
timestamp 1677622389
transform 1 0 4448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_395
timestamp 1677622389
transform 1 0 4456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_397
timestamp 1677622389
transform 1 0 4464 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1677622389
transform 1 0 4472 0 -1 4570
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1677622389
transform 1 0 4568 0 -1 4570
box -9 -3 26 105
use OAI22X1  OAI22X1_19
timestamp 1677622389
transform 1 0 4584 0 -1 4570
box -8 -3 46 105
use FILL  FILL_409
timestamp 1677622389
transform 1 0 4624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_410
timestamp 1677622389
transform 1 0 4632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_411
timestamp 1677622389
transform 1 0 4640 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_36
timestamp 1677622389
transform 1 0 4648 0 -1 4570
box -9 -3 26 105
use OAI22X1  OAI22X1_20
timestamp 1677622389
transform 1 0 4664 0 -1 4570
box -8 -3 46 105
use FILL  FILL_412
timestamp 1677622389
transform 1 0 4704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_413
timestamp 1677622389
transform 1 0 4712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_414
timestamp 1677622389
transform 1 0 4720 0 -1 4570
box -8 -3 16 105
use FILL  FILL_415
timestamp 1677622389
transform 1 0 4728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_416
timestamp 1677622389
transform 1 0 4736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_417
timestamp 1677622389
transform 1 0 4744 0 -1 4570
box -8 -3 16 105
use FILL  FILL_418
timestamp 1677622389
transform 1 0 4752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_419
timestamp 1677622389
transform 1 0 4760 0 -1 4570
box -8 -3 16 105
use FILL  FILL_420
timestamp 1677622389
transform 1 0 4768 0 -1 4570
box -8 -3 16 105
use FILL  FILL_421
timestamp 1677622389
transform 1 0 4776 0 -1 4570
box -8 -3 16 105
use FILL  FILL_422
timestamp 1677622389
transform 1 0 4784 0 -1 4570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_5
timestamp 1677622389
transform 1 0 4843 0 1 4470
box -10 -3 10 3
use M2_M1  M2_M1_448
timestamp 1677622389
transform 1 0 116 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1677622389
transform 1 0 92 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1677622389
transform 1 0 92 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1677622389
transform 1 0 180 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1677622389
transform 1 0 196 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_449
timestamp 1677622389
transform 1 0 196 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_410
timestamp 1677622389
transform 1 0 236 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_450
timestamp 1677622389
transform 1 0 212 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1677622389
transform 1 0 228 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1677622389
transform 1 0 220 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1677622389
transform 1 0 236 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_494
timestamp 1677622389
transform 1 0 220 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1677622389
transform 1 0 236 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1677622389
transform 1 0 356 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_452
timestamp 1677622389
transform 1 0 308 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1677622389
transform 1 0 356 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1677622389
transform 1 0 276 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1677622389
transform 1 0 276 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1677622389
transform 1 0 484 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1677622389
transform 1 0 460 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_454
timestamp 1677622389
transform 1 0 404 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_451
timestamp 1677622389
transform 1 0 412 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_455
timestamp 1677622389
transform 1 0 460 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1677622389
transform 1 0 484 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1677622389
transform 1 0 412 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1677622389
transform 1 0 508 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1677622389
transform 1 0 500 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_456
timestamp 1677622389
transform 1 0 500 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1677622389
transform 1 0 540 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1677622389
transform 1 0 532 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_457
timestamp 1677622389
transform 1 0 540 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1677622389
transform 1 0 556 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_458
timestamp 1677622389
transform 1 0 564 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_452
timestamp 1677622389
transform 1 0 572 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1677622389
transform 1 0 580 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1677622389
transform 1 0 588 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1677622389
transform 1 0 548 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1677622389
transform 1 0 556 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1677622389
transform 1 0 572 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1677622389
transform 1 0 604 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1677622389
transform 1 0 612 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1677622389
transform 1 0 652 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1677622389
transform 1 0 628 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1677622389
transform 1 0 676 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1677622389
transform 1 0 668 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1677622389
transform 1 0 660 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_461
timestamp 1677622389
transform 1 0 628 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1677622389
transform 1 0 644 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_453
timestamp 1677622389
transform 1 0 652 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_463
timestamp 1677622389
transform 1 0 660 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1677622389
transform 1 0 636 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_472
timestamp 1677622389
transform 1 0 644 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_583
timestamp 1677622389
transform 1 0 652 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1677622389
transform 1 0 676 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_396
timestamp 1677622389
transform 1 0 708 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1677622389
transform 1 0 692 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_464
timestamp 1677622389
transform 1 0 708 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_455
timestamp 1677622389
transform 1 0 716 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_585
timestamp 1677622389
transform 1 0 700 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1677622389
transform 1 0 716 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1677622389
transform 1 0 700 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1677622389
transform 1 0 740 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_587
timestamp 1677622389
transform 1 0 740 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1677622389
transform 1 0 764 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1677622389
transform 1 0 780 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_465
timestamp 1677622389
transform 1 0 756 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1677622389
transform 1 0 764 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1677622389
transform 1 0 780 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1677622389
transform 1 0 796 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1677622389
transform 1 0 756 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1677622389
transform 1 0 772 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1677622389
transform 1 0 812 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1677622389
transform 1 0 868 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1677622389
transform 1 0 836 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1677622389
transform 1 0 932 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_473
timestamp 1677622389
transform 1 0 924 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_669
timestamp 1677622389
transform 1 0 924 0 1 4395
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1677622389
transform 1 0 972 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1677622389
transform 1 0 988 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1677622389
transform 1 0 988 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1677622389
transform 1 0 980 0 1 4395
box -2 -2 2 2
use M3_M2  M3_M2_535
timestamp 1677622389
transform 1 0 980 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1677622389
transform 1 0 1044 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_472
timestamp 1677622389
transform 1 0 1044 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1677622389
transform 1 0 1052 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1677622389
transform 1 0 1060 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1677622389
transform 1 0 1100 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1677622389
transform 1 0 1084 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1677622389
transform 1 0 1092 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1677622389
transform 1 0 1108 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_495
timestamp 1677622389
transform 1 0 1116 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_671
timestamp 1677622389
transform 1 0 1124 0 1 4395
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1677622389
transform 1 0 1132 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1677622389
transform 1 0 1164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1677622389
transform 1 0 1180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1677622389
transform 1 0 1156 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_474
timestamp 1677622389
transform 1 0 1164 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_598
timestamp 1677622389
transform 1 0 1172 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1677622389
transform 1 0 1188 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1677622389
transform 1 0 1204 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_599
timestamp 1677622389
transform 1 0 1196 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1677622389
transform 1 0 1236 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1677622389
transform 1 0 1252 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1677622389
transform 1 0 1300 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1677622389
transform 1 0 1308 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1677622389
transform 1 0 1308 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1677622389
transform 1 0 1332 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1677622389
transform 1 0 1356 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_481
timestamp 1677622389
transform 1 0 1364 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1677622389
transform 1 0 1420 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1677622389
transform 1 0 1356 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_476
timestamp 1677622389
transform 1 0 1420 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_603
timestamp 1677622389
transform 1 0 1444 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1677622389
transform 1 0 1460 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1677622389
transform 1 0 1476 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_496
timestamp 1677622389
transform 1 0 1476 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1677622389
transform 1 0 1492 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1677622389
transform 1 0 1540 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_484
timestamp 1677622389
transform 1 0 1508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1677622389
transform 1 0 1516 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1677622389
transform 1 0 1508 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1677622389
transform 1 0 1540 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1677622389
transform 1 0 1556 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1677622389
transform 1 0 1516 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1677622389
transform 1 0 1532 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1677622389
transform 1 0 1548 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1677622389
transform 1 0 1556 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1677622389
transform 1 0 1644 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_488
timestamp 1677622389
transform 1 0 1604 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1677622389
transform 1 0 1660 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1677622389
transform 1 0 1564 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1677622389
transform 1 0 1580 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1677622389
transform 1 0 1532 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1677622389
transform 1 0 1548 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1677622389
transform 1 0 1604 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1677622389
transform 1 0 1564 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1677622389
transform 1 0 1668 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1677622389
transform 1 0 1692 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1677622389
transform 1 0 1684 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1677622389
transform 1 0 1748 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1677622389
transform 1 0 1700 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_490
timestamp 1677622389
transform 1 0 1748 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_457
timestamp 1677622389
transform 1 0 1764 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1677622389
transform 1 0 1788 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_491
timestamp 1677622389
transform 1 0 1780 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1677622389
transform 1 0 1788 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1677622389
transform 1 0 1700 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1677622389
transform 1 0 1780 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_493
timestamp 1677622389
transform 1 0 1804 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1677622389
transform 1 0 1804 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1677622389
transform 1 0 1860 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1677622389
transform 1 0 1844 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1677622389
transform 1 0 1852 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1677622389
transform 1 0 1868 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_501
timestamp 1677622389
transform 1 0 1868 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1677622389
transform 1 0 1884 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_495
timestamp 1677622389
transform 1 0 1884 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1677622389
transform 1 0 1908 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1677622389
transform 1 0 1932 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_496
timestamp 1677622389
transform 1 0 1916 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1677622389
transform 1 0 1932 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1677622389
transform 1 0 1924 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_429
timestamp 1677622389
transform 1 0 1948 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_498
timestamp 1677622389
transform 1 0 1956 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_458
timestamp 1677622389
transform 1 0 1964 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_615
timestamp 1677622389
transform 1 0 1964 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1677622389
transform 1 0 2012 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1677622389
transform 1 0 2052 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_502
timestamp 1677622389
transform 1 0 2052 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_500
timestamp 1677622389
transform 1 0 2068 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_482
timestamp 1677622389
transform 1 0 2068 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_617
timestamp 1677622389
transform 1 0 2092 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_538
timestamp 1677622389
transform 1 0 2092 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1677622389
transform 1 0 2124 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_501
timestamp 1677622389
transform 1 0 2116 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_459
timestamp 1677622389
transform 1 0 2124 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1677622389
transform 1 0 2140 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_502
timestamp 1677622389
transform 1 0 2140 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1677622389
transform 1 0 2124 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1677622389
transform 1 0 2132 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_385
timestamp 1677622389
transform 1 0 2156 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1677622389
transform 1 0 2180 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1677622389
transform 1 0 2188 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1677622389
transform 1 0 2180 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1677622389
transform 1 0 2284 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1677622389
transform 1 0 2220 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1677622389
transform 1 0 2316 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1677622389
transform 1 0 2180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1677622389
transform 1 0 2188 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1677622389
transform 1 0 2220 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1677622389
transform 1 0 2284 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1677622389
transform 1 0 2300 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1677622389
transform 1 0 2172 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1677622389
transform 1 0 2308 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_508
timestamp 1677622389
transform 1 0 2316 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1677622389
transform 1 0 2268 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1677622389
transform 1 0 2284 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1677622389
transform 1 0 2292 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1677622389
transform 1 0 2308 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1677622389
transform 1 0 2316 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1677622389
transform 1 0 2268 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1677622389
transform 1 0 2284 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1677622389
transform 1 0 2340 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1677622389
transform 1 0 2380 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_509
timestamp 1677622389
transform 1 0 2380 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1677622389
transform 1 0 2428 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1677622389
transform 1 0 2420 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1677622389
transform 1 0 2420 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_461
timestamp 1677622389
transform 1 0 2468 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_511
timestamp 1677622389
transform 1 0 2476 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1677622389
transform 1 0 2396 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1677622389
transform 1 0 2396 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1677622389
transform 1 0 2428 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1677622389
transform 1 0 2460 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1677622389
transform 1 0 2508 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1677622389
transform 1 0 2548 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_512
timestamp 1677622389
transform 1 0 2508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1677622389
transform 1 0 2516 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1677622389
transform 1 0 2532 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1677622389
transform 1 0 2540 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_515
timestamp 1677622389
transform 1 0 2548 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_483
timestamp 1677622389
transform 1 0 2516 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_626
timestamp 1677622389
transform 1 0 2524 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1677622389
transform 1 0 2540 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1677622389
transform 1 0 2548 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1677622389
transform 1 0 2516 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1677622389
transform 1 0 2564 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1677622389
transform 1 0 2580 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1677622389
transform 1 0 2580 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_437
timestamp 1677622389
transform 1 0 2620 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_517
timestamp 1677622389
transform 1 0 2620 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1677622389
transform 1 0 2668 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_518
timestamp 1677622389
transform 1 0 2676 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1677622389
transform 1 0 2596 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_401
timestamp 1677622389
transform 1 0 2692 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_519
timestamp 1677622389
transform 1 0 2692 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1677622389
transform 1 0 2684 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1677622389
transform 1 0 2596 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1677622389
transform 1 0 2676 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1677622389
transform 1 0 2724 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1677622389
transform 1 0 2716 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1677622389
transform 1 0 2740 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1677622389
transform 1 0 2724 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1677622389
transform 1 0 2732 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_367
timestamp 1677622389
transform 1 0 2828 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1677622389
transform 1 0 2844 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1677622389
transform 1 0 2868 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1677622389
transform 1 0 2748 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1677622389
transform 1 0 2788 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1677622389
transform 1 0 2836 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_442
timestamp 1677622389
transform 1 0 2876 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_441
timestamp 1677622389
transform 1 0 2884 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_522
timestamp 1677622389
transform 1 0 2748 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1677622389
transform 1 0 2788 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1677622389
transform 1 0 2844 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1677622389
transform 1 0 2860 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1677622389
transform 1 0 2764 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1677622389
transform 1 0 2852 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_508
timestamp 1677622389
transform 1 0 2804 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1677622389
transform 1 0 2852 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1677622389
transform 1 0 2884 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1677622389
transform 1 0 2892 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1677622389
transform 1 0 2884 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1677622389
transform 1 0 2876 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_443
timestamp 1677622389
transform 1 0 2916 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_464
timestamp 1677622389
transform 1 0 2916 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1677622389
transform 1 0 2908 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1677622389
transform 1 0 2884 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1677622389
transform 1 0 2916 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_484
timestamp 1677622389
transform 1 0 2924 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_672
timestamp 1677622389
transform 1 0 2924 0 1 4395
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1677622389
transform 1 0 2948 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1677622389
transform 1 0 2940 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_465
timestamp 1677622389
transform 1 0 2948 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1677622389
transform 1 0 2940 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1677622389
transform 1 0 2948 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1677622389
transform 1 0 2940 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1677622389
transform 1 0 2980 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1677622389
transform 1 0 2972 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_445
timestamp 1677622389
transform 1 0 2988 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1677622389
transform 1 0 2972 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1677622389
transform 1 0 2980 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_443
timestamp 1677622389
transform 1 0 3004 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1677622389
transform 1 0 3004 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1677622389
transform 1 0 2980 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_485
timestamp 1677622389
transform 1 0 2988 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1677622389
transform 1 0 3036 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_640
timestamp 1677622389
transform 1 0 3020 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1677622389
transform 1 0 3028 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1677622389
transform 1 0 3076 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_532
timestamp 1677622389
transform 1 0 3044 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1677622389
transform 1 0 3060 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1677622389
transform 1 0 3076 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1677622389
transform 1 0 3108 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1677622389
transform 1 0 3036 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1677622389
transform 1 0 3052 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1677622389
transform 1 0 3060 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1677622389
transform 1 0 3156 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_643
timestamp 1677622389
transform 1 0 3068 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1677622389
transform 1 0 3156 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_512
timestamp 1677622389
transform 1 0 3052 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1677622389
transform 1 0 3108 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1677622389
transform 1 0 3188 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1677622389
transform 1 0 3308 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1677622389
transform 1 0 3340 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1677622389
transform 1 0 3284 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1677622389
transform 1 0 3356 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1677622389
transform 1 0 3212 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1677622389
transform 1 0 3268 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1677622389
transform 1 0 3332 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1677622389
transform 1 0 3364 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1677622389
transform 1 0 3188 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_514
timestamp 1677622389
transform 1 0 3188 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1677622389
transform 1 0 3212 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_646
timestamp 1677622389
transform 1 0 3284 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1677622389
transform 1 0 3332 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1677622389
transform 1 0 3348 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_446
timestamp 1677622389
transform 1 0 3404 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_368
timestamp 1677622389
transform 1 0 3420 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1677622389
transform 1 0 3420 0 1 4435
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1677622389
transform 1 0 3428 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1677622389
transform 1 0 3444 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_447
timestamp 1677622389
transform 1 0 3444 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1677622389
transform 1 0 3436 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1677622389
transform 1 0 3428 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1677622389
transform 1 0 3532 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_541
timestamp 1677622389
transform 1 0 3452 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1677622389
transform 1 0 3508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1677622389
transform 1 0 3532 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_518
timestamp 1677622389
transform 1 0 3508 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1677622389
transform 1 0 3548 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1677622389
transform 1 0 3572 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_543
timestamp 1677622389
transform 1 0 3628 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_468
timestamp 1677622389
transform 1 0 3636 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1677622389
transform 1 0 3684 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1677622389
transform 1 0 3604 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1677622389
transform 1 0 3772 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1677622389
transform 1 0 3724 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_520
timestamp 1677622389
transform 1 0 3772 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1677622389
transform 1 0 3804 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_546
timestamp 1677622389
transform 1 0 3836 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_382
timestamp 1677622389
transform 1 0 3908 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1677622389
transform 1 0 3932 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_547
timestamp 1677622389
transform 1 0 3892 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1677622389
transform 1 0 3908 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1677622389
transform 1 0 3924 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1677622389
transform 1 0 3900 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1677622389
transform 1 0 3932 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1677622389
transform 1 0 3940 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1677622389
transform 1 0 3940 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_652
timestamp 1677622389
transform 1 0 3948 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_445
timestamp 1677622389
transform 1 0 4004 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_551
timestamp 1677622389
transform 1 0 4004 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_469
timestamp 1677622389
transform 1 0 4012 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_653
timestamp 1677622389
transform 1 0 3996 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1677622389
transform 1 0 4012 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_522
timestamp 1677622389
transform 1 0 3996 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1677622389
transform 1 0 4020 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1677622389
transform 1 0 4036 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1677622389
transform 1 0 4084 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_552
timestamp 1677622389
transform 1 0 4084 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1677622389
transform 1 0 4140 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1677622389
transform 1 0 4060 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_523
timestamp 1677622389
transform 1 0 4084 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1677622389
transform 1 0 4148 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1677622389
transform 1 0 4220 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1677622389
transform 1 0 4212 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1677622389
transform 1 0 4252 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1677622389
transform 1 0 4172 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_369
timestamp 1677622389
transform 1 0 4348 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1677622389
transform 1 0 4300 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_556
timestamp 1677622389
transform 1 0 4340 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1677622389
transform 1 0 4300 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_447
timestamp 1677622389
transform 1 0 4396 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_557
timestamp 1677622389
transform 1 0 4396 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_389
timestamp 1677622389
transform 1 0 4428 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1677622389
transform 1 0 4444 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1677622389
transform 1 0 4412 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1677622389
transform 1 0 4428 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1677622389
transform 1 0 4444 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1677622389
transform 1 0 4420 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1677622389
transform 1 0 4460 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_548
timestamp 1677622389
transform 1 0 4460 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1677622389
transform 1 0 4476 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1677622389
transform 1 0 4508 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1677622389
transform 1 0 4492 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1677622389
transform 1 0 4508 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1677622389
transform 1 0 4476 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1677622389
transform 1 0 4484 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1677622389
transform 1 0 4500 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1677622389
transform 1 0 4516 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1677622389
transform 1 0 4484 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1677622389
transform 1 0 4500 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1677622389
transform 1 0 4564 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1677622389
transform 1 0 4580 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1677622389
transform 1 0 4668 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1677622389
transform 1 0 4636 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_565
timestamp 1677622389
transform 1 0 4636 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1677622389
transform 1 0 4644 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1677622389
transform 1 0 4668 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1677622389
transform 1 0 4540 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1677622389
transform 1 0 4620 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1677622389
transform 1 0 4636 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1677622389
transform 1 0 4692 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1677622389
transform 1 0 4708 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1677622389
transform 1 0 4716 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1677622389
transform 1 0 4772 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1677622389
transform 1 0 4788 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1677622389
transform 1 0 4644 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1677622389
transform 1 0 4660 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1677622389
transform 1 0 4676 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1677622389
transform 1 0 4692 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1677622389
transform 1 0 4780 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1677622389
transform 1 0 4564 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1677622389
transform 1 0 4540 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1677622389
transform 1 0 4572 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1677622389
transform 1 0 4660 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1677622389
transform 1 0 4716 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1677622389
transform 1 0 4676 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1677622389
transform 1 0 4724 0 1 4385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_6
timestamp 1677622389
transform 1 0 48 0 1 4370
box -10 -3 10 3
use FILL  FILL_423
timestamp 1677622389
transform 1 0 72 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1677622389
transform 1 0 80 0 1 4370
box -8 -3 104 105
use FILL  FILL_425
timestamp 1677622389
transform 1 0 176 0 1 4370
box -8 -3 16 105
use FILL  FILL_439
timestamp 1677622389
transform 1 0 184 0 1 4370
box -8 -3 16 105
use FILL  FILL_441
timestamp 1677622389
transform 1 0 192 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_21
timestamp 1677622389
transform 1 0 200 0 1 4370
box -8 -3 46 105
use FILL  FILL_443
timestamp 1677622389
transform 1 0 240 0 1 4370
box -8 -3 16 105
use FILL  FILL_445
timestamp 1677622389
transform 1 0 248 0 1 4370
box -8 -3 16 105
use FILL  FILL_447
timestamp 1677622389
transform 1 0 256 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1677622389
transform 1 0 264 0 1 4370
box -8 -3 104 105
use FILL  FILL_449
timestamp 1677622389
transform 1 0 360 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_553
timestamp 1677622389
transform 1 0 380 0 1 4375
box -3 -3 3 3
use FILL  FILL_450
timestamp 1677622389
transform 1 0 368 0 1 4370
box -8 -3 16 105
use FILL  FILL_451
timestamp 1677622389
transform 1 0 376 0 1 4370
box -8 -3 16 105
use FILL  FILL_452
timestamp 1677622389
transform 1 0 384 0 1 4370
box -8 -3 16 105
use FILL  FILL_460
timestamp 1677622389
transform 1 0 392 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1677622389
transform -1 0 496 0 1 4370
box -8 -3 104 105
use FILL  FILL_461
timestamp 1677622389
transform 1 0 496 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_39
timestamp 1677622389
transform -1 0 520 0 1 4370
box -9 -3 26 105
use FILL  FILL_464
timestamp 1677622389
transform 1 0 520 0 1 4370
box -8 -3 16 105
use FILL  FILL_466
timestamp 1677622389
transform 1 0 528 0 1 4370
box -8 -3 16 105
use FILL  FILL_468
timestamp 1677622389
transform 1 0 536 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_22
timestamp 1677622389
transform 1 0 544 0 1 4370
box -8 -3 46 105
use FILL  FILL_469
timestamp 1677622389
transform 1 0 584 0 1 4370
box -8 -3 16 105
use FILL  FILL_472
timestamp 1677622389
transform 1 0 592 0 1 4370
box -8 -3 16 105
use FILL  FILL_474
timestamp 1677622389
transform 1 0 600 0 1 4370
box -8 -3 16 105
use FILL  FILL_476
timestamp 1677622389
transform 1 0 608 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_23
timestamp 1677622389
transform 1 0 616 0 1 4370
box -8 -3 46 105
use FILL  FILL_478
timestamp 1677622389
transform 1 0 656 0 1 4370
box -8 -3 16 105
use FILL  FILL_479
timestamp 1677622389
transform 1 0 664 0 1 4370
box -8 -3 16 105
use FILL  FILL_480
timestamp 1677622389
transform 1 0 672 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_24
timestamp 1677622389
transform 1 0 680 0 1 4370
box -8 -3 46 105
use FILL  FILL_482
timestamp 1677622389
transform 1 0 720 0 1 4370
box -8 -3 16 105
use FILL  FILL_483
timestamp 1677622389
transform 1 0 728 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1677622389
transform 1 0 736 0 1 4370
box -9 -3 26 105
use FILL  FILL_484
timestamp 1677622389
transform 1 0 752 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_25
timestamp 1677622389
transform 1 0 760 0 1 4370
box -8 -3 46 105
use FILL  FILL_485
timestamp 1677622389
transform 1 0 800 0 1 4370
box -8 -3 16 105
use FILL  FILL_490
timestamp 1677622389
transform 1 0 808 0 1 4370
box -8 -3 16 105
use FILL  FILL_492
timestamp 1677622389
transform 1 0 816 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1677622389
transform 1 0 824 0 1 4370
box -8 -3 104 105
use FILL  FILL_493
timestamp 1677622389
transform 1 0 920 0 1 4370
box -8 -3 16 105
use FILL  FILL_494
timestamp 1677622389
transform 1 0 928 0 1 4370
box -8 -3 16 105
use FILL  FILL_495
timestamp 1677622389
transform 1 0 936 0 1 4370
box -8 -3 16 105
use FILL  FILL_496
timestamp 1677622389
transform 1 0 944 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1677622389
transform 1 0 952 0 1 4370
box -8 -3 32 105
use FILL  FILL_502
timestamp 1677622389
transform 1 0 976 0 1 4370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1677622389
transform 1 0 984 0 1 4370
box -8 -3 16 105
use FILL  FILL_508
timestamp 1677622389
transform 1 0 992 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1677622389
transform 1 0 1000 0 1 4370
box -8 -3 32 105
use FILL  FILL_509
timestamp 1677622389
transform 1 0 1024 0 1 4370
box -8 -3 16 105
use FILL  FILL_512
timestamp 1677622389
transform 1 0 1032 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_554
timestamp 1677622389
transform 1 0 1060 0 1 4375
box -3 -3 3 3
use FILL  FILL_514
timestamp 1677622389
transform 1 0 1040 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1677622389
transform -1 0 1064 0 1 4370
box -9 -3 26 105
use FILL  FILL_515
timestamp 1677622389
transform 1 0 1064 0 1 4370
box -8 -3 16 105
use FILL  FILL_516
timestamp 1677622389
transform 1 0 1072 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_27
timestamp 1677622389
transform 1 0 1080 0 1 4370
box -8 -3 46 105
use FILL  FILL_517
timestamp 1677622389
transform 1 0 1120 0 1 4370
box -8 -3 16 105
use FILL  FILL_526
timestamp 1677622389
transform 1 0 1128 0 1 4370
box -8 -3 16 105
use FILL  FILL_527
timestamp 1677622389
transform 1 0 1136 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_555
timestamp 1677622389
transform 1 0 1156 0 1 4375
box -3 -3 3 3
use NOR2X1  NOR2X1_6
timestamp 1677622389
transform 1 0 1144 0 1 4370
box -8 -3 32 105
use M3_M2  M3_M2_556
timestamp 1677622389
transform 1 0 1204 0 1 4375
box -3 -3 3 3
use OAI21X1  OAI21X1_13
timestamp 1677622389
transform 1 0 1168 0 1 4370
box -8 -3 34 105
use FILL  FILL_528
timestamp 1677622389
transform 1 0 1200 0 1 4370
box -8 -3 16 105
use FILL  FILL_529
timestamp 1677622389
transform 1 0 1208 0 1 4370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1677622389
transform 1 0 1216 0 1 4370
box -8 -3 16 105
use FILL  FILL_531
timestamp 1677622389
transform 1 0 1224 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_14
timestamp 1677622389
transform -1 0 1264 0 1 4370
box -8 -3 34 105
use FILL  FILL_532
timestamp 1677622389
transform 1 0 1264 0 1 4370
box -8 -3 16 105
use FILL  FILL_533
timestamp 1677622389
transform 1 0 1272 0 1 4370
box -8 -3 16 105
use FILL  FILL_534
timestamp 1677622389
transform 1 0 1280 0 1 4370
box -8 -3 16 105
use FILL  FILL_535
timestamp 1677622389
transform 1 0 1288 0 1 4370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1677622389
transform 1 0 1296 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_15
timestamp 1677622389
transform -1 0 1336 0 1 4370
box -8 -3 34 105
use FILL  FILL_537
timestamp 1677622389
transform 1 0 1336 0 1 4370
box -8 -3 16 105
use FILL  FILL_538
timestamp 1677622389
transform 1 0 1344 0 1 4370
box -8 -3 16 105
use FILL  FILL_539
timestamp 1677622389
transform 1 0 1352 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1677622389
transform -1 0 1456 0 1 4370
box -8 -3 104 105
use FILL  FILL_540
timestamp 1677622389
transform 1 0 1456 0 1 4370
box -8 -3 16 105
use FILL  FILL_561
timestamp 1677622389
transform 1 0 1464 0 1 4370
box -8 -3 16 105
use FILL  FILL_562
timestamp 1677622389
transform 1 0 1472 0 1 4370
box -8 -3 16 105
use FILL  FILL_563
timestamp 1677622389
transform 1 0 1480 0 1 4370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1677622389
transform 1 0 1488 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1677622389
transform 1 0 1496 0 1 4370
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1677622389
transform 1 0 1512 0 1 4370
box -9 -3 26 105
use OAI22X1  OAI22X1_26
timestamp 1677622389
transform -1 0 1568 0 1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1677622389
transform 1 0 1568 0 1 4370
box -8 -3 104 105
use FILL  FILL_565
timestamp 1677622389
transform 1 0 1664 0 1 4370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1677622389
transform 1 0 1672 0 1 4370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1677622389
transform 1 0 1680 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1677622389
transform 1 0 1688 0 1 4370
box -8 -3 104 105
use FILL  FILL_576
timestamp 1677622389
transform 1 0 1784 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1677622389
transform -1 0 1808 0 1 4370
box -9 -3 26 105
use FILL  FILL_577
timestamp 1677622389
transform 1 0 1808 0 1 4370
box -8 -3 16 105
use FILL  FILL_578
timestamp 1677622389
transform 1 0 1816 0 1 4370
box -8 -3 16 105
use FILL  FILL_581
timestamp 1677622389
transform 1 0 1824 0 1 4370
box -8 -3 16 105
use FILL  FILL_583
timestamp 1677622389
transform 1 0 1832 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_28
timestamp 1677622389
transform 1 0 1840 0 1 4370
box -8 -3 46 105
use FILL  FILL_585
timestamp 1677622389
transform 1 0 1880 0 1 4370
box -8 -3 16 105
use FILL  FILL_587
timestamp 1677622389
transform 1 0 1888 0 1 4370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1677622389
transform 1 0 1896 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_28
timestamp 1677622389
transform 1 0 1904 0 1 4370
box -8 -3 46 105
use FILL  FILL_591
timestamp 1677622389
transform 1 0 1944 0 1 4370
box -8 -3 16 105
use FILL  FILL_592
timestamp 1677622389
transform 1 0 1952 0 1 4370
box -8 -3 16 105
use FILL  FILL_595
timestamp 1677622389
transform 1 0 1960 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_557
timestamp 1677622389
transform 1 0 2004 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_46
timestamp 1677622389
transform -1 0 2064 0 1 4370
box -8 -3 104 105
use FILL  FILL_596
timestamp 1677622389
transform 1 0 2064 0 1 4370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1677622389
transform 1 0 2072 0 1 4370
box -8 -3 16 105
use FILL  FILL_605
timestamp 1677622389
transform 1 0 2080 0 1 4370
box -8 -3 16 105
use FILL  FILL_606
timestamp 1677622389
transform 1 0 2088 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_31
timestamp 1677622389
transform 1 0 2096 0 1 4370
box -8 -3 46 105
use FILL  FILL_607
timestamp 1677622389
transform 1 0 2136 0 1 4370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1677622389
transform 1 0 2144 0 1 4370
box -8 -3 16 105
use FILL  FILL_615
timestamp 1677622389
transform 1 0 2152 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_55
timestamp 1677622389
transform 1 0 2160 0 1 4370
box -9 -3 26 105
use FILL  FILL_617
timestamp 1677622389
transform 1 0 2176 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1677622389
transform -1 0 2280 0 1 4370
box -8 -3 104 105
use AOI22X1  AOI22X1_32
timestamp 1677622389
transform 1 0 2280 0 1 4370
box -8 -3 46 105
use FILL  FILL_618
timestamp 1677622389
transform 1 0 2320 0 1 4370
box -8 -3 16 105
use FILL  FILL_619
timestamp 1677622389
transform 1 0 2328 0 1 4370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1677622389
transform 1 0 2336 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_56
timestamp 1677622389
transform 1 0 2344 0 1 4370
box -9 -3 26 105
use FILL  FILL_621
timestamp 1677622389
transform 1 0 2360 0 1 4370
box -8 -3 16 105
use FILL  FILL_629
timestamp 1677622389
transform 1 0 2368 0 1 4370
box -8 -3 16 105
use FILL  FILL_631
timestamp 1677622389
transform 1 0 2376 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1677622389
transform 1 0 2384 0 1 4370
box -8 -3 104 105
use FILL  FILL_633
timestamp 1677622389
transform 1 0 2480 0 1 4370
box -8 -3 16 105
use FILL  FILL_634
timestamp 1677622389
transform 1 0 2488 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_58
timestamp 1677622389
transform -1 0 2512 0 1 4370
box -9 -3 26 105
use AOI22X1  AOI22X1_34
timestamp 1677622389
transform 1 0 2512 0 1 4370
box -8 -3 46 105
use INVX2  INVX2_59
timestamp 1677622389
transform 1 0 2552 0 1 4370
box -9 -3 26 105
use FILL  FILL_635
timestamp 1677622389
transform 1 0 2568 0 1 4370
box -8 -3 16 105
use FILL  FILL_636
timestamp 1677622389
transform 1 0 2576 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_558
timestamp 1677622389
transform 1 0 2612 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1677622389
transform 1 0 2644 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_50
timestamp 1677622389
transform 1 0 2584 0 1 4370
box -8 -3 104 105
use FILL  FILL_637
timestamp 1677622389
transform 1 0 2680 0 1 4370
box -8 -3 16 105
use FILL  FILL_638
timestamp 1677622389
transform 1 0 2688 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_35
timestamp 1677622389
transform 1 0 2696 0 1 4370
box -8 -3 46 105
use INVX2  INVX2_60
timestamp 1677622389
transform 1 0 2736 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1677622389
transform 1 0 2752 0 1 4370
box -8 -3 104 105
use OAI21X1  OAI21X1_18
timestamp 1677622389
transform 1 0 2848 0 1 4370
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1677622389
transform 1 0 2880 0 1 4370
box -8 -3 34 105
use FILL  FILL_639
timestamp 1677622389
transform 1 0 2912 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_560
timestamp 1677622389
transform 1 0 2932 0 1 4375
box -3 -3 3 3
use NOR2X1  NOR2X1_7
timestamp 1677622389
transform 1 0 2920 0 1 4370
box -8 -3 32 105
use FILL  FILL_640
timestamp 1677622389
transform 1 0 2944 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1677622389
transform -1 0 2984 0 1 4370
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1677622389
transform -1 0 3016 0 1 4370
box -8 -3 34 105
use FILL  FILL_641
timestamp 1677622389
transform 1 0 3016 0 1 4370
box -8 -3 16 105
use FILL  FILL_642
timestamp 1677622389
transform 1 0 3024 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_30
timestamp 1677622389
transform 1 0 3032 0 1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1677622389
transform -1 0 3168 0 1 4370
box -8 -3 104 105
use FILL  FILL_643
timestamp 1677622389
transform 1 0 3168 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1677622389
transform 1 0 3176 0 1 4370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1677622389
transform 1 0 3272 0 1 4370
box -8 -3 104 105
use FILL  FILL_644
timestamp 1677622389
transform 1 0 3368 0 1 4370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1677622389
transform 1 0 3376 0 1 4370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1677622389
transform 1 0 3384 0 1 4370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1677622389
transform 1 0 3392 0 1 4370
box -8 -3 16 105
use FILL  FILL_702
timestamp 1677622389
transform 1 0 3400 0 1 4370
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1677622389
transform -1 0 3440 0 1 4370
box -8 -3 40 105
use FILL  FILL_703
timestamp 1677622389
transform 1 0 3440 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1677622389
transform -1 0 3544 0 1 4370
box -8 -3 104 105
use FILL  FILL_704
timestamp 1677622389
transform 1 0 3544 0 1 4370
box -8 -3 16 105
use FILL  FILL_705
timestamp 1677622389
transform 1 0 3552 0 1 4370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1677622389
transform 1 0 3560 0 1 4370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1677622389
transform 1 0 3568 0 1 4370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1677622389
transform 1 0 3576 0 1 4370
box -8 -3 16 105
use FILL  FILL_720
timestamp 1677622389
transform 1 0 3584 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1677622389
transform 1 0 3592 0 1 4370
box -8 -3 104 105
use FILL  FILL_722
timestamp 1677622389
transform 1 0 3688 0 1 4370
box -8 -3 16 105
use FILL  FILL_729
timestamp 1677622389
transform 1 0 3696 0 1 4370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1677622389
transform 1 0 3704 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1677622389
transform 1 0 3712 0 1 4370
box -8 -3 104 105
use FILL  FILL_732
timestamp 1677622389
transform 1 0 3808 0 1 4370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1677622389
transform 1 0 3816 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_561
timestamp 1677622389
transform 1 0 3844 0 1 4375
box -3 -3 3 3
use INVX2  INVX2_69
timestamp 1677622389
transform 1 0 3824 0 1 4370
box -9 -3 26 105
use FILL  FILL_734
timestamp 1677622389
transform 1 0 3840 0 1 4370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1677622389
transform 1 0 3848 0 1 4370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1677622389
transform 1 0 3856 0 1 4370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1677622389
transform 1 0 3864 0 1 4370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1677622389
transform 1 0 3872 0 1 4370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1677622389
transform 1 0 3880 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_562
timestamp 1677622389
transform 1 0 3924 0 1 4375
box -3 -3 3 3
use AOI22X1  AOI22X1_39
timestamp 1677622389
transform 1 0 3888 0 1 4370
box -8 -3 46 105
use FILL  FILL_751
timestamp 1677622389
transform 1 0 3928 0 1 4370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1677622389
transform 1 0 3936 0 1 4370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1677622389
transform 1 0 3944 0 1 4370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1677622389
transform 1 0 3952 0 1 4370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1677622389
transform 1 0 3960 0 1 4370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1677622389
transform 1 0 3968 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_563
timestamp 1677622389
transform 1 0 3996 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_37
timestamp 1677622389
transform 1 0 3976 0 1 4370
box -8 -3 46 105
use FILL  FILL_757
timestamp 1677622389
transform 1 0 4016 0 1 4370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1677622389
transform 1 0 4024 0 1 4370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1677622389
transform 1 0 4032 0 1 4370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1677622389
transform 1 0 4040 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1677622389
transform 1 0 4048 0 1 4370
box -8 -3 104 105
use FILL  FILL_765
timestamp 1677622389
transform 1 0 4144 0 1 4370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1677622389
transform 1 0 4152 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1677622389
transform 1 0 4160 0 1 4370
box -8 -3 104 105
use FILL  FILL_767
timestamp 1677622389
transform 1 0 4256 0 1 4370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1677622389
transform 1 0 4264 0 1 4370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1677622389
transform 1 0 4272 0 1 4370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1677622389
transform 1 0 4280 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1677622389
transform 1 0 4288 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_73
timestamp 1677622389
transform 1 0 4384 0 1 4370
box -9 -3 26 105
use FILL  FILL_778
timestamp 1677622389
transform 1 0 4400 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_40
timestamp 1677622389
transform -1 0 4448 0 1 4370
box -8 -3 46 105
use FILL  FILL_779
timestamp 1677622389
transform 1 0 4448 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_564
timestamp 1677622389
transform 1 0 4468 0 1 4375
box -3 -3 3 3
use FILL  FILL_780
timestamp 1677622389
transform 1 0 4456 0 1 4370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1677622389
transform 1 0 4464 0 1 4370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1677622389
transform 1 0 4472 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_39
timestamp 1677622389
transform 1 0 4480 0 1 4370
box -8 -3 46 105
use FILL  FILL_783
timestamp 1677622389
transform 1 0 4520 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1677622389
transform 1 0 4528 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_74
timestamp 1677622389
transform 1 0 4624 0 1 4370
box -9 -3 26 105
use OAI22X1  OAI22X1_42
timestamp 1677622389
transform 1 0 4640 0 1 4370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1677622389
transform 1 0 4680 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_75
timestamp 1677622389
transform 1 0 4776 0 1 4370
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_7
timestamp 1677622389
transform 1 0 4819 0 1 4370
box -10 -3 10 3
use M2_M1  M2_M1_790
timestamp 1677622389
transform 1 0 164 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_581
timestamp 1677622389
transform 1 0 220 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_678
timestamp 1677622389
transform 1 0 220 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1677622389
transform 1 0 212 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1677622389
transform 1 0 228 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_676
timestamp 1677622389
transform 1 0 228 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_679
timestamp 1677622389
transform 1 0 244 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_623
timestamp 1677622389
transform 1 0 252 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1677622389
transform 1 0 244 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1677622389
transform 1 0 252 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_602
timestamp 1677622389
transform 1 0 260 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_680
timestamp 1677622389
transform 1 0 260 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1677622389
transform 1 0 284 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1677622389
transform 1 0 300 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_794
timestamp 1677622389
transform 1 0 308 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_625
timestamp 1677622389
transform 1 0 324 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_795
timestamp 1677622389
transform 1 0 324 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_603
timestamp 1677622389
transform 1 0 372 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1677622389
transform 1 0 348 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1677622389
transform 1 0 356 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1677622389
transform 1 0 372 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_658
timestamp 1677622389
transform 1 0 356 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_796
timestamp 1677622389
transform 1 0 364 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1677622389
transform 1 0 380 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1677622389
transform 1 0 412 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1677622389
transform 1 0 460 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1677622389
transform 1 0 492 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1677622389
transform 1 0 500 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_678
timestamp 1677622389
transform 1 0 460 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1677622389
transform 1 0 500 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1677622389
transform 1 0 492 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_801
timestamp 1677622389
transform 1 0 516 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1677622389
transform 1 0 532 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_685
timestamp 1677622389
transform 1 0 548 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1677622389
transform 1 0 556 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1677622389
transform 1 0 572 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_659
timestamp 1677622389
transform 1 0 556 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_802
timestamp 1677622389
transform 1 0 564 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_701
timestamp 1677622389
transform 1 0 556 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1677622389
transform 1 0 612 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1677622389
transform 1 0 612 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1677622389
transform 1 0 644 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1677622389
transform 1 0 652 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1677622389
transform 1 0 620 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1677622389
transform 1 0 636 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1677622389
transform 1 0 652 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_702
timestamp 1677622389
transform 1 0 644 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1677622389
transform 1 0 620 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1677622389
transform 1 0 700 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_680
timestamp 1677622389
transform 1 0 700 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_691
timestamp 1677622389
transform 1 0 716 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_626
timestamp 1677622389
transform 1 0 748 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1677622389
transform 1 0 796 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_692
timestamp 1677622389
transform 1 0 812 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1677622389
transform 1 0 740 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1677622389
transform 1 0 796 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1677622389
transform 1 0 804 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_681
timestamp 1677622389
transform 1 0 740 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1677622389
transform 1 0 756 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1677622389
transform 1 0 796 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1677622389
transform 1 0 812 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_693
timestamp 1677622389
transform 1 0 836 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1677622389
transform 1 0 852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1677622389
transform 1 0 844 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_628
timestamp 1677622389
transform 1 0 860 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1677622389
transform 1 0 852 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_811
timestamp 1677622389
transform 1 0 868 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1677622389
transform 1 0 884 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1677622389
transform 1 0 884 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_695
timestamp 1677622389
transform 1 0 908 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1677622389
transform 1 0 916 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1677622389
transform 1 0 932 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_629
timestamp 1677622389
transform 1 0 940 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_813
timestamp 1677622389
transform 1 0 924 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1677622389
transform 1 0 940 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1677622389
transform 1 0 916 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1677622389
transform 1 0 1020 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_698
timestamp 1677622389
transform 1 0 1012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1677622389
transform 1 0 996 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1677622389
transform 1 0 996 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1677622389
transform 1 0 1020 0 1 4345
box -2 -2 2 2
use M3_M2  M3_M2_630
timestamp 1677622389
transform 1 0 1036 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1677622389
transform 1 0 1052 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_909
timestamp 1677622389
transform 1 0 1052 0 1 4315
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1677622389
transform 1 0 1084 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1677622389
transform 1 0 1076 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_700
timestamp 1677622389
transform 1 0 1108 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1677622389
transform 1 0 1124 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1677622389
transform 1 0 1156 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1677622389
transform 1 0 1132 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1677622389
transform 1 0 1148 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_701
timestamp 1677622389
transform 1 0 1156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1677622389
transform 1 0 1124 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1677622389
transform 1 0 1132 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1677622389
transform 1 0 1132 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1677622389
transform 1 0 1180 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1677622389
transform 1 0 1180 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_910
timestamp 1677622389
transform 1 0 1196 0 1 4315
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1677622389
transform 1 0 1260 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1677622389
transform 1 0 1252 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1677622389
transform 1 0 1260 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1677622389
transform 1 0 1308 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1677622389
transform 1 0 1276 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_703
timestamp 1677622389
transform 1 0 1276 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_633
timestamp 1677622389
transform 1 0 1300 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_819
timestamp 1677622389
transform 1 0 1324 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_688
timestamp 1677622389
transform 1 0 1324 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1677622389
transform 1 0 1380 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1677622389
transform 1 0 1364 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_634
timestamp 1677622389
transform 1 0 1372 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_820
timestamp 1677622389
transform 1 0 1364 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1677622389
transform 1 0 1372 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_689
timestamp 1677622389
transform 1 0 1412 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1677622389
transform 1 0 1444 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_705
timestamp 1677622389
transform 1 0 1460 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1677622389
transform 1 0 1476 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1677622389
transform 1 0 1492 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1677622389
transform 1 0 1468 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1677622389
transform 1 0 1484 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1677622389
transform 1 0 1508 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1677622389
transform 1 0 1500 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1677622389
transform 1 0 1492 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1677622389
transform 1 0 1580 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1677622389
transform 1 0 1628 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_708
timestamp 1677622389
transform 1 0 1540 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_635
timestamp 1677622389
transform 1 0 1548 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1677622389
transform 1 0 1628 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1677622389
transform 1 0 1548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1677622389
transform 1 0 1580 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1677622389
transform 1 0 1580 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_827
timestamp 1677622389
transform 1 0 1644 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_613
timestamp 1677622389
transform 1 0 1668 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_710
timestamp 1677622389
transform 1 0 1660 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1677622389
transform 1 0 1676 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_711
timestamp 1677622389
transform 1 0 1684 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1677622389
transform 1 0 1676 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_692
timestamp 1677622389
transform 1 0 1676 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_712
timestamp 1677622389
transform 1 0 1716 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_637
timestamp 1677622389
transform 1 0 1764 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1677622389
transform 1 0 1804 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_829
timestamp 1677622389
transform 1 0 1764 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1677622389
transform 1 0 1796 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1677622389
transform 1 0 1804 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1677622389
transform 1 0 1812 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_725
timestamp 1677622389
transform 1 0 1708 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1677622389
transform 1 0 1796 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1677622389
transform 1 0 1812 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_713
timestamp 1677622389
transform 1 0 1844 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1677622389
transform 1 0 1852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1677622389
transform 1 0 1868 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1677622389
transform 1 0 1860 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_708
timestamp 1677622389
transform 1 0 1868 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1677622389
transform 1 0 1884 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1677622389
transform 1 0 1932 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1677622389
transform 1 0 1916 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1677622389
transform 1 0 1940 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1677622389
transform 1 0 1956 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_717
timestamp 1677622389
transform 1 0 1956 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_583
timestamp 1677622389
transform 1 0 1988 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_718
timestamp 1677622389
transform 1 0 1996 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1677622389
transform 1 0 1988 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_661
timestamp 1677622389
transform 1 0 1996 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_911
timestamp 1677622389
transform 1 0 1996 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_709
timestamp 1677622389
transform 1 0 1996 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1677622389
transform 1 0 2020 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1677622389
transform 1 0 2012 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_719
timestamp 1677622389
transform 1 0 2012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1677622389
transform 1 0 2028 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_639
timestamp 1677622389
transform 1 0 2036 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1677622389
transform 1 0 2012 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1677622389
transform 1 0 2020 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1677622389
transform 1 0 2036 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1677622389
transform 1 0 2044 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_840
timestamp 1677622389
transform 1 0 2052 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1677622389
transform 1 0 2036 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1677622389
transform 1 0 2052 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_721
timestamp 1677622389
transform 1 0 2076 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1677622389
transform 1 0 2092 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1677622389
transform 1 0 2100 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1677622389
transform 1 0 2100 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_841
timestamp 1677622389
transform 1 0 2148 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_711
timestamp 1677622389
transform 1 0 2140 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_724
timestamp 1677622389
transform 1 0 2172 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1677622389
transform 1 0 2220 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1677622389
transform 1 0 2244 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_843
timestamp 1677622389
transform 1 0 2252 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1677622389
transform 1 0 2260 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_712
timestamp 1677622389
transform 1 0 2220 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1677622389
transform 1 0 2260 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_725
timestamp 1677622389
transform 1 0 2316 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1677622389
transform 1 0 2324 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1677622389
transform 1 0 2340 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1677622389
transform 1 0 2308 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1677622389
transform 1 0 2324 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1677622389
transform 1 0 2332 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1677622389
transform 1 0 2380 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1677622389
transform 1 0 2484 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1677622389
transform 1 0 2388 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1677622389
transform 1 0 2396 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1677622389
transform 1 0 2404 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1677622389
transform 1 0 2412 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_850
timestamp 1677622389
transform 1 0 2436 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_714
timestamp 1677622389
transform 1 0 2396 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1677622389
transform 1 0 2436 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1677622389
transform 1 0 2524 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_730
timestamp 1677622389
transform 1 0 2532 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_640
timestamp 1677622389
transform 1 0 2540 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1677622389
transform 1 0 2532 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1677622389
transform 1 0 2556 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1677622389
transform 1 0 2556 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_851
timestamp 1677622389
transform 1 0 2540 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1677622389
transform 1 0 2548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1677622389
transform 1 0 2556 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1677622389
transform 1 0 2604 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1677622389
transform 1 0 2596 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1677622389
transform 1 0 2604 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1677622389
transform 1 0 2580 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_853
timestamp 1677622389
transform 1 0 2588 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_716
timestamp 1677622389
transform 1 0 2596 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_854
timestamp 1677622389
transform 1 0 2612 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1677622389
transform 1 0 2628 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1677622389
transform 1 0 2628 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1677622389
transform 1 0 2676 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_735
timestamp 1677622389
transform 1 0 2660 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1677622389
transform 1 0 2668 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1677622389
transform 1 0 2652 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_670
timestamp 1677622389
transform 1 0 2660 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1677622389
transform 1 0 2684 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_856
timestamp 1677622389
transform 1 0 2676 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_641
timestamp 1677622389
transform 1 0 2708 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_857
timestamp 1677622389
transform 1 0 2708 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_572
timestamp 1677622389
transform 1 0 2740 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1677622389
transform 1 0 2724 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1677622389
transform 1 0 2764 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1677622389
transform 1 0 2724 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_642
timestamp 1677622389
transform 1 0 2748 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_858
timestamp 1677622389
transform 1 0 2748 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_671
timestamp 1677622389
transform 1 0 2796 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_674
timestamp 1677622389
transform 1 0 2812 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1677622389
transform 1 0 2804 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1677622389
transform 1 0 2836 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1677622389
transform 1 0 2836 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1677622389
transform 1 0 2852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1677622389
transform 1 0 2844 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1677622389
transform 1 0 2852 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1677622389
transform 1 0 2844 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_861
timestamp 1677622389
transform 1 0 2868 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1677622389
transform 1 0 2868 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_675
timestamp 1677622389
transform 1 0 2900 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1677622389
transform 1 0 2908 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1677622389
transform 1 0 2908 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_912
timestamp 1677622389
transform 1 0 2900 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1677622389
transform 1 0 2900 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1677622389
transform 1 0 2892 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_676
timestamp 1677622389
transform 1 0 2932 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1677622389
transform 1 0 2924 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1677622389
transform 1 0 2932 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1677622389
transform 1 0 2956 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_673
timestamp 1677622389
transform 1 0 2964 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1677622389
transform 1 0 2980 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1677622389
transform 1 0 2972 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1677622389
transform 1 0 2996 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1677622389
transform 1 0 2988 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1677622389
transform 1 0 2980 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1677622389
transform 1 0 3020 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_864
timestamp 1677622389
transform 1 0 3020 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_694
timestamp 1677622389
transform 1 0 3036 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1677622389
transform 1 0 3044 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1677622389
transform 1 0 3036 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1677622389
transform 1 0 3076 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1677622389
transform 1 0 3116 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_743
timestamp 1677622389
transform 1 0 3068 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1677622389
transform 1 0 3076 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1677622389
transform 1 0 3092 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1677622389
transform 1 0 3108 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1677622389
transform 1 0 3116 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1677622389
transform 1 0 3084 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1677622389
transform 1 0 3100 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_721
timestamp 1677622389
transform 1 0 3100 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1677622389
transform 1 0 3156 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1677622389
transform 1 0 3204 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1677622389
transform 1 0 3180 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_748
timestamp 1677622389
transform 1 0 3188 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1677622389
transform 1 0 3204 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_645
timestamp 1677622389
transform 1 0 3212 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1677622389
transform 1 0 3180 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_675
timestamp 1677622389
transform 1 0 3188 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_868
timestamp 1677622389
transform 1 0 3196 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1677622389
transform 1 0 3212 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1677622389
transform 1 0 3196 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_870
timestamp 1677622389
transform 1 0 3236 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1677622389
transform 1 0 3260 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1677622389
transform 1 0 3276 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1677622389
transform 1 0 3356 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1677622389
transform 1 0 3420 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1677622389
transform 1 0 3412 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_646
timestamp 1677622389
transform 1 0 3428 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_754
timestamp 1677622389
transform 1 0 3436 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1677622389
transform 1 0 3452 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1677622389
transform 1 0 3460 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1677622389
transform 1 0 3428 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1677622389
transform 1 0 3500 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_873
timestamp 1677622389
transform 1 0 3492 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_736
timestamp 1677622389
transform 1 0 3492 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1677622389
transform 1 0 3532 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1677622389
transform 1 0 3524 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_648
timestamp 1677622389
transform 1 0 3540 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_758
timestamp 1677622389
transform 1 0 3548 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1677622389
transform 1 0 3540 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1677622389
transform 1 0 3564 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1677622389
transform 1 0 3572 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_695
timestamp 1677622389
transform 1 0 3540 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1677622389
transform 1 0 3588 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1677622389
transform 1 0 3580 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1677622389
transform 1 0 3612 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1677622389
transform 1 0 3604 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1677622389
transform 1 0 3620 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1677622389
transform 1 0 3636 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1677622389
transform 1 0 3628 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1677622389
transform 1 0 3644 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1677622389
transform 1 0 3684 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1677622389
transform 1 0 3708 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_738
timestamp 1677622389
transform 1 0 3708 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1677622389
transform 1 0 3748 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1677622389
transform 1 0 3732 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_763
timestamp 1677622389
transform 1 0 3740 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1677622389
transform 1 0 3748 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1677622389
transform 1 0 3732 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1677622389
transform 1 0 3804 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_651
timestamp 1677622389
transform 1 0 3812 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_766
timestamp 1677622389
transform 1 0 3820 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1677622389
transform 1 0 3788 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1677622389
transform 1 0 3796 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1677622389
transform 1 0 3812 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_652
timestamp 1677622389
transform 1 0 3836 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1677622389
transform 1 0 3836 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1677622389
transform 1 0 3860 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_767
timestamp 1677622389
transform 1 0 3860 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_574
timestamp 1677622389
transform 1 0 3892 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1677622389
transform 1 0 3900 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1677622389
transform 1 0 3948 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_768
timestamp 1677622389
transform 1 0 3996 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1677622389
transform 1 0 4012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1677622389
transform 1 0 3900 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1677622389
transform 1 0 3916 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1677622389
transform 1 0 3948 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1677622389
transform 1 0 3884 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_740
timestamp 1677622389
transform 1 0 3876 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_915
timestamp 1677622389
transform 1 0 3908 0 1 4315
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1677622389
transform 1 0 3892 0 1 4305
box -2 -2 2 2
use M3_M2  M3_M2_596
timestamp 1677622389
transform 1 0 4028 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_770
timestamp 1677622389
transform 1 0 4028 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1677622389
transform 1 0 4020 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1677622389
transform 1 0 4028 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_741
timestamp 1677622389
transform 1 0 3948 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1677622389
transform 1 0 3980 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1677622389
transform 1 0 4012 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1677622389
transform 1 0 4028 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1677622389
transform 1 0 4060 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1677622389
transform 1 0 4084 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_771
timestamp 1677622389
transform 1 0 4084 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1677622389
transform 1 0 4108 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_732
timestamp 1677622389
transform 1 0 4076 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1677622389
transform 1 0 4156 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1677622389
transform 1 0 4180 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1677622389
transform 1 0 4180 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1677622389
transform 1 0 4172 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1677622389
transform 1 0 4180 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1677622389
transform 1 0 4196 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1677622389
transform 1 0 4188 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1677622389
transform 1 0 4180 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1677622389
transform 1 0 4228 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_773
timestamp 1677622389
transform 1 0 4212 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1677622389
transform 1 0 4220 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1677622389
transform 1 0 4228 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1677622389
transform 1 0 4220 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1677622389
transform 1 0 4236 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1677622389
transform 1 0 4252 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1677622389
transform 1 0 4252 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_747
timestamp 1677622389
transform 1 0 4252 0 1 4285
box -3 -3 3 3
use M2_M1  M2_M1_776
timestamp 1677622389
transform 1 0 4268 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_577
timestamp 1677622389
transform 1 0 4316 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1677622389
transform 1 0 4348 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1677622389
transform 1 0 4364 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1677622389
transform 1 0 4308 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_777
timestamp 1677622389
transform 1 0 4292 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_655
timestamp 1677622389
transform 1 0 4300 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1677622389
transform 1 0 4316 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1677622389
transform 1 0 4348 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_778
timestamp 1677622389
transform 1 0 4308 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1677622389
transform 1 0 4316 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1677622389
transform 1 0 4300 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1677622389
transform 1 0 4332 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_780
timestamp 1677622389
transform 1 0 4340 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1677622389
transform 1 0 4324 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1677622389
transform 1 0 4348 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1677622389
transform 1 0 4364 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1677622389
transform 1 0 4364 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_619
timestamp 1677622389
transform 1 0 4380 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_782
timestamp 1677622389
transform 1 0 4380 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1677622389
transform 1 0 4388 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_696
timestamp 1677622389
transform 1 0 4364 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1677622389
transform 1 0 4356 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1677622389
transform 1 0 4420 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_783
timestamp 1677622389
transform 1 0 4420 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_697
timestamp 1677622389
transform 1 0 4412 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_901
timestamp 1677622389
transform 1 0 4428 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_620
timestamp 1677622389
transform 1 0 4452 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_784
timestamp 1677622389
transform 1 0 4444 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1677622389
transform 1 0 4452 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1677622389
transform 1 0 4460 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1677622389
transform 1 0 4476 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_698
timestamp 1677622389
transform 1 0 4476 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1677622389
transform 1 0 4516 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_786
timestamp 1677622389
transform 1 0 4508 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_699
timestamp 1677622389
transform 1 0 4532 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1677622389
transform 1 0 4572 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1677622389
transform 1 0 4596 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1677622389
transform 1 0 4652 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_621
timestamp 1677622389
transform 1 0 4668 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_788
timestamp 1677622389
transform 1 0 4684 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_601
timestamp 1677622389
transform 1 0 4788 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1677622389
transform 1 0 4780 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_789
timestamp 1677622389
transform 1 0 4772 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1677622389
transform 1 0 4708 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1677622389
transform 1 0 4764 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1677622389
transform 1 0 4780 0 1 4325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_8
timestamp 1677622389
transform 1 0 24 0 1 4270
box -10 -3 10 3
use FILL  FILL_424
timestamp 1677622389
transform 1 0 72 0 -1 4370
box -8 -3 16 105
use FILL  FILL_426
timestamp 1677622389
transform 1 0 80 0 -1 4370
box -8 -3 16 105
use FILL  FILL_427
timestamp 1677622389
transform 1 0 88 0 -1 4370
box -8 -3 16 105
use FILL  FILL_428
timestamp 1677622389
transform 1 0 96 0 -1 4370
box -8 -3 16 105
use FILL  FILL_429
timestamp 1677622389
transform 1 0 104 0 -1 4370
box -8 -3 16 105
use FILL  FILL_430
timestamp 1677622389
transform 1 0 112 0 -1 4370
box -8 -3 16 105
use FILL  FILL_431
timestamp 1677622389
transform 1 0 120 0 -1 4370
box -8 -3 16 105
use FILL  FILL_432
timestamp 1677622389
transform 1 0 128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_433
timestamp 1677622389
transform 1 0 136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_434
timestamp 1677622389
transform 1 0 144 0 -1 4370
box -8 -3 16 105
use FILL  FILL_435
timestamp 1677622389
transform 1 0 152 0 -1 4370
box -8 -3 16 105
use FILL  FILL_436
timestamp 1677622389
transform 1 0 160 0 -1 4370
box -8 -3 16 105
use FILL  FILL_437
timestamp 1677622389
transform 1 0 168 0 -1 4370
box -8 -3 16 105
use FILL  FILL_438
timestamp 1677622389
transform 1 0 176 0 -1 4370
box -8 -3 16 105
use FILL  FILL_440
timestamp 1677622389
transform 1 0 184 0 -1 4370
box -8 -3 16 105
use FILL  FILL_442
timestamp 1677622389
transform 1 0 192 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_22
timestamp 1677622389
transform 1 0 200 0 -1 4370
box -8 -3 46 105
use FILL  FILL_444
timestamp 1677622389
transform 1 0 240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_446
timestamp 1677622389
transform 1 0 248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_448
timestamp 1677622389
transform 1 0 256 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_37
timestamp 1677622389
transform 1 0 264 0 -1 4370
box -9 -3 26 105
use FILL  FILL_453
timestamp 1677622389
transform 1 0 280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_454
timestamp 1677622389
transform 1 0 288 0 -1 4370
box -8 -3 16 105
use FILL  FILL_455
timestamp 1677622389
transform 1 0 296 0 -1 4370
box -8 -3 16 105
use FILL  FILL_456
timestamp 1677622389
transform 1 0 304 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_38
timestamp 1677622389
transform -1 0 328 0 -1 4370
box -9 -3 26 105
use FILL  FILL_457
timestamp 1677622389
transform 1 0 328 0 -1 4370
box -8 -3 16 105
use FILL  FILL_458
timestamp 1677622389
transform 1 0 336 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_21
timestamp 1677622389
transform -1 0 384 0 -1 4370
box -8 -3 46 105
use FILL  FILL_459
timestamp 1677622389
transform 1 0 384 0 -1 4370
box -8 -3 16 105
use FILL  FILL_462
timestamp 1677622389
transform 1 0 392 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1677622389
transform 1 0 400 0 -1 4370
box -8 -3 104 105
use FILL  FILL_463
timestamp 1677622389
transform 1 0 496 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_40
timestamp 1677622389
transform -1 0 520 0 -1 4370
box -9 -3 26 105
use FILL  FILL_465
timestamp 1677622389
transform 1 0 520 0 -1 4370
box -8 -3 16 105
use FILL  FILL_467
timestamp 1677622389
transform 1 0 528 0 -1 4370
box -8 -3 16 105
use FILL  FILL_470
timestamp 1677622389
transform 1 0 536 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_23
timestamp 1677622389
transform -1 0 584 0 -1 4370
box -8 -3 46 105
use FILL  FILL_471
timestamp 1677622389
transform 1 0 584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_473
timestamp 1677622389
transform 1 0 592 0 -1 4370
box -8 -3 16 105
use FILL  FILL_475
timestamp 1677622389
transform 1 0 600 0 -1 4370
box -8 -3 16 105
use FILL  FILL_477
timestamp 1677622389
transform 1 0 608 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_24
timestamp 1677622389
transform 1 0 616 0 -1 4370
box -8 -3 46 105
use INVX2  INVX2_41
timestamp 1677622389
transform 1 0 656 0 -1 4370
box -9 -3 26 105
use FILL  FILL_481
timestamp 1677622389
transform 1 0 672 0 -1 4370
box -8 -3 16 105
use FILL  FILL_486
timestamp 1677622389
transform 1 0 680 0 -1 4370
box -8 -3 16 105
use FILL  FILL_487
timestamp 1677622389
transform 1 0 688 0 -1 4370
box -8 -3 16 105
use FILL  FILL_488
timestamp 1677622389
transform 1 0 696 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_748
timestamp 1677622389
transform 1 0 772 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1677622389
transform 1 0 804 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_38
timestamp 1677622389
transform 1 0 704 0 -1 4370
box -8 -3 104 105
use FILL  FILL_489
timestamp 1677622389
transform 1 0 800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_491
timestamp 1677622389
transform 1 0 808 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_750
timestamp 1677622389
transform 1 0 844 0 1 4275
box -3 -3 3 3
use OAI22X1  OAI22X1_25
timestamp 1677622389
transform 1 0 816 0 -1 4370
box -8 -3 46 105
use FILL  FILL_497
timestamp 1677622389
transform 1 0 856 0 -1 4370
box -8 -3 16 105
use FILL  FILL_498
timestamp 1677622389
transform 1 0 864 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1677622389
transform -1 0 888 0 -1 4370
box -9 -3 26 105
use FILL  FILL_499
timestamp 1677622389
transform 1 0 888 0 -1 4370
box -8 -3 16 105
use FILL  FILL_500
timestamp 1677622389
transform 1 0 896 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_26
timestamp 1677622389
transform 1 0 904 0 -1 4370
box -8 -3 46 105
use FILL  FILL_501
timestamp 1677622389
transform 1 0 944 0 -1 4370
box -8 -3 16 105
use FILL  FILL_503
timestamp 1677622389
transform 1 0 952 0 -1 4370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1677622389
transform 1 0 960 0 -1 4370
box -8 -3 16 105
use FILL  FILL_505
timestamp 1677622389
transform 1 0 968 0 -1 4370
box -8 -3 16 105
use FILL  FILL_506
timestamp 1677622389
transform 1 0 976 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_12
timestamp 1677622389
transform 1 0 984 0 -1 4370
box -8 -3 34 105
use FILL  FILL_510
timestamp 1677622389
transform 1 0 1016 0 -1 4370
box -8 -3 16 105
use FILL  FILL_511
timestamp 1677622389
transform 1 0 1024 0 -1 4370
box -8 -3 16 105
use FILL  FILL_513
timestamp 1677622389
transform 1 0 1032 0 -1 4370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1677622389
transform 1 0 1040 0 -1 4370
box -8 -3 16 105
use FILL  FILL_519
timestamp 1677622389
transform 1 0 1048 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1677622389
transform 1 0 1056 0 -1 4370
box -8 -3 32 105
use FILL  FILL_520
timestamp 1677622389
transform 1 0 1080 0 -1 4370
box -8 -3 16 105
use FILL  FILL_521
timestamp 1677622389
transform 1 0 1088 0 -1 4370
box -8 -3 16 105
use FILL  FILL_522
timestamp 1677622389
transform 1 0 1096 0 -1 4370
box -8 -3 16 105
use FILL  FILL_523
timestamp 1677622389
transform 1 0 1104 0 -1 4370
box -8 -3 16 105
use FILL  FILL_524
timestamp 1677622389
transform 1 0 1112 0 -1 4370
box -8 -3 16 105
use FILL  FILL_525
timestamp 1677622389
transform 1 0 1120 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_16
timestamp 1677622389
transform 1 0 1128 0 -1 4370
box -8 -3 34 105
use FILL  FILL_541
timestamp 1677622389
transform 1 0 1160 0 -1 4370
box -8 -3 16 105
use FILL  FILL_542
timestamp 1677622389
transform 1 0 1168 0 -1 4370
box -8 -3 16 105
use FILL  FILL_543
timestamp 1677622389
transform 1 0 1176 0 -1 4370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1677622389
transform 1 0 1184 0 -1 4370
box -8 -3 16 105
use FILL  FILL_545
timestamp 1677622389
transform 1 0 1192 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1677622389
transform -1 0 1232 0 -1 4370
box -8 -3 34 105
use FILL  FILL_546
timestamp 1677622389
transform 1 0 1232 0 -1 4370
box -8 -3 16 105
use FILL  FILL_547
timestamp 1677622389
transform 1 0 1240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_548
timestamp 1677622389
transform 1 0 1248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_549
timestamp 1677622389
transform 1 0 1256 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1677622389
transform 1 0 1264 0 -1 4370
box -8 -3 104 105
use FILL  FILL_550
timestamp 1677622389
transform 1 0 1360 0 -1 4370
box -8 -3 16 105
use FILL  FILL_551
timestamp 1677622389
transform 1 0 1368 0 -1 4370
box -8 -3 16 105
use FILL  FILL_552
timestamp 1677622389
transform 1 0 1376 0 -1 4370
box -8 -3 16 105
use FILL  FILL_553
timestamp 1677622389
transform 1 0 1384 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_45
timestamp 1677622389
transform 1 0 1392 0 -1 4370
box -9 -3 26 105
use FILL  FILL_554
timestamp 1677622389
transform 1 0 1408 0 -1 4370
box -8 -3 16 105
use FILL  FILL_555
timestamp 1677622389
transform 1 0 1416 0 -1 4370
box -8 -3 16 105
use FILL  FILL_556
timestamp 1677622389
transform 1 0 1424 0 -1 4370
box -8 -3 16 105
use FILL  FILL_557
timestamp 1677622389
transform 1 0 1432 0 -1 4370
box -8 -3 16 105
use FILL  FILL_558
timestamp 1677622389
transform 1 0 1440 0 -1 4370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1677622389
transform 1 0 1448 0 -1 4370
box -8 -3 16 105
use FILL  FILL_560
timestamp 1677622389
transform 1 0 1456 0 -1 4370
box -8 -3 16 105
use FILL  FILL_567
timestamp 1677622389
transform 1 0 1464 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_27
timestamp 1677622389
transform -1 0 1512 0 -1 4370
box -8 -3 46 105
use FILL  FILL_568
timestamp 1677622389
transform 1 0 1512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1677622389
transform 1 0 1520 0 -1 4370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1677622389
transform 1 0 1528 0 -1 4370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1677622389
transform 1 0 1536 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_751
timestamp 1677622389
transform 1 0 1604 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_43
timestamp 1677622389
transform -1 0 1640 0 -1 4370
box -8 -3 104 105
use FILL  FILL_572
timestamp 1677622389
transform 1 0 1640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_573
timestamp 1677622389
transform 1 0 1648 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_48
timestamp 1677622389
transform 1 0 1656 0 -1 4370
box -9 -3 26 105
use FILL  FILL_574
timestamp 1677622389
transform 1 0 1672 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_50
timestamp 1677622389
transform 1 0 1680 0 -1 4370
box -9 -3 26 105
use FILL  FILL_579
timestamp 1677622389
transform 1 0 1696 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1677622389
transform 1 0 1704 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_51
timestamp 1677622389
transform -1 0 1816 0 -1 4370
box -9 -3 26 105
use FILL  FILL_580
timestamp 1677622389
transform 1 0 1816 0 -1 4370
box -8 -3 16 105
use FILL  FILL_582
timestamp 1677622389
transform 1 0 1824 0 -1 4370
box -8 -3 16 105
use FILL  FILL_584
timestamp 1677622389
transform 1 0 1832 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_29
timestamp 1677622389
transform 1 0 1840 0 -1 4370
box -8 -3 46 105
use FILL  FILL_586
timestamp 1677622389
transform 1 0 1880 0 -1 4370
box -8 -3 16 105
use FILL  FILL_588
timestamp 1677622389
transform 1 0 1888 0 -1 4370
box -8 -3 16 105
use FILL  FILL_590
timestamp 1677622389
transform 1 0 1896 0 -1 4370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1677622389
transform 1 0 1904 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_29
timestamp 1677622389
transform 1 0 1912 0 -1 4370
box -8 -3 46 105
use FILL  FILL_594
timestamp 1677622389
transform 1 0 1952 0 -1 4370
box -8 -3 16 105
use FILL  FILL_597
timestamp 1677622389
transform 1 0 1960 0 -1 4370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1677622389
transform 1 0 1968 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_752
timestamp 1677622389
transform 1 0 1988 0 1 4275
box -3 -3 3 3
use INVX2  INVX2_52
timestamp 1677622389
transform -1 0 1992 0 -1 4370
box -9 -3 26 105
use FILL  FILL_599
timestamp 1677622389
transform 1 0 1992 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_30
timestamp 1677622389
transform -1 0 2040 0 -1 4370
box -8 -3 46 105
use FILL  FILL_600
timestamp 1677622389
transform 1 0 2040 0 -1 4370
box -8 -3 16 105
use FILL  FILL_601
timestamp 1677622389
transform 1 0 2048 0 -1 4370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1677622389
transform 1 0 2056 0 -1 4370
box -8 -3 16 105
use FILL  FILL_603
timestamp 1677622389
transform 1 0 2064 0 -1 4370
box -8 -3 16 105
use FILL  FILL_608
timestamp 1677622389
transform 1 0 2072 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1677622389
transform -1 0 2096 0 -1 4370
box -9 -3 26 105
use FILL  FILL_609
timestamp 1677622389
transform 1 0 2096 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1677622389
transform 1 0 2104 0 -1 4370
box -9 -3 26 105
use FILL  FILL_610
timestamp 1677622389
transform 1 0 2120 0 -1 4370
box -8 -3 16 105
use FILL  FILL_611
timestamp 1677622389
transform 1 0 2128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_612
timestamp 1677622389
transform 1 0 2136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_614
timestamp 1677622389
transform 1 0 2144 0 -1 4370
box -8 -3 16 105
use FILL  FILL_616
timestamp 1677622389
transform 1 0 2152 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1677622389
transform 1 0 2160 0 -1 4370
box -8 -3 104 105
use FILL  FILL_622
timestamp 1677622389
transform 1 0 2256 0 -1 4370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1677622389
transform 1 0 2264 0 -1 4370
box -8 -3 16 105
use FILL  FILL_624
timestamp 1677622389
transform 1 0 2272 0 -1 4370
box -8 -3 16 105
use FILL  FILL_625
timestamp 1677622389
transform 1 0 2280 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1677622389
transform -1 0 2304 0 -1 4370
box -9 -3 26 105
use FILL  FILL_626
timestamp 1677622389
transform 1 0 2304 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_33
timestamp 1677622389
transform -1 0 2352 0 -1 4370
box -8 -3 46 105
use FILL  FILL_627
timestamp 1677622389
transform 1 0 2352 0 -1 4370
box -8 -3 16 105
use FILL  FILL_628
timestamp 1677622389
transform 1 0 2360 0 -1 4370
box -8 -3 16 105
use FILL  FILL_630
timestamp 1677622389
transform 1 0 2368 0 -1 4370
box -8 -3 16 105
use FILL  FILL_632
timestamp 1677622389
transform 1 0 2376 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1677622389
transform 1 0 2384 0 -1 4370
box -9 -3 26 105
use M3_M2  M3_M2_753
timestamp 1677622389
transform 1 0 2452 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_55
timestamp 1677622389
transform -1 0 2496 0 -1 4370
box -8 -3 104 105
use FILL  FILL_645
timestamp 1677622389
transform 1 0 2496 0 -1 4370
box -8 -3 16 105
use FILL  FILL_646
timestamp 1677622389
transform 1 0 2504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_647
timestamp 1677622389
transform 1 0 2512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_648
timestamp 1677622389
transform 1 0 2520 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_62
timestamp 1677622389
transform 1 0 2528 0 -1 4370
box -9 -3 26 105
use FILL  FILL_649
timestamp 1677622389
transform 1 0 2544 0 -1 4370
box -8 -3 16 105
use FILL  FILL_650
timestamp 1677622389
transform 1 0 2552 0 -1 4370
box -8 -3 16 105
use FILL  FILL_651
timestamp 1677622389
transform 1 0 2560 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_36
timestamp 1677622389
transform 1 0 2568 0 -1 4370
box -8 -3 46 105
use FILL  FILL_652
timestamp 1677622389
transform 1 0 2608 0 -1 4370
box -8 -3 16 105
use FILL  FILL_653
timestamp 1677622389
transform 1 0 2616 0 -1 4370
box -8 -3 16 105
use FILL  FILL_654
timestamp 1677622389
transform 1 0 2624 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1677622389
transform 1 0 2632 0 -1 4370
box -8 -3 46 105
use FILL  FILL_655
timestamp 1677622389
transform 1 0 2672 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_63
timestamp 1677622389
transform 1 0 2680 0 -1 4370
box -9 -3 26 105
use FILL  FILL_656
timestamp 1677622389
transform 1 0 2696 0 -1 4370
box -8 -3 16 105
use FILL  FILL_657
timestamp 1677622389
transform 1 0 2704 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1677622389
transform 1 0 2712 0 -1 4370
box -8 -3 104 105
use FILL  FILL_658
timestamp 1677622389
transform 1 0 2808 0 -1 4370
box -8 -3 16 105
use FILL  FILL_659
timestamp 1677622389
transform 1 0 2816 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1677622389
transform 1 0 2824 0 -1 4370
box -8 -3 32 105
use FILL  FILL_660
timestamp 1677622389
transform 1 0 2848 0 -1 4370
box -8 -3 16 105
use FILL  FILL_661
timestamp 1677622389
transform 1 0 2856 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_22
timestamp 1677622389
transform 1 0 2864 0 -1 4370
box -8 -3 34 105
use FILL  FILL_662
timestamp 1677622389
transform 1 0 2896 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1677622389
transform 1 0 2904 0 -1 4370
box -8 -3 32 105
use FILL  FILL_663
timestamp 1677622389
transform 1 0 2928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_664
timestamp 1677622389
transform 1 0 2936 0 -1 4370
box -8 -3 16 105
use FILL  FILL_665
timestamp 1677622389
transform 1 0 2944 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1677622389
transform 1 0 2952 0 -1 4370
box -8 -3 32 105
use FILL  FILL_666
timestamp 1677622389
transform 1 0 2976 0 -1 4370
box -8 -3 16 105
use FILL  FILL_667
timestamp 1677622389
transform 1 0 2984 0 -1 4370
box -8 -3 16 105
use FILL  FILL_668
timestamp 1677622389
transform 1 0 2992 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1677622389
transform -1 0 3032 0 -1 4370
box -8 -3 34 105
use FILL  FILL_669
timestamp 1677622389
transform 1 0 3032 0 -1 4370
box -8 -3 16 105
use FILL  FILL_670
timestamp 1677622389
transform 1 0 3040 0 -1 4370
box -8 -3 16 105
use FILL  FILL_671
timestamp 1677622389
transform 1 0 3048 0 -1 4370
box -8 -3 16 105
use FILL  FILL_672
timestamp 1677622389
transform 1 0 3056 0 -1 4370
box -8 -3 16 105
use FILL  FILL_673
timestamp 1677622389
transform 1 0 3064 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_31
timestamp 1677622389
transform -1 0 3112 0 -1 4370
box -8 -3 46 105
use FILL  FILL_674
timestamp 1677622389
transform 1 0 3112 0 -1 4370
box -8 -3 16 105
use FILL  FILL_675
timestamp 1677622389
transform 1 0 3120 0 -1 4370
box -8 -3 16 105
use FILL  FILL_676
timestamp 1677622389
transform 1 0 3128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_677
timestamp 1677622389
transform 1 0 3136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_678
timestamp 1677622389
transform 1 0 3144 0 -1 4370
box -8 -3 16 105
use FILL  FILL_679
timestamp 1677622389
transform 1 0 3152 0 -1 4370
box -8 -3 16 105
use FILL  FILL_680
timestamp 1677622389
transform 1 0 3160 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_32
timestamp 1677622389
transform -1 0 3208 0 -1 4370
box -8 -3 46 105
use INVX2  INVX2_64
timestamp 1677622389
transform -1 0 3224 0 -1 4370
box -9 -3 26 105
use FILL  FILL_681
timestamp 1677622389
transform 1 0 3224 0 -1 4370
box -8 -3 16 105
use FILL  FILL_682
timestamp 1677622389
transform 1 0 3232 0 -1 4370
box -8 -3 16 105
use FILL  FILL_683
timestamp 1677622389
transform 1 0 3240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_684
timestamp 1677622389
transform 1 0 3248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_685
timestamp 1677622389
transform 1 0 3256 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_65
timestamp 1677622389
transform -1 0 3280 0 -1 4370
box -9 -3 26 105
use FILL  FILL_686
timestamp 1677622389
transform 1 0 3280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_687
timestamp 1677622389
transform 1 0 3288 0 -1 4370
box -8 -3 16 105
use FILL  FILL_688
timestamp 1677622389
transform 1 0 3296 0 -1 4370
box -8 -3 16 105
use FILL  FILL_689
timestamp 1677622389
transform 1 0 3304 0 -1 4370
box -8 -3 16 105
use FILL  FILL_690
timestamp 1677622389
transform 1 0 3312 0 -1 4370
box -8 -3 16 105
use FILL  FILL_691
timestamp 1677622389
transform 1 0 3320 0 -1 4370
box -8 -3 16 105
use FILL  FILL_692
timestamp 1677622389
transform 1 0 3328 0 -1 4370
box -8 -3 16 105
use FILL  FILL_693
timestamp 1677622389
transform 1 0 3336 0 -1 4370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1677622389
transform 1 0 3344 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_66
timestamp 1677622389
transform 1 0 3352 0 -1 4370
box -9 -3 26 105
use FILL  FILL_695
timestamp 1677622389
transform 1 0 3368 0 -1 4370
box -8 -3 16 105
use FILL  FILL_697
timestamp 1677622389
transform 1 0 3376 0 -1 4370
box -8 -3 16 105
use FILL  FILL_699
timestamp 1677622389
transform 1 0 3384 0 -1 4370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1677622389
transform 1 0 3392 0 -1 4370
box -8 -3 16 105
use FILL  FILL_708
timestamp 1677622389
transform 1 0 3400 0 -1 4370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1677622389
transform 1 0 3408 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_33
timestamp 1677622389
transform -1 0 3456 0 -1 4370
box -8 -3 46 105
use FILL  FILL_710
timestamp 1677622389
transform 1 0 3456 0 -1 4370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1677622389
transform 1 0 3464 0 -1 4370
box -8 -3 16 105
use FILL  FILL_712
timestamp 1677622389
transform 1 0 3472 0 -1 4370
box -8 -3 16 105
use FILL  FILL_713
timestamp 1677622389
transform 1 0 3480 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_67
timestamp 1677622389
transform 1 0 3488 0 -1 4370
box -9 -3 26 105
use FILL  FILL_714
timestamp 1677622389
transform 1 0 3504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1677622389
transform 1 0 3512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_716
timestamp 1677622389
transform 1 0 3520 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_34
timestamp 1677622389
transform -1 0 3568 0 -1 4370
box -8 -3 46 105
use FILL  FILL_717
timestamp 1677622389
transform 1 0 3568 0 -1 4370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1677622389
transform 1 0 3576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_721
timestamp 1677622389
transform 1 0 3584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1677622389
transform 1 0 3592 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_35
timestamp 1677622389
transform 1 0 3600 0 -1 4370
box -8 -3 46 105
use FILL  FILL_724
timestamp 1677622389
transform 1 0 3640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1677622389
transform 1 0 3648 0 -1 4370
box -8 -3 16 105
use FILL  FILL_726
timestamp 1677622389
transform 1 0 3656 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_68
timestamp 1677622389
transform -1 0 3680 0 -1 4370
box -9 -3 26 105
use FILL  FILL_727
timestamp 1677622389
transform 1 0 3680 0 -1 4370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1677622389
transform 1 0 3688 0 -1 4370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1677622389
transform 1 0 3696 0 -1 4370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1677622389
transform 1 0 3704 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_38
timestamp 1677622389
transform -1 0 3752 0 -1 4370
box -8 -3 46 105
use FILL  FILL_736
timestamp 1677622389
transform 1 0 3752 0 -1 4370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1677622389
transform 1 0 3760 0 -1 4370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1677622389
transform 1 0 3768 0 -1 4370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1677622389
transform 1 0 3776 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_36
timestamp 1677622389
transform 1 0 3784 0 -1 4370
box -8 -3 46 105
use FILL  FILL_740
timestamp 1677622389
transform 1 0 3824 0 -1 4370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1677622389
transform 1 0 3832 0 -1 4370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1677622389
transform 1 0 3840 0 -1 4370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1677622389
transform 1 0 3848 0 -1 4370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1677622389
transform 1 0 3856 0 -1 4370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1677622389
transform 1 0 3864 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_754
timestamp 1677622389
transform 1 0 3884 0 1 4275
box -3 -3 3 3
use FILL  FILL_759
timestamp 1677622389
transform 1 0 3872 0 -1 4370
box -8 -3 16 105
use NAND3X1  NAND3X1_3
timestamp 1677622389
transform -1 0 3912 0 -1 4370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1677622389
transform -1 0 4008 0 -1 4370
box -8 -3 104 105
use M3_M2  M3_M2_755
timestamp 1677622389
transform 1 0 4028 0 1 4275
box -3 -3 3 3
use INVX2  INVX2_70
timestamp 1677622389
transform 1 0 4008 0 -1 4370
box -9 -3 26 105
use FILL  FILL_760
timestamp 1677622389
transform 1 0 4024 0 -1 4370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1677622389
transform 1 0 4032 0 -1 4370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1677622389
transform 1 0 4040 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1677622389
transform 1 0 4048 0 -1 4370
box -9 -3 26 105
use FILL  FILL_768
timestamp 1677622389
transform 1 0 4064 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_756
timestamp 1677622389
transform 1 0 4084 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_63
timestamp 1677622389
transform 1 0 4072 0 -1 4370
box -8 -3 104 105
use FILL  FILL_769
timestamp 1677622389
transform 1 0 4168 0 -1 4370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1677622389
transform 1 0 4176 0 -1 4370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1677622389
transform 1 0 4184 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_757
timestamp 1677622389
transform 1 0 4220 0 1 4275
box -3 -3 3 3
use OAI22X1  OAI22X1_38
timestamp 1677622389
transform 1 0 4192 0 -1 4370
box -8 -3 46 105
use FILL  FILL_772
timestamp 1677622389
transform 1 0 4232 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_72
timestamp 1677622389
transform -1 0 4256 0 -1 4370
box -9 -3 26 105
use FILL  FILL_773
timestamp 1677622389
transform 1 0 4256 0 -1 4370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1677622389
transform 1 0 4264 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_40
timestamp 1677622389
transform 1 0 4272 0 -1 4370
box -8 -3 46 105
use FILL  FILL_784
timestamp 1677622389
transform 1 0 4312 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_41
timestamp 1677622389
transform 1 0 4320 0 -1 4370
box -8 -3 46 105
use FILL  FILL_785
timestamp 1677622389
transform 1 0 4360 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_41
timestamp 1677622389
transform -1 0 4408 0 -1 4370
box -8 -3 46 105
use FILL  FILL_786
timestamp 1677622389
transform 1 0 4408 0 -1 4370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1677622389
transform 1 0 4416 0 -1 4370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1677622389
transform 1 0 4424 0 -1 4370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1677622389
transform 1 0 4432 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1677622389
transform 1 0 4440 0 -1 4370
box -8 -3 46 105
use FILL  FILL_790
timestamp 1677622389
transform 1 0 4480 0 -1 4370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1677622389
transform 1 0 4488 0 -1 4370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1677622389
transform 1 0 4496 0 -1 4370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1677622389
transform 1 0 4504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1677622389
transform 1 0 4512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1677622389
transform 1 0 4520 0 -1 4370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1677622389
transform 1 0 4528 0 -1 4370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1677622389
transform 1 0 4536 0 -1 4370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1677622389
transform 1 0 4544 0 -1 4370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1677622389
transform 1 0 4552 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1677622389
transform 1 0 4560 0 -1 4370
box -8 -3 104 105
use FILL  FILL_800
timestamp 1677622389
transform 1 0 4656 0 -1 4370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1677622389
transform 1 0 4664 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1677622389
transform 1 0 4672 0 -1 4370
box -8 -3 104 105
use FILL  FILL_802
timestamp 1677622389
transform 1 0 4768 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1677622389
transform 1 0 4776 0 -1 4370
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_9
timestamp 1677622389
transform 1 0 4843 0 1 4270
box -10 -3 10 3
use M3_M2  M3_M2_869
timestamp 1677622389
transform 1 0 84 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1677622389
transform 1 0 116 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1677622389
transform 1 0 164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1677622389
transform 1 0 84 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_778
timestamp 1677622389
transform 1 0 188 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_934
timestamp 1677622389
transform 1 0 244 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_904
timestamp 1677622389
transform 1 0 244 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1677622389
transform 1 0 300 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_935
timestamp 1677622389
transform 1 0 308 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1677622389
transform 1 0 332 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_905
timestamp 1677622389
transform 1 0 332 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1677622389
transform 1 0 380 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1677622389
transform 1 0 364 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_936
timestamp 1677622389
transform 1 0 396 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_871
timestamp 1677622389
transform 1 0 412 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1054
timestamp 1677622389
transform 1 0 364 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_906
timestamp 1677622389
transform 1 0 388 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1055
timestamp 1677622389
transform 1 0 460 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1677622389
transform 1 0 500 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_907
timestamp 1677622389
transform 1 0 500 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_938
timestamp 1677622389
transform 1 0 532 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1677622389
transform 1 0 548 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1677622389
transform 1 0 524 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1677622389
transform 1 0 556 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1677622389
transform 1 0 572 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1677622389
transform 1 0 572 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_940
timestamp 1677622389
transform 1 0 572 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1677622389
transform 1 0 540 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1677622389
transform 1 0 556 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1677622389
transform 1 0 564 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_955
timestamp 1677622389
transform 1 0 532 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1677622389
transform 1 0 596 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1677622389
transform 1 0 604 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1677622389
transform 1 0 612 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_941
timestamp 1677622389
transform 1 0 612 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_758
timestamp 1677622389
transform 1 0 628 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1677622389
transform 1 0 652 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1677622389
transform 1 0 652 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1677622389
transform 1 0 652 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1677622389
transform 1 0 700 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1677622389
transform 1 0 716 0 1 4265
box -3 -3 3 3
use M2_M1  M2_M1_943
timestamp 1677622389
transform 1 0 708 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1677622389
transform 1 0 628 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_822
timestamp 1677622389
transform 1 0 740 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1677622389
transform 1 0 748 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1677622389
transform 1 0 740 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1677622389
transform 1 0 748 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_908
timestamp 1677622389
transform 1 0 748 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1677622389
transform 1 0 756 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_945
timestamp 1677622389
transform 1 0 772 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1677622389
transform 1 0 788 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_874
timestamp 1677622389
transform 1 0 796 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1677622389
transform 1 0 780 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_891
timestamp 1677622389
transform 1 0 788 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1677622389
transform 1 0 796 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_772
timestamp 1677622389
transform 1 0 812 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1677622389
transform 1 0 844 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1677622389
transform 1 0 836 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_947
timestamp 1677622389
transform 1 0 868 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1677622389
transform 1 0 836 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_825
timestamp 1677622389
transform 1 0 924 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1160
timestamp 1677622389
transform 1 0 924 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1677622389
transform 1 0 948 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_892
timestamp 1677622389
transform 1 0 964 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1161
timestamp 1677622389
transform 1 0 964 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1677622389
transform 1 0 1004 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1677622389
transform 1 0 1004 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1677622389
transform 1 0 1028 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_760
timestamp 1677622389
transform 1 0 1060 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1677622389
transform 1 0 1076 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1677622389
transform 1 0 1060 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1677622389
transform 1 0 1076 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1677622389
transform 1 0 1060 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1677622389
transform 1 0 1100 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1677622389
transform 1 0 1092 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1068
timestamp 1677622389
transform 1 0 1092 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1677622389
transform 1 0 1108 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_951
timestamp 1677622389
transform 1 0 1108 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_783
timestamp 1677622389
transform 1 0 1132 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1677622389
transform 1 0 1140 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_952
timestamp 1677622389
transform 1 0 1132 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1677622389
transform 1 0 1148 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1677622389
transform 1 0 1116 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1677622389
transform 1 0 1140 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1677622389
transform 1 0 1148 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_956
timestamp 1677622389
transform 1 0 1108 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1677622389
transform 1 0 1188 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_920
timestamp 1677622389
transform 1 0 1196 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1677622389
transform 1 0 1196 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_910
timestamp 1677622389
transform 1 0 1196 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1677622389
transform 1 0 1236 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_921
timestamp 1677622389
transform 1 0 1236 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_829
timestamp 1677622389
transform 1 0 1252 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_954
timestamp 1677622389
transform 1 0 1252 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_830
timestamp 1677622389
transform 1 0 1276 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_955
timestamp 1677622389
transform 1 0 1276 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_785
timestamp 1677622389
transform 1 0 1292 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_922
timestamp 1677622389
transform 1 0 1292 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1677622389
transform 1 0 1316 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_831
timestamp 1677622389
transform 1 0 1324 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1073
timestamp 1677622389
transform 1 0 1324 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_832
timestamp 1677622389
transform 1 0 1356 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_956
timestamp 1677622389
transform 1 0 1332 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1677622389
transform 1 0 1348 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1677622389
transform 1 0 1356 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1677622389
transform 1 0 1332 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1677622389
transform 1 0 1356 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1677622389
transform 1 0 1364 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_911
timestamp 1677622389
transform 1 0 1356 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1677622389
transform 1 0 1404 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1677622389
transform 1 0 1404 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1677622389
transform 1 0 1428 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1677622389
transform 1 0 1436 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1677622389
transform 1 0 1396 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1677622389
transform 1 0 1412 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1677622389
transform 1 0 1420 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1677622389
transform 1 0 1428 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_912
timestamp 1677622389
transform 1 0 1404 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1677622389
transform 1 0 1436 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1080
timestamp 1677622389
transform 1 0 1452 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_957
timestamp 1677622389
transform 1 0 1444 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1081
timestamp 1677622389
transform 1 0 1460 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_834
timestamp 1677622389
transform 1 0 1492 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1677622389
transform 1 0 1516 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_962
timestamp 1677622389
transform 1 0 1492 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1677622389
transform 1 0 1508 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1677622389
transform 1 0 1516 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1677622389
transform 1 0 1500 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_958
timestamp 1677622389
transform 1 0 1508 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1677622389
transform 1 0 1540 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1677622389
transform 1 0 1564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1677622389
transform 1 0 1556 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_761
timestamp 1677622389
transform 1 0 1572 0 1 4265
box -3 -3 3 3
use M2_M1  M2_M1_1085
timestamp 1677622389
transform 1 0 1572 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_775
timestamp 1677622389
transform 1 0 1692 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_966
timestamp 1677622389
transform 1 0 1612 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1677622389
transform 1 0 1644 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1677622389
transform 1 0 1692 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1677622389
transform 1 0 1620 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1677622389
transform 1 0 1644 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1677622389
transform 1 0 1708 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1677622389
transform 1 0 1716 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1677622389
transform 1 0 1812 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1677622389
transform 1 0 1860 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1677622389
transform 1 0 1828 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1677622389
transform 1 0 1844 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_968
timestamp 1677622389
transform 1 0 1788 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1677622389
transform 1 0 1820 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1677622389
transform 1 0 1828 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1677622389
transform 1 0 1844 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1677622389
transform 1 0 1860 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1677622389
transform 1 0 1868 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1677622389
transform 1 0 1740 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1677622389
transform 1 0 1828 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1677622389
transform 1 0 1836 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1677622389
transform 1 0 1852 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1677622389
transform 1 0 1740 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1677622389
transform 1 0 1788 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1677622389
transform 1 0 1820 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1677622389
transform 1 0 1852 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1677622389
transform 1 0 1868 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1677622389
transform 1 0 1884 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1677622389
transform 1 0 1900 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_974
timestamp 1677622389
transform 1 0 1908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1677622389
transform 1 0 1900 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_894
timestamp 1677622389
transform 1 0 1908 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1677622389
transform 1 0 1932 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1677622389
transform 1 0 1924 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1092
timestamp 1677622389
transform 1 0 1924 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1677622389
transform 1 0 1940 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1677622389
transform 1 0 1980 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1677622389
transform 1 0 1964 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_976
timestamp 1677622389
transform 1 0 1988 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1677622389
transform 1 0 1956 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_961
timestamp 1677622389
transform 1 0 1956 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1677622389
transform 1 0 1996 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_977
timestamp 1677622389
transform 1 0 2004 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_895
timestamp 1677622389
transform 1 0 1972 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1094
timestamp 1677622389
transform 1 0 1980 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_962
timestamp 1677622389
transform 1 0 1972 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1677622389
transform 1 0 2012 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_978
timestamp 1677622389
transform 1 0 2044 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1677622389
transform 1 0 2060 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1677622389
transform 1 0 2028 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1677622389
transform 1 0 2036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1677622389
transform 1 0 2052 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1677622389
transform 1 0 2148 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1677622389
transform 1 0 2180 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_920
timestamp 1677622389
transform 1 0 2180 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1677622389
transform 1 0 2204 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_921
timestamp 1677622389
transform 1 0 2220 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1677622389
transform 1 0 2244 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1677622389
transform 1 0 2244 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_897
timestamp 1677622389
transform 1 0 2244 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1677622389
transform 1 0 2260 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1677622389
transform 1 0 2284 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1677622389
transform 1 0 2260 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1677622389
transform 1 0 2284 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1677622389
transform 1 0 2340 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1677622389
transform 1 0 2260 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_766
timestamp 1677622389
transform 1 0 2396 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1677622389
transform 1 0 2396 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1677622389
transform 1 0 2364 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1677622389
transform 1 0 2380 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1677622389
transform 1 0 2396 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1677622389
transform 1 0 2372 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1677622389
transform 1 0 2388 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_922
timestamp 1677622389
transform 1 0 2372 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1677622389
transform 1 0 2412 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1677622389
transform 1 0 2404 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_987
timestamp 1677622389
transform 1 0 2452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1677622389
transform 1 0 2468 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1677622389
transform 1 0 2460 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1677622389
transform 1 0 2476 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_924
timestamp 1677622389
transform 1 0 2476 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1677622389
transform 1 0 2604 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_989
timestamp 1677622389
transform 1 0 2540 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1677622389
transform 1 0 2596 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1677622389
transform 1 0 2604 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1677622389
transform 1 0 2516 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_925
timestamp 1677622389
transform 1 0 2532 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1677622389
transform 1 0 2644 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1677622389
transform 1 0 2636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1677622389
transform 1 0 2660 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1677622389
transform 1 0 2628 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1677622389
transform 1 0 2644 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1677622389
transform 1 0 2652 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1677622389
transform 1 0 2676 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_843
timestamp 1677622389
transform 1 0 2708 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1677622389
transform 1 0 2708 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_790
timestamp 1677622389
transform 1 0 2804 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1677622389
transform 1 0 2748 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1677622389
transform 1 0 2812 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_996
timestamp 1677622389
transform 1 0 2748 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1677622389
transform 1 0 2804 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1677622389
transform 1 0 2724 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_926
timestamp 1677622389
transform 1 0 2740 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1677622389
transform 1 0 2820 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1677622389
transform 1 0 2820 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_846
timestamp 1677622389
transform 1 0 2860 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_924
timestamp 1677622389
transform 1 0 2868 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_878
timestamp 1677622389
transform 1 0 2868 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1111
timestamp 1677622389
transform 1 0 2868 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1677622389
transform 1 0 2860 0 1 4195
box -2 -2 2 2
use M3_M2  M3_M2_927
timestamp 1677622389
transform 1 0 2868 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1677622389
transform 1 0 2884 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_999
timestamp 1677622389
transform 1 0 2892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1677622389
transform 1 0 2884 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1677622389
transform 1 0 2900 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_928
timestamp 1677622389
transform 1 0 2892 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1677622389
transform 1 0 2924 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_847
timestamp 1677622389
transform 1 0 2940 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1677622389
transform 1 0 2940 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_929
timestamp 1677622389
transform 1 0 2924 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1677622389
transform 1 0 2956 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1677622389
transform 1 0 2964 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_926
timestamp 1677622389
transform 1 0 2972 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_879
timestamp 1677622389
transform 1 0 2956 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1114
timestamp 1677622389
transform 1 0 2956 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1677622389
transform 1 0 2980 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_849
timestamp 1677622389
transform 1 0 2996 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1677622389
transform 1 0 2980 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1677622389
transform 1 0 2996 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1677622389
transform 1 0 2980 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1677622389
transform 1 0 2972 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1677622389
transform 1 0 3020 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1677622389
transform 1 0 3036 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1677622389
transform 1 0 3028 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1677622389
transform 1 0 3044 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1677622389
transform 1 0 3060 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1677622389
transform 1 0 3028 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1677622389
transform 1 0 3036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1677622389
transform 1 0 3052 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1677622389
transform 1 0 3060 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1677622389
transform 1 0 3092 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1005
timestamp 1677622389
transform 1 0 3084 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1677622389
transform 1 0 3084 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_931
timestamp 1677622389
transform 1 0 3084 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1677622389
transform 1 0 3148 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1677622389
transform 1 0 3204 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1006
timestamp 1677622389
transform 1 0 3148 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1677622389
transform 1 0 3204 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1677622389
transform 1 0 3188 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1677622389
transform 1 0 3204 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_881
timestamp 1677622389
transform 1 0 3228 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1677622389
transform 1 0 3260 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1008
timestamp 1677622389
transform 1 0 3236 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1677622389
transform 1 0 3260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1677622389
transform 1 0 3220 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_932
timestamp 1677622389
transform 1 0 3116 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1677622389
transform 1 0 3204 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1677622389
transform 1 0 3220 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1677622389
transform 1 0 3244 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1677622389
transform 1 0 3244 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1677622389
transform 1 0 3276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1677622389
transform 1 0 3276 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_963
timestamp 1677622389
transform 1 0 3276 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1677622389
transform 1 0 3316 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1677622389
transform 1 0 3364 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_936
timestamp 1677622389
transform 1 0 3316 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1677622389
transform 1 0 3388 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1677622389
transform 1 0 3412 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_917
timestamp 1677622389
transform 1 0 3412 0 1 4235
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1677622389
transform 1 0 3412 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1012
timestamp 1677622389
transform 1 0 3412 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_882
timestamp 1677622389
transform 1 0 3428 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1677622389
transform 1 0 3452 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1125
timestamp 1677622389
transform 1 0 3436 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_900
timestamp 1677622389
transform 1 0 3444 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1677622389
transform 1 0 3468 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_929
timestamp 1677622389
transform 1 0 3460 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1677622389
transform 1 0 3468 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_883
timestamp 1677622389
transform 1 0 3476 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1677622389
transform 1 0 3484 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_884
timestamp 1677622389
transform 1 0 3500 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1126
timestamp 1677622389
transform 1 0 3500 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_937
timestamp 1677622389
transform 1 0 3468 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1677622389
transform 1 0 3492 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1677622389
transform 1 0 3516 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1677622389
transform 1 0 3532 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1677622389
transform 1 0 3524 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_856
timestamp 1677622389
transform 1 0 3556 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1677622389
transform 1 0 3540 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1677622389
transform 1 0 3556 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1677622389
transform 1 0 3572 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1677622389
transform 1 0 3580 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1677622389
transform 1 0 3540 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1677622389
transform 1 0 3572 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1677622389
transform 1 0 3596 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1677622389
transform 1 0 3596 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1677622389
transform 1 0 3628 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1677622389
transform 1 0 3644 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1019
timestamp 1677622389
transform 1 0 3612 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1677622389
transform 1 0 3628 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_886
timestamp 1677622389
transform 1 0 3636 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1677622389
transform 1 0 3644 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1677622389
transform 1 0 3596 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1677622389
transform 1 0 3604 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1677622389
transform 1 0 3620 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1677622389
transform 1 0 3636 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_940
timestamp 1677622389
transform 1 0 3604 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1677622389
transform 1 0 3620 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1677622389
transform 1 0 3612 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1677622389
transform 1 0 3652 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_794
timestamp 1677622389
transform 1 0 3732 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1677622389
transform 1 0 3772 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1677622389
transform 1 0 3724 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1022
timestamp 1677622389
transform 1 0 3724 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1677622389
transform 1 0 3772 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_942
timestamp 1677622389
transform 1 0 3724 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1677622389
transform 1 0 3796 0 1 4265
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1677622389
transform 1 0 3788 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1677622389
transform 1 0 3812 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1677622389
transform 1 0 3820 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_887
timestamp 1677622389
transform 1 0 3828 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1677622389
transform 1 0 3844 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1677622389
transform 1 0 3836 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1677622389
transform 1 0 3812 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_901
timestamp 1677622389
transform 1 0 3820 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1677622389
transform 1 0 3884 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1677622389
transform 1 0 3900 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1677622389
transform 1 0 3868 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1677622389
transform 1 0 3892 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1026
timestamp 1677622389
transform 1 0 3868 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1677622389
transform 1 0 3884 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1677622389
transform 1 0 3892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1677622389
transform 1 0 3852 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1677622389
transform 1 0 3860 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1677622389
transform 1 0 3876 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1677622389
transform 1 0 3892 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_943
timestamp 1677622389
transform 1 0 3852 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1677622389
transform 1 0 3900 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1029
timestamp 1677622389
transform 1 0 3932 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1677622389
transform 1 0 3924 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_945
timestamp 1677622389
transform 1 0 3932 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1677622389
transform 1 0 3996 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1677622389
transform 1 0 4020 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1677622389
transform 1 0 4092 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_1140
timestamp 1677622389
transform 1 0 3988 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_946
timestamp 1677622389
transform 1 0 3988 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1030
timestamp 1677622389
transform 1 0 4052 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1677622389
transform 1 0 4084 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1677622389
transform 1 0 4092 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1677622389
transform 1 0 4100 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1677622389
transform 1 0 4116 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1677622389
transform 1 0 4132 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1677622389
transform 1 0 4004 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1677622389
transform 1 0 4092 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1677622389
transform 1 0 4108 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1677622389
transform 1 0 4124 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_947
timestamp 1677622389
transform 1 0 4028 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1677622389
transform 1 0 4052 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1677622389
transform 1 0 4108 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1145
timestamp 1677622389
transform 1 0 4172 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_888
timestamp 1677622389
transform 1 0 4204 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1036
timestamp 1677622389
transform 1 0 4212 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_863
timestamp 1677622389
transform 1 0 4244 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1037
timestamp 1677622389
transform 1 0 4244 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1677622389
transform 1 0 4260 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_799
timestamp 1677622389
transform 1 0 4276 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1677622389
transform 1 0 4308 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1677622389
transform 1 0 4300 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1677622389
transform 1 0 4292 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_918
timestamp 1677622389
transform 1 0 4308 0 1 4235
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1677622389
transform 1 0 4284 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1677622389
transform 1 0 4276 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_950
timestamp 1677622389
transform 1 0 4268 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1677622389
transform 1 0 4300 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_931
timestamp 1677622389
transform 1 0 4308 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1677622389
transform 1 0 4308 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_902
timestamp 1677622389
transform 1 0 4308 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1677622389
transform 1 0 4388 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1677622389
transform 1 0 4380 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1040
timestamp 1677622389
transform 1 0 4380 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1677622389
transform 1 0 4356 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1677622389
transform 1 0 4452 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1677622389
transform 1 0 4460 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_1041
timestamp 1677622389
transform 1 0 4452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1677622389
transform 1 0 4460 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1677622389
transform 1 0 4476 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_819
timestamp 1677622389
transform 1 0 4516 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1677622389
transform 1 0 4508 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1677622389
transform 1 0 4492 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_889
timestamp 1677622389
transform 1 0 4500 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1044
timestamp 1677622389
transform 1 0 4508 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1677622389
transform 1 0 4532 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1677622389
transform 1 0 4548 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1677622389
transform 1 0 4484 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1677622389
transform 1 0 4500 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1677622389
transform 1 0 4516 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1677622389
transform 1 0 4524 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_951
timestamp 1677622389
transform 1 0 4484 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1677622389
transform 1 0 4548 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1153
timestamp 1677622389
transform 1 0 4556 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1677622389
transform 1 0 4556 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1677622389
transform 1 0 4580 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1047
timestamp 1677622389
transform 1 0 4580 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1677622389
transform 1 0 4572 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_890
timestamp 1677622389
transform 1 0 4596 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1048
timestamp 1677622389
transform 1 0 4604 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_953
timestamp 1677622389
transform 1 0 4612 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1677622389
transform 1 0 4604 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1677622389
transform 1 0 4684 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1677622389
transform 1 0 4668 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1049
timestamp 1677622389
transform 1 0 4668 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1677622389
transform 1 0 4692 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1677622389
transform 1 0 4652 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1677622389
transform 1 0 4660 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_967
timestamp 1677622389
transform 1 0 4652 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1677622389
transform 1 0 4716 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1677622389
transform 1 0 4708 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1051
timestamp 1677622389
transform 1 0 4708 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1677622389
transform 1 0 4684 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1677622389
transform 1 0 4700 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_954
timestamp 1677622389
transform 1 0 4692 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1159
timestamp 1677622389
transform 1 0 4724 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_968
timestamp 1677622389
transform 1 0 4764 0 1 4185
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_10
timestamp 1677622389
transform 1 0 48 0 1 4170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1677622389
transform 1 0 72 0 1 4170
box -8 -3 104 105
use FILL  FILL_803
timestamp 1677622389
transform 1 0 168 0 1 4170
box -8 -3 16 105
use FILL  FILL_804
timestamp 1677622389
transform 1 0 176 0 1 4170
box -8 -3 16 105
use FILL  FILL_805
timestamp 1677622389
transform 1 0 184 0 1 4170
box -8 -3 16 105
use FILL  FILL_806
timestamp 1677622389
transform 1 0 192 0 1 4170
box -8 -3 16 105
use FILL  FILL_807
timestamp 1677622389
transform 1 0 200 0 1 4170
box -8 -3 16 105
use FILL  FILL_818
timestamp 1677622389
transform 1 0 208 0 1 4170
box -8 -3 16 105
use FILL  FILL_819
timestamp 1677622389
transform 1 0 216 0 1 4170
box -8 -3 16 105
use FILL  FILL_820
timestamp 1677622389
transform 1 0 224 0 1 4170
box -8 -3 16 105
use FILL  FILL_821
timestamp 1677622389
transform 1 0 232 0 1 4170
box -8 -3 16 105
use FILL  FILL_822
timestamp 1677622389
transform 1 0 240 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1677622389
transform -1 0 344 0 1 4170
box -8 -3 104 105
use FILL  FILL_823
timestamp 1677622389
transform 1 0 344 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1677622389
transform 1 0 352 0 1 4170
box -8 -3 104 105
use FILL  FILL_826
timestamp 1677622389
transform 1 0 448 0 1 4170
box -8 -3 16 105
use FILL  FILL_838
timestamp 1677622389
transform 1 0 456 0 1 4170
box -8 -3 16 105
use FILL  FILL_840
timestamp 1677622389
transform 1 0 464 0 1 4170
box -8 -3 16 105
use FILL  FILL_841
timestamp 1677622389
transform 1 0 472 0 1 4170
box -8 -3 16 105
use FILL  FILL_842
timestamp 1677622389
transform 1 0 480 0 1 4170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1677622389
transform 1 0 488 0 1 4170
box -8 -3 16 105
use FILL  FILL_844
timestamp 1677622389
transform 1 0 496 0 1 4170
box -8 -3 16 105
use FILL  FILL_845
timestamp 1677622389
transform 1 0 504 0 1 4170
box -8 -3 16 105
use FILL  FILL_847
timestamp 1677622389
transform 1 0 512 0 1 4170
box -8 -3 16 105
use FILL  FILL_849
timestamp 1677622389
transform 1 0 520 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_45
timestamp 1677622389
transform 1 0 528 0 1 4170
box -8 -3 46 105
use FILL  FILL_851
timestamp 1677622389
transform 1 0 568 0 1 4170
box -8 -3 16 105
use FILL  FILL_853
timestamp 1677622389
transform 1 0 576 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_81
timestamp 1677622389
transform 1 0 584 0 1 4170
box -9 -3 26 105
use FILL  FILL_855
timestamp 1677622389
transform 1 0 600 0 1 4170
box -8 -3 16 105
use FILL  FILL_857
timestamp 1677622389
transform 1 0 608 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1677622389
transform 1 0 616 0 1 4170
box -8 -3 104 105
use FILL  FILL_859
timestamp 1677622389
transform 1 0 712 0 1 4170
box -8 -3 16 105
use FILL  FILL_860
timestamp 1677622389
transform 1 0 720 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_83
timestamp 1677622389
transform -1 0 744 0 1 4170
box -9 -3 26 105
use FILL  FILL_861
timestamp 1677622389
transform 1 0 744 0 1 4170
box -8 -3 16 105
use FILL  FILL_867
timestamp 1677622389
transform 1 0 752 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_43
timestamp 1677622389
transform 1 0 760 0 1 4170
box -8 -3 46 105
use FILL  FILL_869
timestamp 1677622389
transform 1 0 800 0 1 4170
box -8 -3 16 105
use FILL  FILL_870
timestamp 1677622389
transform 1 0 808 0 1 4170
box -8 -3 16 105
use FILL  FILL_871
timestamp 1677622389
transform 1 0 816 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1677622389
transform 1 0 824 0 1 4170
box -8 -3 104 105
use FILL  FILL_872
timestamp 1677622389
transform 1 0 920 0 1 4170
box -8 -3 16 105
use FILL  FILL_887
timestamp 1677622389
transform 1 0 928 0 1 4170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1677622389
transform 1 0 936 0 1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1677622389
transform 1 0 944 0 1 4170
box -8 -3 32 105
use FILL  FILL_890
timestamp 1677622389
transform 1 0 968 0 1 4170
box -8 -3 16 105
use FILL  FILL_891
timestamp 1677622389
transform 1 0 976 0 1 4170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1677622389
transform 1 0 984 0 1 4170
box -8 -3 16 105
use FILL  FILL_895
timestamp 1677622389
transform 1 0 992 0 1 4170
box -8 -3 16 105
use FILL  FILL_897
timestamp 1677622389
transform 1 0 1000 0 1 4170
box -8 -3 16 105
use FILL  FILL_899
timestamp 1677622389
transform 1 0 1008 0 1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1677622389
transform 1 0 1016 0 1 4170
box -8 -3 32 105
use FILL  FILL_900
timestamp 1677622389
transform 1 0 1040 0 1 4170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1677622389
transform 1 0 1048 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1677622389
transform -1 0 1088 0 1 4170
box -8 -3 34 105
use FILL  FILL_903
timestamp 1677622389
transform 1 0 1088 0 1 4170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1677622389
transform 1 0 1096 0 1 4170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1677622389
transform 1 0 1104 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_48
timestamp 1677622389
transform 1 0 1112 0 1 4170
box -8 -3 46 105
use FILL  FILL_906
timestamp 1677622389
transform 1 0 1152 0 1 4170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1677622389
transform 1 0 1160 0 1 4170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1677622389
transform 1 0 1168 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_85
timestamp 1677622389
transform 1 0 1176 0 1 4170
box -9 -3 26 105
use FILL  FILL_909
timestamp 1677622389
transform 1 0 1192 0 1 4170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1677622389
transform 1 0 1200 0 1 4170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1677622389
transform 1 0 1208 0 1 4170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1677622389
transform 1 0 1216 0 1 4170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1677622389
transform 1 0 1224 0 1 4170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1677622389
transform 1 0 1232 0 1 4170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1677622389
transform 1 0 1240 0 1 4170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1677622389
transform 1 0 1248 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1677622389
transform -1 0 1288 0 1 4170
box -8 -3 34 105
use FILL  FILL_917
timestamp 1677622389
transform 1 0 1288 0 1 4170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1677622389
transform 1 0 1296 0 1 4170
box -8 -3 16 105
use FILL  FILL_932
timestamp 1677622389
transform 1 0 1304 0 1 4170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1677622389
transform 1 0 1312 0 1 4170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1677622389
transform 1 0 1320 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_28
timestamp 1677622389
transform -1 0 1360 0 1 4170
box -8 -3 34 105
use INVX2  INVX2_86
timestamp 1677622389
transform 1 0 1360 0 1 4170
box -9 -3 26 105
use FILL  FILL_937
timestamp 1677622389
transform 1 0 1376 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_969
timestamp 1677622389
transform 1 0 1396 0 1 4175
box -3 -3 3 3
use FILL  FILL_942
timestamp 1677622389
transform 1 0 1384 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_45
timestamp 1677622389
transform -1 0 1432 0 1 4170
box -8 -3 46 105
use INVX2  INVX2_87
timestamp 1677622389
transform -1 0 1448 0 1 4170
box -9 -3 26 105
use M3_M2  M3_M2_970
timestamp 1677622389
transform 1 0 1460 0 1 4175
box -3 -3 3 3
use FILL  FILL_944
timestamp 1677622389
transform 1 0 1448 0 1 4170
box -8 -3 16 105
use FILL  FILL_945
timestamp 1677622389
transform 1 0 1456 0 1 4170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1677622389
transform 1 0 1464 0 1 4170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1677622389
transform 1 0 1472 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_46
timestamp 1677622389
transform -1 0 1520 0 1 4170
box -8 -3 46 105
use FILL  FILL_948
timestamp 1677622389
transform 1 0 1520 0 1 4170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1677622389
transform 1 0 1528 0 1 4170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1677622389
transform 1 0 1536 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_88
timestamp 1677622389
transform -1 0 1560 0 1 4170
box -9 -3 26 105
use FILL  FILL_951
timestamp 1677622389
transform 1 0 1560 0 1 4170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1677622389
transform 1 0 1568 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_89
timestamp 1677622389
transform 1 0 1576 0 1 4170
box -9 -3 26 105
use FILL  FILL_959
timestamp 1677622389
transform 1 0 1592 0 1 4170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1677622389
transform 1 0 1600 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1677622389
transform -1 0 1704 0 1 4170
box -8 -3 104 105
use FILL  FILL_961
timestamp 1677622389
transform 1 0 1704 0 1 4170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1677622389
transform 1 0 1712 0 1 4170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1677622389
transform 1 0 1720 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_971
timestamp 1677622389
transform 1 0 1772 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1677622389
transform 1 0 1828 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_79
timestamp 1677622389
transform 1 0 1728 0 1 4170
box -8 -3 104 105
use AOI22X1  AOI22X1_49
timestamp 1677622389
transform 1 0 1824 0 1 4170
box -8 -3 46 105
use FILL  FILL_976
timestamp 1677622389
transform 1 0 1864 0 1 4170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1677622389
transform 1 0 1872 0 1 4170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1677622389
transform 1 0 1880 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_91
timestamp 1677622389
transform -1 0 1904 0 1 4170
box -9 -3 26 105
use FILL  FILL_979
timestamp 1677622389
transform 1 0 1904 0 1 4170
box -8 -3 16 105
use FILL  FILL_996
timestamp 1677622389
transform 1 0 1912 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_93
timestamp 1677622389
transform 1 0 1920 0 1 4170
box -9 -3 26 105
use FILL  FILL_998
timestamp 1677622389
transform 1 0 1936 0 1 4170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1677622389
transform 1 0 1944 0 1 4170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1677622389
transform 1 0 1952 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_49
timestamp 1677622389
transform 1 0 1960 0 1 4170
box -8 -3 46 105
use FILL  FILL_1001
timestamp 1677622389
transform 1 0 2000 0 1 4170
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1677622389
transform 1 0 2008 0 1 4170
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1677622389
transform 1 0 2016 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_51
timestamp 1677622389
transform 1 0 2024 0 1 4170
box -8 -3 46 105
use FILL  FILL_1011
timestamp 1677622389
transform 1 0 2064 0 1 4170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1677622389
transform 1 0 2072 0 1 4170
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1677622389
transform 1 0 2080 0 1 4170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1677622389
transform 1 0 2088 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_973
timestamp 1677622389
transform 1 0 2180 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_80
timestamp 1677622389
transform -1 0 2192 0 1 4170
box -8 -3 104 105
use M3_M2  M3_M2_974
timestamp 1677622389
transform 1 0 2204 0 1 4175
box -3 -3 3 3
use FILL  FILL_1015
timestamp 1677622389
transform 1 0 2192 0 1 4170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1677622389
transform 1 0 2200 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_94
timestamp 1677622389
transform 1 0 2208 0 1 4170
box -9 -3 26 105
use FILL  FILL_1024
timestamp 1677622389
transform 1 0 2224 0 1 4170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1677622389
transform 1 0 2232 0 1 4170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1677622389
transform 1 0 2240 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1677622389
transform 1 0 2248 0 1 4170
box -8 -3 104 105
use FILL  FILL_1031
timestamp 1677622389
transform 1 0 2344 0 1 4170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1677622389
transform 1 0 2352 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_53
timestamp 1677622389
transform -1 0 2400 0 1 4170
box -8 -3 46 105
use FILL  FILL_1033
timestamp 1677622389
transform 1 0 2400 0 1 4170
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1677622389
transform 1 0 2408 0 1 4170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1677622389
transform 1 0 2416 0 1 4170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1677622389
transform 1 0 2424 0 1 4170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1677622389
transform 1 0 2432 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_975
timestamp 1677622389
transform 1 0 2460 0 1 4175
box -3 -3 3 3
use OAI22X1  OAI22X1_51
timestamp 1677622389
transform -1 0 2480 0 1 4170
box -8 -3 46 105
use FILL  FILL_1038
timestamp 1677622389
transform 1 0 2480 0 1 4170
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1677622389
transform 1 0 2488 0 1 4170
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1677622389
transform 1 0 2496 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1677622389
transform 1 0 2504 0 1 4170
box -8 -3 104 105
use FILL  FILL_1041
timestamp 1677622389
transform 1 0 2600 0 1 4170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1677622389
transform 1 0 2608 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_54
timestamp 1677622389
transform 1 0 2616 0 1 4170
box -8 -3 46 105
use FILL  FILL_1043
timestamp 1677622389
transform 1 0 2656 0 1 4170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1677622389
transform 1 0 2664 0 1 4170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1677622389
transform 1 0 2672 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_95
timestamp 1677622389
transform 1 0 2680 0 1 4170
box -9 -3 26 105
use FILL  FILL_1046
timestamp 1677622389
transform 1 0 2696 0 1 4170
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1677622389
transform 1 0 2704 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1677622389
transform 1 0 2712 0 1 4170
box -8 -3 104 105
use FILL  FILL_1063
timestamp 1677622389
transform 1 0 2808 0 1 4170
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1677622389
transform 1 0 2816 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_976
timestamp 1677622389
transform 1 0 2860 0 1 4175
box -3 -3 3 3
use OAI21X1  OAI21X1_30
timestamp 1677622389
transform 1 0 2824 0 1 4170
box -8 -3 34 105
use FILL  FILL_1066
timestamp 1677622389
transform 1 0 2856 0 1 4170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1677622389
transform 1 0 2864 0 1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1677622389
transform 1 0 2872 0 1 4170
box -8 -3 32 105
use FILL  FILL_1070
timestamp 1677622389
transform 1 0 2896 0 1 4170
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1677622389
transform 1 0 2904 0 1 4170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1677622389
transform 1 0 2912 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1677622389
transform -1 0 2952 0 1 4170
box -8 -3 34 105
use FILL  FILL_1075
timestamp 1677622389
transform 1 0 2952 0 1 4170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1677622389
transform 1 0 2960 0 1 4170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1677622389
transform 1 0 2968 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_33
timestamp 1677622389
transform -1 0 3008 0 1 4170
box -8 -3 34 105
use FILL  FILL_1078
timestamp 1677622389
transform 1 0 3008 0 1 4170
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1677622389
transform 1 0 3016 0 1 4170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1677622389
transform 1 0 3024 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_53
timestamp 1677622389
transform 1 0 3032 0 1 4170
box -8 -3 46 105
use FILL  FILL_1090
timestamp 1677622389
transform 1 0 3072 0 1 4170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1677622389
transform 1 0 3080 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_100
timestamp 1677622389
transform -1 0 3104 0 1 4170
box -9 -3 26 105
use M3_M2  M3_M2_977
timestamp 1677622389
transform 1 0 3188 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_88
timestamp 1677622389
transform -1 0 3200 0 1 4170
box -8 -3 104 105
use M3_M2  M3_M2_978
timestamp 1677622389
transform 1 0 3220 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_101
timestamp 1677622389
transform 1 0 3200 0 1 4170
box -9 -3 26 105
use FILL  FILL_1098
timestamp 1677622389
transform 1 0 3216 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_54
timestamp 1677622389
transform -1 0 3264 0 1 4170
box -8 -3 46 105
use FILL  FILL_1099
timestamp 1677622389
transform 1 0 3264 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_979
timestamp 1677622389
transform 1 0 3284 0 1 4175
box -3 -3 3 3
use FILL  FILL_1100
timestamp 1677622389
transform 1 0 3272 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_980
timestamp 1677622389
transform 1 0 3356 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_89
timestamp 1677622389
transform -1 0 3376 0 1 4170
box -8 -3 104 105
use FILL  FILL_1101
timestamp 1677622389
transform 1 0 3376 0 1 4170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1677622389
transform 1 0 3384 0 1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1677622389
transform -1 0 3424 0 1 4170
box -8 -3 40 105
use FILL  FILL_1103
timestamp 1677622389
transform 1 0 3424 0 1 4170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1677622389
transform 1 0 3432 0 1 4170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1677622389
transform 1 0 3440 0 1 4170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1677622389
transform 1 0 3448 0 1 4170
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1677622389
transform 1 0 3456 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_57
timestamp 1677622389
transform 1 0 3464 0 1 4170
box -8 -3 46 105
use FILL  FILL_1108
timestamp 1677622389
transform 1 0 3504 0 1 4170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1677622389
transform 1 0 3512 0 1 4170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1677622389
transform 1 0 3520 0 1 4170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1677622389
transform 1 0 3528 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_58
timestamp 1677622389
transform -1 0 3576 0 1 4170
box -8 -3 46 105
use FILL  FILL_1112
timestamp 1677622389
transform 1 0 3576 0 1 4170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1677622389
transform 1 0 3584 0 1 4170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1677622389
transform 1 0 3592 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_57
timestamp 1677622389
transform 1 0 3600 0 1 4170
box -8 -3 46 105
use FILL  FILL_1140
timestamp 1677622389
transform 1 0 3640 0 1 4170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1677622389
transform 1 0 3648 0 1 4170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1677622389
transform 1 0 3656 0 1 4170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1677622389
transform 1 0 3664 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_103
timestamp 1677622389
transform -1 0 3688 0 1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1677622389
transform -1 0 3784 0 1 4170
box -8 -3 104 105
use FILL  FILL_1144
timestamp 1677622389
transform 1 0 3784 0 1 4170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1677622389
transform 1 0 3792 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_59
timestamp 1677622389
transform 1 0 3800 0 1 4170
box -8 -3 46 105
use M3_M2  M3_M2_981
timestamp 1677622389
transform 1 0 3852 0 1 4175
box -3 -3 3 3
use FILL  FILL_1154
timestamp 1677622389
transform 1 0 3840 0 1 4170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1677622389
transform 1 0 3848 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_982
timestamp 1677622389
transform 1 0 3892 0 1 4175
box -3 -3 3 3
use OAI22X1  OAI22X1_58
timestamp 1677622389
transform -1 0 3896 0 1 4170
box -8 -3 46 105
use FILL  FILL_1156
timestamp 1677622389
transform 1 0 3896 0 1 4170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1677622389
transform 1 0 3904 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_105
timestamp 1677622389
transform -1 0 3928 0 1 4170
box -9 -3 26 105
use FILL  FILL_1158
timestamp 1677622389
transform 1 0 3928 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_983
timestamp 1677622389
transform 1 0 3948 0 1 4175
box -3 -3 3 3
use FILL  FILL_1168
timestamp 1677622389
transform 1 0 3936 0 1 4170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1677622389
transform 1 0 3944 0 1 4170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1677622389
transform 1 0 3952 0 1 4170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1677622389
transform 1 0 3960 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_106
timestamp 1677622389
transform -1 0 3984 0 1 4170
box -9 -3 26 105
use FILL  FILL_1172
timestamp 1677622389
transform 1 0 3984 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_984
timestamp 1677622389
transform 1 0 4004 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1677622389
transform 1 0 4076 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1677622389
transform 1 0 4092 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_93
timestamp 1677622389
transform 1 0 3992 0 1 4170
box -8 -3 104 105
use OAI22X1  OAI22X1_60
timestamp 1677622389
transform 1 0 4088 0 1 4170
box -8 -3 46 105
use FILL  FILL_1180
timestamp 1677622389
transform 1 0 4128 0 1 4170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1677622389
transform 1 0 4136 0 1 4170
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1677622389
transform 1 0 4144 0 1 4170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1677622389
transform 1 0 4152 0 1 4170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1677622389
transform 1 0 4160 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_107
timestamp 1677622389
transform 1 0 4168 0 1 4170
box -9 -3 26 105
use FILL  FILL_1189
timestamp 1677622389
transform 1 0 4184 0 1 4170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1677622389
transform 1 0 4192 0 1 4170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1677622389
transform 1 0 4200 0 1 4170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1677622389
transform 1 0 4208 0 1 4170
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1677622389
transform 1 0 4216 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_987
timestamp 1677622389
transform 1 0 4268 0 1 4175
box -3 -3 3 3
use AOI22X1  AOI22X1_60
timestamp 1677622389
transform -1 0 4264 0 1 4170
box -8 -3 46 105
use FILL  FILL_1199
timestamp 1677622389
transform 1 0 4264 0 1 4170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1677622389
transform 1 0 4272 0 1 4170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1677622389
transform 1 0 4280 0 1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1677622389
transform -1 0 4320 0 1 4170
box -8 -3 40 105
use FILL  FILL_1210
timestamp 1677622389
transform 1 0 4320 0 1 4170
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1677622389
transform 1 0 4328 0 1 4170
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1677622389
transform 1 0 4336 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1677622389
transform 1 0 4344 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_109
timestamp 1677622389
transform 1 0 4440 0 1 4170
box -9 -3 26 105
use M3_M2  M3_M2_988
timestamp 1677622389
transform 1 0 4484 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_110
timestamp 1677622389
transform 1 0 4456 0 1 4170
box -9 -3 26 105
use FILL  FILL_1223
timestamp 1677622389
transform 1 0 4472 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_62
timestamp 1677622389
transform 1 0 4480 0 1 4170
box -8 -3 46 105
use FILL  FILL_1225
timestamp 1677622389
transform 1 0 4520 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_61
timestamp 1677622389
transform -1 0 4568 0 1 4170
box -8 -3 46 105
use FILL  FILL_1226
timestamp 1677622389
transform 1 0 4568 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1677622389
transform -1 0 4592 0 1 4170
box -9 -3 26 105
use FILL  FILL_1227
timestamp 1677622389
transform 1 0 4592 0 1 4170
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1677622389
transform 1 0 4600 0 1 4170
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1677622389
transform 1 0 4608 0 1 4170
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1677622389
transform 1 0 4616 0 1 4170
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1677622389
transform 1 0 4624 0 1 4170
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1677622389
transform 1 0 4632 0 1 4170
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1677622389
transform 1 0 4640 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_989
timestamp 1677622389
transform 1 0 4660 0 1 4175
box -3 -3 3 3
use FILL  FILL_1241
timestamp 1677622389
transform 1 0 4648 0 1 4170
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1677622389
transform 1 0 4656 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_63
timestamp 1677622389
transform 1 0 4664 0 1 4170
box -8 -3 46 105
use FILL  FILL_1243
timestamp 1677622389
transform 1 0 4704 0 1 4170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1677622389
transform 1 0 4712 0 1 4170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1677622389
transform 1 0 4720 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_115
timestamp 1677622389
transform 1 0 4728 0 1 4170
box -9 -3 26 105
use FILL  FILL_1252
timestamp 1677622389
transform 1 0 4744 0 1 4170
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1677622389
transform 1 0 4752 0 1 4170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1677622389
transform 1 0 4760 0 1 4170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1677622389
transform 1 0 4768 0 1 4170
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1677622389
transform 1 0 4776 0 1 4170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1677622389
transform 1 0 4784 0 1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_11
timestamp 1677622389
transform 1 0 4819 0 1 4170
box -10 -3 10 3
use M2_M1  M2_M1_1257
timestamp 1677622389
transform 1 0 116 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1677622389
transform 1 0 156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1677622389
transform 1 0 164 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1049
timestamp 1677622389
transform 1 0 156 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1677622389
transform 1 0 196 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1167
timestamp 1677622389
transform 1 0 196 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1677622389
transform 1 0 164 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1677622389
transform 1 0 172 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1677622389
transform 1 0 180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1677622389
transform 1 0 196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1677622389
transform 1 0 204 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1677622389
transform 1 0 164 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1677622389
transform 1 0 212 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1677622389
transform 1 0 204 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1677622389
transform 1 0 204 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1677622389
transform 1 0 228 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1168
timestamp 1677622389
transform 1 0 228 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1677622389
transform 1 0 244 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1052
timestamp 1677622389
transform 1 0 244 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1262
timestamp 1677622389
transform 1 0 292 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1677622389
transform 1 0 324 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1677622389
transform 1 0 332 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1085
timestamp 1677622389
transform 1 0 292 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1677622389
transform 1 0 332 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1677622389
transform 1 0 284 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1677622389
transform 1 0 348 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1677622389
transform 1 0 396 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1677622389
transform 1 0 468 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1677622389
transform 1 0 476 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1677622389
transform 1 0 500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1677622389
transform 1 0 508 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1677622389
transform 1 0 460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1677622389
transform 1 0 468 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1677622389
transform 1 0 476 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1268
timestamp 1677622389
transform 1 0 484 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1677622389
transform 1 0 500 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1054
timestamp 1677622389
transform 1 0 508 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1677622389
transform 1 0 500 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1677622389
transform 1 0 500 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1677622389
transform 1 0 516 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1175
timestamp 1677622389
transform 1 0 556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1677622389
transform 1 0 564 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1677622389
transform 1 0 532 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1677622389
transform 1 0 548 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1677622389
transform 1 0 564 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1140
timestamp 1677622389
transform 1 0 524 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1677622389
transform 1 0 564 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1677622389
transform 1 0 556 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1677622389
transform 1 0 556 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1677622389
transform 1 0 596 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1677622389
transform 1 0 620 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1177
timestamp 1677622389
transform 1 0 724 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1677622389
transform 1 0 636 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1677622389
transform 1 0 644 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1677622389
transform 1 0 676 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1091
timestamp 1677622389
transform 1 0 636 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1677622389
transform 1 0 676 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1677622389
transform 1 0 644 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1677622389
transform 1 0 772 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1276
timestamp 1677622389
transform 1 0 772 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1677622389
transform 1 0 788 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1677622389
transform 1 0 804 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1677622389
transform 1 0 820 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1677622389
transform 1 0 812 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1123
timestamp 1677622389
transform 1 0 788 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1278
timestamp 1677622389
transform 1 0 868 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1677622389
transform 1 0 892 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1056
timestamp 1677622389
transform 1 0 916 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1181
timestamp 1677622389
transform 1 0 940 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1677622389
transform 1 0 948 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1677622389
transform 1 0 964 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1677622389
transform 1 0 948 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1280
timestamp 1677622389
transform 1 0 956 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1058
timestamp 1677622389
transform 1 0 964 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1184
timestamp 1677622389
transform 1 0 980 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1034
timestamp 1677622389
transform 1 0 1020 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1281
timestamp 1677622389
transform 1 0 1012 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1677622389
transform 1 0 1020 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1093
timestamp 1677622389
transform 1 0 1012 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1677622389
transform 1 0 1036 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1185
timestamp 1677622389
transform 1 0 1044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1677622389
transform 1 0 1052 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1059
timestamp 1677622389
transform 1 0 1052 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1677622389
transform 1 0 1052 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1677622389
transform 1 0 1076 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1677622389
transform 1 0 1076 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1124
timestamp 1677622389
transform 1 0 1076 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1283
timestamp 1677622389
transform 1 0 1100 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1677622389
transform 1 0 1124 0 1 4145
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1677622389
transform 1 0 1124 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1187
timestamp 1677622389
transform 1 0 1156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1677622389
transform 1 0 1164 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1677622389
transform 1 0 1148 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1364
timestamp 1677622389
transform 1 0 1148 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1677622389
transform 1 0 1172 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1677622389
transform 1 0 1188 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1677622389
transform 1 0 1284 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1677622389
transform 1 0 1252 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1150
timestamp 1677622389
transform 1 0 1284 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1190
timestamp 1677622389
transform 1 0 1300 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1677622389
transform 1 0 1300 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1677622389
transform 1 0 1316 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1677622389
transform 1 0 1308 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1677622389
transform 1 0 1332 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1287
timestamp 1677622389
transform 1 0 1356 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1677622389
transform 1 0 1388 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1677622389
transform 1 0 1396 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1677622389
transform 1 0 1412 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1126
timestamp 1677622389
transform 1 0 1388 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1288
timestamp 1677622389
transform 1 0 1404 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1677622389
transform 1 0 1412 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1677622389
transform 1 0 1436 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1062
timestamp 1677622389
transform 1 0 1436 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1289
timestamp 1677622389
transform 1 0 1444 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1677622389
transform 1 0 1452 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1677622389
transform 1 0 1540 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1677622389
transform 1 0 1500 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1097
timestamp 1677622389
transform 1 0 1500 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1196
timestamp 1677622389
transform 1 0 1564 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1142
timestamp 1677622389
transform 1 0 1556 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1677622389
transform 1 0 1612 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1197
timestamp 1677622389
transform 1 0 1620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1677622389
transform 1 0 1636 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1677622389
transform 1 0 1612 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1677622389
transform 1 0 1628 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1037
timestamp 1677622389
transform 1 0 1644 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1677622389
transform 1 0 1612 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1677622389
transform 1 0 1636 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1677622389
transform 1 0 1660 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1677622389
transform 1 0 1676 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1294
timestamp 1677622389
transform 1 0 1668 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1677622389
transform 1 0 1692 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1199
timestamp 1677622389
transform 1 0 1708 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1129
timestamp 1677622389
transform 1 0 1732 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1677622389
transform 1 0 1772 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1677622389
transform 1 0 1788 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1677622389
transform 1 0 1756 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1677622389
transform 1 0 1764 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1063
timestamp 1677622389
transform 1 0 1772 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1297
timestamp 1677622389
transform 1 0 1780 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1064
timestamp 1677622389
transform 1 0 1788 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1298
timestamp 1677622389
transform 1 0 1804 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1677622389
transform 1 0 1812 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1130
timestamp 1677622389
transform 1 0 1828 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1677622389
transform 1 0 1836 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1299
timestamp 1677622389
transform 1 0 1860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1677622389
transform 1 0 1868 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1098
timestamp 1677622389
transform 1 0 1868 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1203
timestamp 1677622389
transform 1 0 1884 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1065
timestamp 1677622389
transform 1 0 1884 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1301
timestamp 1677622389
transform 1 0 1916 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_990
timestamp 1677622389
transform 1 0 1940 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1677622389
transform 1 0 1940 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1677622389
transform 1 0 1940 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1204
timestamp 1677622389
transform 1 0 1940 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1677622389
transform 1 0 1948 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_991
timestamp 1677622389
transform 1 0 2012 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1677622389
transform 1 0 2108 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1677622389
transform 1 0 2108 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1677622389
transform 1 0 2028 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1677622389
transform 1 0 2084 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1099
timestamp 1677622389
transform 1 0 2060 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1305
timestamp 1677622389
transform 1 0 2124 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1677622389
transform 1 0 2140 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1677622389
transform 1 0 2132 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1677622389
transform 1 0 2124 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1677622389
transform 1 0 2188 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1677622389
transform 1 0 2188 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1677622389
transform 1 0 2180 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1066
timestamp 1677622389
transform 1 0 2188 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1677622389
transform 1 0 2204 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1067
timestamp 1677622389
transform 1 0 2204 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1307
timestamp 1677622389
transform 1 0 2212 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1068
timestamp 1677622389
transform 1 0 2220 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1677622389
transform 1 0 2212 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1677622389
transform 1 0 2260 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1677622389
transform 1 0 2308 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1677622389
transform 1 0 2244 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1677622389
transform 1 0 2340 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1677622389
transform 1 0 2340 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1677622389
transform 1 0 2252 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1677622389
transform 1 0 2260 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1677622389
transform 1 0 2292 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1069
timestamp 1677622389
transform 1 0 2340 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1677622389
transform 1 0 2252 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1677622389
transform 1 0 2292 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1677622389
transform 1 0 2316 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1677622389
transform 1 0 2364 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1210
timestamp 1677622389
transform 1 0 2364 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_995
timestamp 1677622389
transform 1 0 2412 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1677622389
transform 1 0 2404 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1211
timestamp 1677622389
transform 1 0 2412 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1677622389
transform 1 0 2428 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1677622389
transform 1 0 2404 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1021
timestamp 1677622389
transform 1 0 2452 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1677622389
transform 1 0 2444 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1677622389
transform 1 0 2468 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1677622389
transform 1 0 2532 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1677622389
transform 1 0 2444 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1677622389
transform 1 0 2452 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1677622389
transform 1 0 2460 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1314
timestamp 1677622389
transform 1 0 2508 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1677622389
transform 1 0 2548 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1677622389
transform 1 0 2556 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1103
timestamp 1677622389
transform 1 0 2508 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1677622389
transform 1 0 2548 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1677622389
transform 1 0 2556 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1677622389
transform 1 0 2620 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1214
timestamp 1677622389
transform 1 0 2596 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1677622389
transform 1 0 2604 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1677622389
transform 1 0 2620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1677622389
transform 1 0 2628 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1677622389
transform 1 0 2612 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1677622389
transform 1 0 2620 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1677622389
transform 1 0 2604 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1677622389
transform 1 0 2628 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1677622389
transform 1 0 2652 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1677622389
transform 1 0 2668 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1677622389
transform 1 0 2684 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1677622389
transform 1 0 2692 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1677622389
transform 1 0 2652 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1677622389
transform 1 0 2660 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1677622389
transform 1 0 2676 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1072
timestamp 1677622389
transform 1 0 2684 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1677622389
transform 1 0 2668 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1677622389
transform 1 0 2700 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1321
timestamp 1677622389
transform 1 0 2700 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1004
timestamp 1677622389
transform 1 0 2796 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1221
timestamp 1677622389
transform 1 0 2732 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1677622389
transform 1 0 2716 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1677622389
transform 1 0 2756 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1073
timestamp 1677622389
transform 1 0 2804 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1324
timestamp 1677622389
transform 1 0 2812 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1677622389
transform 1 0 2716 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1677622389
transform 1 0 2756 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1677622389
transform 1 0 2828 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1164
timestamp 1677622389
transform 1 0 2828 0 1 4145
box -2 -2 2 2
use M3_M2  M3_M2_997
timestamp 1677622389
transform 1 0 2844 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1677622389
transform 1 0 2844 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1222
timestamp 1677622389
transform 1 0 2836 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1677622389
transform 1 0 2844 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1677622389
transform 1 0 2836 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1677622389
transform 1 0 2868 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1325
timestamp 1677622389
transform 1 0 2860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1677622389
transform 1 0 2868 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1677622389
transform 1 0 2892 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1677622389
transform 1 0 2924 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1677622389
transform 1 0 2940 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1677622389
transform 1 0 2964 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1677622389
transform 1 0 2980 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1677622389
transform 1 0 3004 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1225
timestamp 1677622389
transform 1 0 3020 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1074
timestamp 1677622389
transform 1 0 3020 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1677622389
transform 1 0 3020 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1329
timestamp 1677622389
transform 1 0 3044 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1677622389
transform 1 0 3100 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1677622389
transform 1 0 3116 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1144
timestamp 1677622389
transform 1 0 3108 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1677622389
transform 1 0 3156 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1228
timestamp 1677622389
transform 1 0 3156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1677622389
transform 1 0 3148 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1075
timestamp 1677622389
transform 1 0 3156 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1331
timestamp 1677622389
transform 1 0 3164 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1677622389
transform 1 0 3180 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1677622389
transform 1 0 3204 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1005
timestamp 1677622389
transform 1 0 3220 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1677622389
transform 1 0 3244 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1231
timestamp 1677622389
transform 1 0 3220 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1677622389
transform 1 0 3244 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1006
timestamp 1677622389
transform 1 0 3364 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1232
timestamp 1677622389
transform 1 0 3356 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1076
timestamp 1677622389
transform 1 0 3340 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1333
timestamp 1677622389
transform 1 0 3348 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1677622389
transform 1 0 3396 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1133
timestamp 1677622389
transform 1 0 3396 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1677622389
transform 1 0 3436 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1335
timestamp 1677622389
transform 1 0 3428 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1677622389
transform 1 0 3412 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1026
timestamp 1677622389
transform 1 0 3452 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1233
timestamp 1677622389
transform 1 0 3452 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1677622389
transform 1 0 3444 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1677622389
transform 1 0 3420 0 1 4105
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1677622389
transform 1 0 3420 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1336
timestamp 1677622389
transform 1 0 3468 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1134
timestamp 1677622389
transform 1 0 3468 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1677622389
transform 1 0 3500 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1677622389
transform 1 0 3484 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1677622389
transform 1 0 3508 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1234
timestamp 1677622389
transform 1 0 3500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1677622389
transform 1 0 3484 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1677622389
transform 1 0 3524 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1677622389
transform 1 0 3532 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1677622389
transform 1 0 3508 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1077
timestamp 1677622389
transform 1 0 3532 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1677622389
transform 1 0 3524 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1677622389
transform 1 0 3508 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1677622389
transform 1 0 3580 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1677622389
transform 1 0 3572 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1237
timestamp 1677622389
transform 1 0 3572 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1677622389
transform 1 0 3588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1677622389
transform 1 0 3564 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1677622389
transform 1 0 3580 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1677622389
transform 1 0 3596 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1677622389
transform 1 0 3644 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1239
timestamp 1677622389
transform 1 0 3620 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1047
timestamp 1677622389
transform 1 0 3652 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1677622389
transform 1 0 3644 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1677622389
transform 1 0 3620 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1677622389
transform 1 0 3740 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1342
timestamp 1677622389
transform 1 0 3740 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1677622389
transform 1 0 3748 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1677622389
transform 1 0 3748 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1240
timestamp 1677622389
transform 1 0 3772 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1677622389
transform 1 0 3804 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1137
timestamp 1677622389
transform 1 0 3804 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1241
timestamp 1677622389
transform 1 0 3844 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1677622389
transform 1 0 3852 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1078
timestamp 1677622389
transform 1 0 3852 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1677622389
transform 1 0 3892 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1243
timestamp 1677622389
transform 1 0 3892 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1677622389
transform 1 0 3876 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1677622389
transform 1 0 3900 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1010
timestamp 1677622389
transform 1 0 3932 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1677622389
transform 1 0 3932 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1011
timestamp 1677622389
transform 1 0 3980 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1677622389
transform 1 0 3972 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1245
timestamp 1677622389
transform 1 0 3948 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1677622389
transform 1 0 3972 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1677622389
transform 1 0 4028 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1032
timestamp 1677622389
transform 1 0 4084 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1677622389
transform 1 0 4124 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1677622389
transform 1 0 4132 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1677622389
transform 1 0 4092 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1677622389
transform 1 0 4108 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1677622389
transform 1 0 4124 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1677622389
transform 1 0 4132 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1079
timestamp 1677622389
transform 1 0 4092 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1349
timestamp 1677622389
transform 1 0 4100 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1677622389
transform 1 0 4116 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1145
timestamp 1677622389
transform 1 0 4092 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1677622389
transform 1 0 4132 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1013
timestamp 1677622389
transform 1 0 4148 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1352
timestamp 1677622389
transform 1 0 4204 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1138
timestamp 1677622389
transform 1 0 4228 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1677622389
transform 1 0 4268 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1677622389
transform 1 0 4300 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1250
timestamp 1677622389
transform 1 0 4356 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1677622389
transform 1 0 4380 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1114
timestamp 1677622389
transform 1 0 4380 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1677622389
transform 1 0 4468 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1677622389
transform 1 0 4484 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1000
timestamp 1677622389
transform 1 0 4500 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1677622389
transform 1 0 4508 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1115
timestamp 1677622389
transform 1 0 4508 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1371
timestamp 1677622389
transform 1 0 4516 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1677622389
transform 1 0 4500 0 1 4105
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1677622389
transform 1 0 4516 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1356
timestamp 1677622389
transform 1 0 4532 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1146
timestamp 1677622389
transform 1 0 4532 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1251
timestamp 1677622389
transform 1 0 4556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1677622389
transform 1 0 4572 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1677622389
transform 1 0 4588 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1116
timestamp 1677622389
transform 1 0 4572 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1677622389
transform 1 0 4604 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1677622389
transform 1 0 4612 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1252
timestamp 1677622389
transform 1 0 4628 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1081
timestamp 1677622389
transform 1 0 4628 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1359
timestamp 1677622389
transform 1 0 4636 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1117
timestamp 1677622389
transform 1 0 4636 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1253
timestamp 1677622389
transform 1 0 4652 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1677622389
transform 1 0 4660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1677622389
transform 1 0 4676 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1048
timestamp 1677622389
transform 1 0 4684 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1256
timestamp 1677622389
transform 1 0 4692 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1677622389
transform 1 0 4652 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1677622389
transform 1 0 4668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1677622389
transform 1 0 4684 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1118
timestamp 1677622389
transform 1 0 4684 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1677622389
transform 1 0 4652 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1677622389
transform 1 0 4788 0 1 4125
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_12
timestamp 1677622389
transform 1 0 24 0 1 4070
box -10 -3 10 3
use FILL  FILL_808
timestamp 1677622389
transform 1 0 72 0 -1 4170
box -8 -3 16 105
use FILL  FILL_809
timestamp 1677622389
transform 1 0 80 0 -1 4170
box -8 -3 16 105
use FILL  FILL_810
timestamp 1677622389
transform 1 0 88 0 -1 4170
box -8 -3 16 105
use FILL  FILL_811
timestamp 1677622389
transform 1 0 96 0 -1 4170
box -8 -3 16 105
use FILL  FILL_812
timestamp 1677622389
transform 1 0 104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_813
timestamp 1677622389
transform 1 0 112 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_77
timestamp 1677622389
transform -1 0 136 0 -1 4170
box -9 -3 26 105
use FILL  FILL_814
timestamp 1677622389
transform 1 0 136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_815
timestamp 1677622389
transform 1 0 144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_816
timestamp 1677622389
transform 1 0 152 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_43
timestamp 1677622389
transform -1 0 200 0 -1 4170
box -8 -3 46 105
use FILL  FILL_817
timestamp 1677622389
transform 1 0 200 0 -1 4170
box -8 -3 16 105
use FILL  FILL_824
timestamp 1677622389
transform 1 0 208 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_78
timestamp 1677622389
transform -1 0 232 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1677622389
transform 1 0 232 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_79
timestamp 1677622389
transform -1 0 344 0 -1 4170
box -9 -3 26 105
use FILL  FILL_825
timestamp 1677622389
transform 1 0 344 0 -1 4170
box -8 -3 16 105
use FILL  FILL_827
timestamp 1677622389
transform 1 0 352 0 -1 4170
box -8 -3 16 105
use FILL  FILL_828
timestamp 1677622389
transform 1 0 360 0 -1 4170
box -8 -3 16 105
use FILL  FILL_829
timestamp 1677622389
transform 1 0 368 0 -1 4170
box -8 -3 16 105
use FILL  FILL_830
timestamp 1677622389
transform 1 0 376 0 -1 4170
box -8 -3 16 105
use FILL  FILL_831
timestamp 1677622389
transform 1 0 384 0 -1 4170
box -8 -3 16 105
use FILL  FILL_832
timestamp 1677622389
transform 1 0 392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_833
timestamp 1677622389
transform 1 0 400 0 -1 4170
box -8 -3 16 105
use FILL  FILL_834
timestamp 1677622389
transform 1 0 408 0 -1 4170
box -8 -3 16 105
use FILL  FILL_835
timestamp 1677622389
transform 1 0 416 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_80
timestamp 1677622389
transform -1 0 440 0 -1 4170
box -9 -3 26 105
use FILL  FILL_836
timestamp 1677622389
transform 1 0 440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_837
timestamp 1677622389
transform 1 0 448 0 -1 4170
box -8 -3 16 105
use FILL  FILL_839
timestamp 1677622389
transform 1 0 456 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_44
timestamp 1677622389
transform 1 0 464 0 -1 4170
box -8 -3 46 105
use FILL  FILL_846
timestamp 1677622389
transform 1 0 504 0 -1 4170
box -8 -3 16 105
use FILL  FILL_848
timestamp 1677622389
transform 1 0 512 0 -1 4170
box -8 -3 16 105
use FILL  FILL_850
timestamp 1677622389
transform 1 0 520 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_46
timestamp 1677622389
transform 1 0 528 0 -1 4170
box -8 -3 46 105
use FILL  FILL_852
timestamp 1677622389
transform 1 0 568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1677622389
transform 1 0 576 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_82
timestamp 1677622389
transform 1 0 584 0 -1 4170
box -9 -3 26 105
use FILL  FILL_856
timestamp 1677622389
transform 1 0 600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1677622389
transform 1 0 608 0 -1 4170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1677622389
transform 1 0 616 0 -1 4170
box -8 -3 16 105
use FILL  FILL_863
timestamp 1677622389
transform 1 0 624 0 -1 4170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1677622389
transform 1 0 632 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1677622389
transform -1 0 736 0 -1 4170
box -8 -3 104 105
use FILL  FILL_865
timestamp 1677622389
transform 1 0 736 0 -1 4170
box -8 -3 16 105
use FILL  FILL_866
timestamp 1677622389
transform 1 0 744 0 -1 4170
box -8 -3 16 105
use FILL  FILL_868
timestamp 1677622389
transform 1 0 752 0 -1 4170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1677622389
transform 1 0 760 0 -1 4170
box -8 -3 16 105
use FILL  FILL_874
timestamp 1677622389
transform 1 0 768 0 -1 4170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1677622389
transform 1 0 776 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_44
timestamp 1677622389
transform 1 0 784 0 -1 4170
box -8 -3 46 105
use FILL  FILL_876
timestamp 1677622389
transform 1 0 824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1677622389
transform 1 0 832 0 -1 4170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1677622389
transform 1 0 840 0 -1 4170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1677622389
transform 1 0 848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1677622389
transform 1 0 856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1677622389
transform 1 0 864 0 -1 4170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1677622389
transform 1 0 872 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_84
timestamp 1677622389
transform -1 0 896 0 -1 4170
box -9 -3 26 105
use FILL  FILL_883
timestamp 1677622389
transform 1 0 896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_884
timestamp 1677622389
transform 1 0 904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1677622389
transform 1 0 912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1677622389
transform 1 0 920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1677622389
transform 1 0 928 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_47
timestamp 1677622389
transform 1 0 936 0 -1 4170
box -8 -3 46 105
use FILL  FILL_892
timestamp 1677622389
transform 1 0 976 0 -1 4170
box -8 -3 16 105
use FILL  FILL_894
timestamp 1677622389
transform 1 0 984 0 -1 4170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1677622389
transform 1 0 992 0 -1 4170
box -8 -3 16 105
use FILL  FILL_898
timestamp 1677622389
transform 1 0 1000 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_24
timestamp 1677622389
transform 1 0 1008 0 -1 4170
box -8 -3 34 105
use FILL  FILL_901
timestamp 1677622389
transform 1 0 1040 0 -1 4170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1677622389
transform 1 0 1048 0 -1 4170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1677622389
transform 1 0 1056 0 -1 4170
box -8 -3 16 105
use FILL  FILL_921
timestamp 1677622389
transform 1 0 1064 0 -1 4170
box -8 -3 16 105
use FILL  FILL_922
timestamp 1677622389
transform 1 0 1072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1677622389
transform 1 0 1080 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_27
timestamp 1677622389
transform 1 0 1088 0 -1 4170
box -8 -3 34 105
use FILL  FILL_924
timestamp 1677622389
transform 1 0 1120 0 -1 4170
box -8 -3 16 105
use FILL  FILL_925
timestamp 1677622389
transform 1 0 1128 0 -1 4170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1677622389
transform 1 0 1136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1677622389
transform 1 0 1144 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1677622389
transform 1 0 1152 0 -1 4170
box -8 -3 32 105
use FILL  FILL_928
timestamp 1677622389
transform 1 0 1176 0 -1 4170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1677622389
transform 1 0 1184 0 -1 4170
box -8 -3 16 105
use FILL  FILL_930
timestamp 1677622389
transform 1 0 1192 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1159
timestamp 1677622389
transform 1 0 1284 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_76
timestamp 1677622389
transform -1 0 1296 0 -1 4170
box -8 -3 104 105
use FILL  FILL_931
timestamp 1677622389
transform 1 0 1296 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1160
timestamp 1677622389
transform 1 0 1316 0 1 4075
box -3 -3 3 3
use FILL  FILL_933
timestamp 1677622389
transform 1 0 1304 0 -1 4170
box -8 -3 16 105
use FILL  FILL_935
timestamp 1677622389
transform 1 0 1312 0 -1 4170
box -8 -3 16 105
use FILL  FILL_938
timestamp 1677622389
transform 1 0 1320 0 -1 4170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1677622389
transform 1 0 1328 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_29
timestamp 1677622389
transform -1 0 1368 0 -1 4170
box -8 -3 34 105
use FILL  FILL_940
timestamp 1677622389
transform 1 0 1368 0 -1 4170
box -8 -3 16 105
use FILL  FILL_941
timestamp 1677622389
transform 1 0 1376 0 -1 4170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1677622389
transform 1 0 1384 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_47
timestamp 1677622389
transform -1 0 1432 0 -1 4170
box -8 -3 46 105
use FILL  FILL_952
timestamp 1677622389
transform 1 0 1432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1677622389
transform 1 0 1440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1677622389
transform 1 0 1448 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1677622389
transform -1 0 1552 0 -1 4170
box -8 -3 104 105
use FILL  FILL_955
timestamp 1677622389
transform 1 0 1552 0 -1 4170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1677622389
transform 1 0 1560 0 -1 4170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1677622389
transform 1 0 1568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1677622389
transform 1 0 1576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1677622389
transform 1 0 1584 0 -1 4170
box -8 -3 16 105
use FILL  FILL_964
timestamp 1677622389
transform 1 0 1592 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_48
timestamp 1677622389
transform -1 0 1640 0 -1 4170
box -8 -3 46 105
use FILL  FILL_965
timestamp 1677622389
transform 1 0 1640 0 -1 4170
box -8 -3 16 105
use FILL  FILL_966
timestamp 1677622389
transform 1 0 1648 0 -1 4170
box -8 -3 16 105
use FILL  FILL_967
timestamp 1677622389
transform 1 0 1656 0 -1 4170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1677622389
transform 1 0 1664 0 -1 4170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1677622389
transform 1 0 1672 0 -1 4170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1677622389
transform 1 0 1680 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_90
timestamp 1677622389
transform -1 0 1704 0 -1 4170
box -9 -3 26 105
use FILL  FILL_971
timestamp 1677622389
transform 1 0 1704 0 -1 4170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1677622389
transform 1 0 1712 0 -1 4170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1677622389
transform 1 0 1720 0 -1 4170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1677622389
transform 1 0 1728 0 -1 4170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1677622389
transform 1 0 1736 0 -1 4170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1677622389
transform 1 0 1744 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1161
timestamp 1677622389
transform 1 0 1764 0 1 4075
box -3 -3 3 3
use FILL  FILL_983
timestamp 1677622389
transform 1 0 1752 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1677622389
transform 1 0 1760 0 -1 4170
box -8 -3 46 105
use M3_M2  M3_M2_1162
timestamp 1677622389
transform 1 0 1812 0 1 4075
box -3 -3 3 3
use FILL  FILL_984
timestamp 1677622389
transform 1 0 1800 0 -1 4170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1677622389
transform 1 0 1808 0 -1 4170
box -8 -3 16 105
use FILL  FILL_986
timestamp 1677622389
transform 1 0 1816 0 -1 4170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1677622389
transform 1 0 1824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1677622389
transform 1 0 1832 0 -1 4170
box -8 -3 16 105
use FILL  FILL_989
timestamp 1677622389
transform 1 0 1840 0 -1 4170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1677622389
transform 1 0 1848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1677622389
transform 1 0 1856 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1163
timestamp 1677622389
transform 1 0 1876 0 1 4075
box -3 -3 3 3
use INVX2  INVX2_92
timestamp 1677622389
transform 1 0 1864 0 -1 4170
box -9 -3 26 105
use FILL  FILL_992
timestamp 1677622389
transform 1 0 1880 0 -1 4170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1677622389
transform 1 0 1888 0 -1 4170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1677622389
transform 1 0 1896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1677622389
transform 1 0 1904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1677622389
transform 1 0 1912 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_50
timestamp 1677622389
transform 1 0 1920 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1002
timestamp 1677622389
transform 1 0 1960 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1677622389
transform 1 0 1968 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1677622389
transform 1 0 1976 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1677622389
transform 1 0 1984 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1677622389
transform 1 0 1992 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1677622389
transform 1 0 2000 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1677622389
transform 1 0 2008 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1677622389
transform 1 0 2016 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1164
timestamp 1677622389
transform 1 0 2100 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_81
timestamp 1677622389
transform -1 0 2120 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1018
timestamp 1677622389
transform 1 0 2120 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1677622389
transform 1 0 2128 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1677622389
transform 1 0 2136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1677622389
transform 1 0 2144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1677622389
transform 1 0 2152 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1677622389
transform 1 0 2160 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1023
timestamp 1677622389
transform 1 0 2200 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1677622389
transform 1 0 2208 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1677622389
transform 1 0 2216 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1677622389
transform 1 0 2224 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1677622389
transform 1 0 2232 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_96
timestamp 1677622389
transform 1 0 2240 0 -1 4170
box -9 -3 26 105
use M3_M2  M3_M2_1165
timestamp 1677622389
transform 1 0 2340 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_84
timestamp 1677622389
transform -1 0 2352 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1047
timestamp 1677622389
transform 1 0 2352 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1677622389
transform 1 0 2360 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1677622389
transform 1 0 2368 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1166
timestamp 1677622389
transform 1 0 2388 0 1 4075
box -3 -3 3 3
use FILL  FILL_1050
timestamp 1677622389
transform 1 0 2376 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1677622389
transform 1 0 2384 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_52
timestamp 1677622389
transform -1 0 2432 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1052
timestamp 1677622389
transform 1 0 2432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1677622389
transform 1 0 2440 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1167
timestamp 1677622389
transform 1 0 2484 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1677622389
transform 1 0 2532 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_85
timestamp 1677622389
transform -1 0 2544 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_97
timestamp 1677622389
transform -1 0 2560 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1054
timestamp 1677622389
transform 1 0 2560 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1677622389
transform 1 0 2568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1677622389
transform 1 0 2576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1677622389
transform 1 0 2584 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_55
timestamp 1677622389
transform 1 0 2592 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1058
timestamp 1677622389
transform 1 0 2632 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1677622389
transform 1 0 2640 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1677622389
transform 1 0 2648 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_56
timestamp 1677622389
transform 1 0 2656 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1061
timestamp 1677622389
transform 1 0 2696 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_98
timestamp 1677622389
transform 1 0 2704 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1677622389
transform 1 0 2720 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1065
timestamp 1677622389
transform 1 0 2816 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1677622389
transform 1 0 2824 0 -1 4170
box -8 -3 32 105
use FILL  FILL_1067
timestamp 1677622389
transform 1 0 2848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1677622389
transform 1 0 2856 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1677622389
transform 1 0 2864 0 -1 4170
box -8 -3 34 105
use FILL  FILL_1071
timestamp 1677622389
transform 1 0 2896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1677622389
transform 1 0 2904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1677622389
transform 1 0 2912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1677622389
transform 1 0 2920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1677622389
transform 1 0 2928 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1677622389
transform 1 0 2936 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_34
timestamp 1677622389
transform -1 0 2976 0 -1 4170
box -8 -3 34 105
use FILL  FILL_1083
timestamp 1677622389
transform 1 0 2976 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1677622389
transform 1 0 2984 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1677622389
transform 1 0 2992 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1677622389
transform 1 0 3000 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1677622389
transform 1 0 3008 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1677622389
transform 1 0 3016 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_99
timestamp 1677622389
transform -1 0 3040 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1092
timestamp 1677622389
transform 1 0 3040 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1677622389
transform 1 0 3048 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1677622389
transform 1 0 3056 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1677622389
transform 1 0 3064 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1677622389
transform 1 0 3072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1677622389
transform 1 0 3080 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1677622389
transform 1 0 3088 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1677622389
transform 1 0 3096 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1677622389
transform 1 0 3104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1677622389
transform 1 0 3112 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1677622389
transform 1 0 3120 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1677622389
transform 1 0 3128 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_55
timestamp 1677622389
transform 1 0 3136 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1122
timestamp 1677622389
transform 1 0 3176 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1677622389
transform 1 0 3184 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1677622389
transform 1 0 3192 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1677622389
transform 1 0 3200 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1677622389
transform 1 0 3208 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1126
timestamp 1677622389
transform 1 0 3304 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1677622389
transform 1 0 3312 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1677622389
transform 1 0 3320 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1677622389
transform 1 0 3328 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_102
timestamp 1677622389
transform 1 0 3336 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1130
timestamp 1677622389
transform 1 0 3352 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_0
timestamp 1677622389
transform -1 0 3384 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1131
timestamp 1677622389
transform 1 0 3384 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1677622389
transform 1 0 3392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1677622389
transform 1 0 3400 0 -1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1677622389
transform -1 0 3440 0 -1 4170
box -8 -3 40 105
use FILL  FILL_1134
timestamp 1677622389
transform 1 0 3440 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_1
timestamp 1677622389
transform -1 0 3472 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1135
timestamp 1677622389
transform 1 0 3472 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_2
timestamp 1677622389
transform 1 0 3480 0 -1 4170
box -5 -3 28 105
use M3_M2  M3_M2_1169
timestamp 1677622389
transform 1 0 3524 0 1 4075
box -3 -3 3 3
use BUFX2  BUFX2_3
timestamp 1677622389
transform 1 0 3504 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1136
timestamp 1677622389
transform 1 0 3528 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1677622389
transform 1 0 3536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1677622389
transform 1 0 3544 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_56
timestamp 1677622389
transform 1 0 3552 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1139
timestamp 1677622389
transform 1 0 3592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1677622389
transform 1 0 3600 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1677622389
transform 1 0 3608 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1146
timestamp 1677622389
transform 1 0 3704 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1677622389
transform 1 0 3712 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1677622389
transform 1 0 3720 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_104
timestamp 1677622389
transform 1 0 3728 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1149
timestamp 1677622389
transform 1 0 3744 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_4
timestamp 1677622389
transform 1 0 3752 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1150
timestamp 1677622389
transform 1 0 3776 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1677622389
transform 1 0 3784 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1677622389
transform 1 0 3792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1677622389
transform 1 0 3800 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1677622389
transform 1 0 3808 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1677622389
transform 1 0 3816 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_5
timestamp 1677622389
transform 1 0 3824 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1162
timestamp 1677622389
transform 1 0 3848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1677622389
transform 1 0 3856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1677622389
transform 1 0 3864 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_59
timestamp 1677622389
transform 1 0 3872 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1165
timestamp 1677622389
transform 1 0 3912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1677622389
transform 1 0 3920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1677622389
transform 1 0 3928 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1677622389
transform 1 0 3936 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1173
timestamp 1677622389
transform 1 0 4032 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1677622389
transform 1 0 4040 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1677622389
transform 1 0 4048 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1677622389
transform 1 0 4056 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1677622389
transform 1 0 4064 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1677622389
transform 1 0 4072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1677622389
transform 1 0 4080 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_61
timestamp 1677622389
transform 1 0 4088 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1181
timestamp 1677622389
transform 1 0 4128 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1677622389
transform 1 0 4136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1677622389
transform 1 0 4144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1677622389
transform 1 0 4152 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_108
timestamp 1677622389
transform 1 0 4160 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1190
timestamp 1677622389
transform 1 0 4176 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1677622389
transform 1 0 4184 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1677622389
transform 1 0 4192 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1677622389
transform 1 0 4200 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1677622389
transform 1 0 4208 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1677622389
transform 1 0 4216 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1677622389
transform 1 0 4224 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1677622389
transform 1 0 4232 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1677622389
transform 1 0 4240 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1677622389
transform 1 0 4248 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1677622389
transform 1 0 4256 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1677622389
transform 1 0 4264 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1677622389
transform 1 0 4272 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1677622389
transform 1 0 4280 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1677622389
transform 1 0 4288 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1677622389
transform 1 0 4296 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1677622389
transform 1 0 4304 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1677622389
transform 1 0 4312 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1677622389
transform 1 0 4320 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1677622389
transform 1 0 4328 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1677622389
transform 1 0 4336 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1677622389
transform 1 0 4344 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1221
timestamp 1677622389
transform 1 0 4440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1677622389
transform 1 0 4448 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_111
timestamp 1677622389
transform 1 0 4456 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1224
timestamp 1677622389
transform 1 0 4472 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1677622389
transform 1 0 4480 0 -1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1677622389
transform -1 0 4520 0 -1 4170
box -8 -3 40 105
use FILL  FILL_1229
timestamp 1677622389
transform 1 0 4520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1677622389
transform 1 0 4528 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1677622389
transform 1 0 4536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1677622389
transform 1 0 4544 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_62
timestamp 1677622389
transform -1 0 4592 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1233
timestamp 1677622389
transform 1 0 4592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1677622389
transform 1 0 4600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1677622389
transform 1 0 4608 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_113
timestamp 1677622389
transform -1 0 4632 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1245
timestamp 1677622389
transform 1 0 4632 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_114
timestamp 1677622389
transform -1 0 4656 0 -1 4170
box -9 -3 26 105
use OAI22X1  OAI22X1_64
timestamp 1677622389
transform 1 0 4656 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1246
timestamp 1677622389
transform 1 0 4696 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1677622389
transform 1 0 4704 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1677622389
transform 1 0 4712 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1677622389
transform 1 0 4720 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1677622389
transform 1 0 4728 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1677622389
transform 1 0 4736 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1677622389
transform 1 0 4744 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1677622389
transform 1 0 4752 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1677622389
transform 1 0 4760 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1677622389
transform 1 0 4768 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1677622389
transform 1 0 4776 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1677622389
transform 1 0 4784 0 -1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_13
timestamp 1677622389
transform 1 0 4843 0 1 4070
box -10 -3 10 3
use M3_M2  M3_M2_1198
timestamp 1677622389
transform 1 0 164 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1677622389
transform 1 0 132 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1677622389
transform 1 0 172 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1376
timestamp 1677622389
transform 1 0 132 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1677622389
transform 1 0 164 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1677622389
transform 1 0 172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1677622389
transform 1 0 84 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1199
timestamp 1677622389
transform 1 0 212 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1677622389
transform 1 0 236 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1379
timestamp 1677622389
transform 1 0 196 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1677622389
transform 1 0 204 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1677622389
transform 1 0 220 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1677622389
transform 1 0 236 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1677622389
transform 1 0 244 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1677622389
transform 1 0 204 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1677622389
transform 1 0 212 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1677622389
transform 1 0 228 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1200
timestamp 1677622389
transform 1 0 268 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1677622389
transform 1 0 292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1677622389
transform 1 0 268 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1677622389
transform 1 0 284 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1677622389
transform 1 0 308 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1266
timestamp 1677622389
transform 1 0 308 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1677622389
transform 1 0 332 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1490
timestamp 1677622389
transform 1 0 324 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1170
timestamp 1677622389
transform 1 0 364 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1677622389
transform 1 0 364 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1386
timestamp 1677622389
transform 1 0 348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1677622389
transform 1 0 364 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1677622389
transform 1 0 356 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1187
timestamp 1677622389
transform 1 0 460 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1677622389
transform 1 0 468 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1677622389
transform 1 0 436 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1677622389
transform 1 0 476 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1388
timestamp 1677622389
transform 1 0 436 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1677622389
transform 1 0 468 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1677622389
transform 1 0 476 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1677622389
transform 1 0 388 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1188
timestamp 1677622389
transform 1 0 492 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1391
timestamp 1677622389
transform 1 0 500 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1267
timestamp 1677622389
transform 1 0 500 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1677622389
transform 1 0 524 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1677622389
transform 1 0 548 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1392
timestamp 1677622389
transform 1 0 532 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1677622389
transform 1 0 548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1677622389
transform 1 0 516 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1677622389
transform 1 0 524 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1677622389
transform 1 0 564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1677622389
transform 1 0 556 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1189
timestamp 1677622389
transform 1 0 628 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1395
timestamp 1677622389
transform 1 0 612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1677622389
transform 1 0 628 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1677622389
transform 1 0 596 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1677622389
transform 1 0 644 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1677622389
transform 1 0 740 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1677622389
transform 1 0 716 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1397
timestamp 1677622389
transform 1 0 708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1677622389
transform 1 0 740 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1222
timestamp 1677622389
transform 1 0 756 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1677622389
transform 1 0 812 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1398
timestamp 1677622389
transform 1 0 796 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1677622389
transform 1 0 852 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1677622389
transform 1 0 772 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1268
timestamp 1677622389
transform 1 0 804 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1677622389
transform 1 0 772 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1677622389
transform 1 0 836 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1677622389
transform 1 0 804 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1677622389
transform 1 0 860 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1677622389
transform 1 0 892 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1400
timestamp 1677622389
transform 1 0 932 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1677622389
transform 1 0 884 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1677622389
transform 1 0 916 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1677622389
transform 1 0 980 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1401
timestamp 1677622389
transform 1 0 980 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1269
timestamp 1677622389
transform 1 0 980 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1570
timestamp 1677622389
transform 1 0 980 0 1 3995
box -2 -2 2 2
use M3_M2  M3_M2_1224
timestamp 1677622389
transform 1 0 1028 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1501
timestamp 1677622389
transform 1 0 1020 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1677622389
transform 1 0 1028 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1225
timestamp 1677622389
transform 1 0 1052 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1402
timestamp 1677622389
transform 1 0 1044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1677622389
transform 1 0 1052 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1204
timestamp 1677622389
transform 1 0 1092 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1404
timestamp 1677622389
transform 1 0 1076 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1245
timestamp 1677622389
transform 1 0 1084 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1405
timestamp 1677622389
transform 1 0 1092 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1677622389
transform 1 0 1100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1677622389
transform 1 0 1084 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1291
timestamp 1677622389
transform 1 0 1084 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1504
timestamp 1677622389
transform 1 0 1116 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1205
timestamp 1677622389
transform 1 0 1156 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1677622389
transform 1 0 1164 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1407
timestamp 1677622389
transform 1 0 1132 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1677622389
transform 1 0 1148 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1677622389
transform 1 0 1164 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1270
timestamp 1677622389
transform 1 0 1132 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1505
timestamp 1677622389
transform 1 0 1156 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1677622389
transform 1 0 1164 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1246
timestamp 1677622389
transform 1 0 1188 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1677622389
transform 1 0 1228 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1677622389
transform 1 0 1220 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1677622389
transform 1 0 1260 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1677622389
transform 1 0 1220 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1677622389
transform 1 0 1228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1677622389
transform 1 0 1260 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1677622389
transform 1 0 1308 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1677622389
transform 1 0 1372 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1413
timestamp 1677622389
transform 1 0 1420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1677622389
transform 1 0 1452 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1677622389
transform 1 0 1372 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1292
timestamp 1677622389
transform 1 0 1420 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1677622389
transform 1 0 1460 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1509
timestamp 1677622389
transform 1 0 1460 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1229
timestamp 1677622389
transform 1 0 1508 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1415
timestamp 1677622389
transform 1 0 1492 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1677622389
transform 1 0 1508 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1248
timestamp 1677622389
transform 1 0 1524 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1510
timestamp 1677622389
transform 1 0 1500 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1677622389
transform 1 0 1516 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1677622389
transform 1 0 1524 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1293
timestamp 1677622389
transform 1 0 1500 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1677622389
transform 1 0 1540 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1677622389
transform 1 0 1588 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1677622389
transform 1 0 1572 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1677622389
transform 1 0 1588 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1249
timestamp 1677622389
transform 1 0 1596 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1513
timestamp 1677622389
transform 1 0 1564 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1677622389
transform 1 0 1580 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1677622389
transform 1 0 1596 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1677622389
transform 1 0 1612 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1231
timestamp 1677622389
transform 1 0 1628 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1516
timestamp 1677622389
transform 1 0 1644 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1232
timestamp 1677622389
transform 1 0 1740 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1677622389
transform 1 0 1780 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1420
timestamp 1677622389
transform 1 0 1740 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1677622389
transform 1 0 1772 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1677622389
transform 1 0 1780 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1677622389
transform 1 0 1692 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1271
timestamp 1677622389
transform 1 0 1724 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1677622389
transform 1 0 1692 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1677622389
transform 1 0 1716 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1518
timestamp 1677622389
transform 1 0 1788 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1677622389
transform 1 0 1804 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1677622389
transform 1 0 1828 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1677622389
transform 1 0 1820 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1191
timestamp 1677622389
transform 1 0 1836 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1520
timestamp 1677622389
transform 1 0 1836 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1307
timestamp 1677622389
transform 1 0 1860 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1677622389
transform 1 0 1884 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1425
timestamp 1677622389
transform 1 0 1884 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1178
timestamp 1677622389
transform 1 0 1916 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1677622389
transform 1 0 1956 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1426
timestamp 1677622389
transform 1 0 1948 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1677622389
transform 1 0 1956 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1677622389
transform 1 0 1996 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1296
timestamp 1677622389
transform 1 0 1996 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1522
timestamp 1677622389
transform 1 0 2012 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1308
timestamp 1677622389
transform 1 0 2012 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1523
timestamp 1677622389
transform 1 0 2028 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1677622389
transform 1 0 2044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1677622389
transform 1 0 2060 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1297
timestamp 1677622389
transform 1 0 2060 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1677622389
transform 1 0 2084 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1677622389
transform 1 0 2076 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1430
timestamp 1677622389
transform 1 0 2084 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1251
timestamp 1677622389
transform 1 0 2092 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1677622389
transform 1 0 2108 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1677622389
transform 1 0 2108 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1431
timestamp 1677622389
transform 1 0 2100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1677622389
transform 1 0 2108 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1677622389
transform 1 0 2092 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1677622389
transform 1 0 2100 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1309
timestamp 1677622389
transform 1 0 2084 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1677622389
transform 1 0 2124 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1677622389
transform 1 0 2140 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1433
timestamp 1677622389
transform 1 0 2148 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1677622389
transform 1 0 2140 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1272
timestamp 1677622389
transform 1 0 2148 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1677622389
transform 1 0 2148 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1434
timestamp 1677622389
transform 1 0 2188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1677622389
transform 1 0 2212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1677622389
transform 1 0 2220 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1677622389
transform 1 0 2260 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1677622389
transform 1 0 2284 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1273
timestamp 1677622389
transform 1 0 2284 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1528
timestamp 1677622389
transform 1 0 2316 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1173
timestamp 1677622389
transform 1 0 2332 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1438
timestamp 1677622389
transform 1 0 2332 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1311
timestamp 1677622389
transform 1 0 2324 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1677622389
transform 1 0 2364 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1439
timestamp 1677622389
transform 1 0 2364 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1677622389
transform 1 0 2380 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1677622389
transform 1 0 2348 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1677622389
transform 1 0 2396 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1253
timestamp 1677622389
transform 1 0 2404 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1677622389
transform 1 0 2396 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1530
timestamp 1677622389
transform 1 0 2404 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1298
timestamp 1677622389
transform 1 0 2388 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1677622389
transform 1 0 2420 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1677622389
transform 1 0 2436 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1677622389
transform 1 0 2428 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1677622389
transform 1 0 2428 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1677622389
transform 1 0 2436 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1210
timestamp 1677622389
transform 1 0 2556 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1442
timestamp 1677622389
transform 1 0 2468 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1677622389
transform 1 0 2476 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1255
timestamp 1677622389
transform 1 0 2484 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1444
timestamp 1677622389
transform 1 0 2508 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1275
timestamp 1677622389
transform 1 0 2468 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1677622389
transform 1 0 2508 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1677622389
transform 1 0 2556 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1299
timestamp 1677622389
transform 1 0 2556 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1534
timestamp 1677622389
transform 1 0 2580 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1182
timestamp 1677622389
transform 1 0 2596 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1677622389
transform 1 0 2660 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1445
timestamp 1677622389
transform 1 0 2604 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1677622389
transform 1 0 2612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1677622389
transform 1 0 2644 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1277
timestamp 1677622389
transform 1 0 2604 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1677622389
transform 1 0 2644 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1535
timestamp 1677622389
transform 1 0 2692 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1312
timestamp 1677622389
transform 1 0 2612 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1448
timestamp 1677622389
transform 1 0 2756 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1256
timestamp 1677622389
transform 1 0 2804 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1449
timestamp 1677622389
transform 1 0 2812 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1677622389
transform 1 0 2820 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1677622389
transform 1 0 2732 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1279
timestamp 1677622389
transform 1 0 2796 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1677622389
transform 1 0 2828 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1677622389
transform 1 0 2820 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1537
timestamp 1677622389
transform 1 0 2828 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1677622389
transform 1 0 2852 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1677622389
transform 1 0 2860 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1677622389
transform 1 0 2884 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1677622389
transform 1 0 2892 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1313
timestamp 1677622389
transform 1 0 2892 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1540
timestamp 1677622389
transform 1 0 2916 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1677622389
transform 1 0 2940 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1677622389
transform 1 0 2964 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1211
timestamp 1677622389
transform 1 0 2988 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1541
timestamp 1677622389
transform 1 0 3004 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1314
timestamp 1677622389
transform 1 0 3004 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1677622389
transform 1 0 3036 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1453
timestamp 1677622389
transform 1 0 3052 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1677622389
transform 1 0 3100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1677622389
transform 1 0 3020 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1235
timestamp 1677622389
transform 1 0 3172 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1677622389
transform 1 0 3172 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1455
timestamp 1677622389
transform 1 0 3236 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1677622389
transform 1 0 3212 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1315
timestamp 1677622389
transform 1 0 3228 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1456
timestamp 1677622389
transform 1 0 3332 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1316
timestamp 1677622389
transform 1 0 3332 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1677622389
transform 1 0 3396 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1544
timestamp 1677622389
transform 1 0 3396 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1258
timestamp 1677622389
transform 1 0 3412 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1457
timestamp 1677622389
transform 1 0 3420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1677622389
transform 1 0 3436 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1183
timestamp 1677622389
transform 1 0 3452 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1677622389
transform 1 0 3452 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1459
timestamp 1677622389
transform 1 0 3460 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1677622389
transform 1 0 3412 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1677622389
transform 1 0 3428 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1677622389
transform 1 0 3444 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1301
timestamp 1677622389
transform 1 0 3444 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1460
timestamp 1677622389
transform 1 0 3484 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1237
timestamp 1677622389
transform 1 0 3516 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1677622389
transform 1 0 3548 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1677622389
transform 1 0 3572 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1677622389
transform 1 0 3556 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1677622389
transform 1 0 3596 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1461
timestamp 1677622389
transform 1 0 3564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1677622389
transform 1 0 3580 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1261
timestamp 1677622389
transform 1 0 3588 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1548
timestamp 1677622389
transform 1 0 3548 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1677622389
transform 1 0 3556 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1677622389
transform 1 0 3572 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1677622389
transform 1 0 3588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1302
timestamp 1677622389
transform 1 0 3588 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1677622389
transform 1 0 3556 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1677622389
transform 1 0 3580 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1463
timestamp 1677622389
transform 1 0 3604 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1262
timestamp 1677622389
transform 1 0 3620 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1677622389
transform 1 0 3612 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1677622389
transform 1 0 3724 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1677622389
transform 1 0 3684 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1677622389
transform 1 0 3684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1677622389
transform 1 0 3724 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1213
timestamp 1677622389
transform 1 0 3740 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1465
timestamp 1677622389
transform 1 0 3740 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1677622389
transform 1 0 3804 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1677622389
transform 1 0 3788 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1677622389
transform 1 0 3796 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1677622389
transform 1 0 3828 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1677622389
transform 1 0 3860 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1303
timestamp 1677622389
transform 1 0 3860 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1467
timestamp 1677622389
transform 1 0 3940 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1677622389
transform 1 0 3892 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1677622389
transform 1 0 4028 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1281
timestamp 1677622389
transform 1 0 4028 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1469
timestamp 1677622389
transform 1 0 4092 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1677622389
transform 1 0 4044 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1282
timestamp 1677622389
transform 1 0 4068 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1677622389
transform 1 0 4092 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1677622389
transform 1 0 4036 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1677622389
transform 1 0 4132 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1470
timestamp 1677622389
transform 1 0 4172 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1677622389
transform 1 0 4252 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1677622389
transform 1 0 4212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1677622389
transform 1 0 4228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1677622389
transform 1 0 4244 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1677622389
transform 1 0 4204 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1677622389
transform 1 0 4260 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1677622389
transform 1 0 4252 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1263
timestamp 1677622389
transform 1 0 4268 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1561
timestamp 1677622389
transform 1 0 4268 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1241
timestamp 1677622389
transform 1 0 4308 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1475
timestamp 1677622389
transform 1 0 4308 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1677622389
transform 1 0 4300 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1285
timestamp 1677622389
transform 1 0 4308 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1563
timestamp 1677622389
transform 1 0 4324 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1677622389
transform 1 0 4380 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1677622389
transform 1 0 4356 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1677622389
transform 1 0 4380 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1677622389
transform 1 0 4468 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1477
timestamp 1677622389
transform 1 0 4468 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1677622389
transform 1 0 4476 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1184
timestamp 1677622389
transform 1 0 4516 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1677622389
transform 1 0 4492 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1479
timestamp 1677622389
transform 1 0 4516 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1185
timestamp 1677622389
transform 1 0 4556 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1677622389
transform 1 0 4540 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1677622389
transform 1 0 4564 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1480
timestamp 1677622389
transform 1 0 4564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1677622389
transform 1 0 4492 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1677622389
transform 1 0 4508 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1677622389
transform 1 0 4524 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1677622389
transform 1 0 4540 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1304
timestamp 1677622389
transform 1 0 4508 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1677622389
transform 1 0 4564 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1677622389
transform 1 0 4660 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1677622389
transform 1 0 4684 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1677622389
transform 1 0 4676 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1481
timestamp 1677622389
transform 1 0 4684 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1244
timestamp 1677622389
transform 1 0 4732 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1482
timestamp 1677622389
transform 1 0 4732 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1677622389
transform 1 0 4788 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1677622389
transform 1 0 4708 0 1 4005
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_14
timestamp 1677622389
transform 1 0 48 0 1 3970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_97
timestamp 1677622389
transform 1 0 72 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_116
timestamp 1677622389
transform -1 0 184 0 1 3970
box -9 -3 26 105
use FILL  FILL_1266
timestamp 1677622389
transform 1 0 184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1677622389
transform 1 0 192 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_63
timestamp 1677622389
transform -1 0 240 0 1 3970
box -8 -3 46 105
use FILL  FILL_1270
timestamp 1677622389
transform 1 0 240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1677622389
transform 1 0 248 0 1 3970
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1677622389
transform 1 0 256 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_65
timestamp 1677622389
transform 1 0 264 0 1 3970
box -8 -3 46 105
use FILL  FILL_1275
timestamp 1677622389
transform 1 0 304 0 1 3970
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1677622389
transform 1 0 312 0 1 3970
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1677622389
transform 1 0 320 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_66
timestamp 1677622389
transform -1 0 368 0 1 3970
box -8 -3 46 105
use FILL  FILL_1281
timestamp 1677622389
transform 1 0 368 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1677622389
transform 1 0 376 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_118
timestamp 1677622389
transform -1 0 488 0 1 3970
box -9 -3 26 105
use FILL  FILL_1282
timestamp 1677622389
transform 1 0 488 0 1 3970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1677622389
transform 1 0 496 0 1 3970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1677622389
transform 1 0 504 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_67
timestamp 1677622389
transform -1 0 552 0 1 3970
box -8 -3 46 105
use FILL  FILL_1292
timestamp 1677622389
transform 1 0 552 0 1 3970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1677622389
transform 1 0 560 0 1 3970
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1677622389
transform 1 0 568 0 1 3970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1677622389
transform 1 0 576 0 1 3970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1677622389
transform 1 0 584 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1321
timestamp 1677622389
transform 1 0 612 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_69
timestamp 1677622389
transform 1 0 592 0 1 3970
box -8 -3 46 105
use FILL  FILL_1303
timestamp 1677622389
transform 1 0 632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1677622389
transform 1 0 640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1677622389
transform 1 0 648 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1322
timestamp 1677622389
transform 1 0 700 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_101
timestamp 1677622389
transform -1 0 752 0 1 3970
box -8 -3 104 105
use FILL  FILL_1306
timestamp 1677622389
transform 1 0 752 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1677622389
transform 1 0 760 0 1 3970
box -8 -3 104 105
use FILL  FILL_1317
timestamp 1677622389
transform 1 0 856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1677622389
transform 1 0 864 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1677622389
transform 1 0 872 0 1 3970
box -8 -3 104 105
use FILL  FILL_1319
timestamp 1677622389
transform 1 0 968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1677622389
transform 1 0 976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1677622389
transform 1 0 984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1677622389
transform 1 0 992 0 1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1677622389
transform 1 0 1000 0 1 3970
box -8 -3 32 105
use FILL  FILL_1323
timestamp 1677622389
transform 1 0 1024 0 1 3970
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1677622389
transform 1 0 1032 0 1 3970
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1677622389
transform 1 0 1040 0 1 3970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1677622389
transform 1 0 1048 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_71
timestamp 1677622389
transform -1 0 1096 0 1 3970
box -8 -3 46 105
use FILL  FILL_1339
timestamp 1677622389
transform 1 0 1096 0 1 3970
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1677622389
transform 1 0 1104 0 1 3970
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1677622389
transform 1 0 1112 0 1 3970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1677622389
transform 1 0 1120 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1323
timestamp 1677622389
transform 1 0 1148 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1677622389
transform 1 0 1172 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_72
timestamp 1677622389
transform 1 0 1128 0 1 3970
box -8 -3 46 105
use FILL  FILL_1351
timestamp 1677622389
transform 1 0 1168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1677622389
transform 1 0 1176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1677622389
transform 1 0 1184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1677622389
transform 1 0 1192 0 1 3970
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1677622389
transform 1 0 1200 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_125
timestamp 1677622389
transform 1 0 1208 0 1 3970
box -9 -3 26 105
use M3_M2  M3_M2_1325
timestamp 1677622389
transform 1 0 1316 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_105
timestamp 1677622389
transform -1 0 1320 0 1 3970
box -8 -3 104 105
use FILL  FILL_1366
timestamp 1677622389
transform 1 0 1320 0 1 3970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1677622389
transform 1 0 1328 0 1 3970
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1677622389
transform 1 0 1336 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1326
timestamp 1677622389
transform 1 0 1356 0 1 3975
box -3 -3 3 3
use FILL  FILL_1378
timestamp 1677622389
transform 1 0 1344 0 1 3970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1677622389
transform 1 0 1352 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1677622389
transform 1 0 1360 0 1 3970
box -8 -3 104 105
use FILL  FILL_1381
timestamp 1677622389
transform 1 0 1456 0 1 3970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1677622389
transform 1 0 1464 0 1 3970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1677622389
transform 1 0 1472 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_67
timestamp 1677622389
transform -1 0 1520 0 1 3970
box -8 -3 46 105
use FILL  FILL_1384
timestamp 1677622389
transform 1 0 1520 0 1 3970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1677622389
transform 1 0 1528 0 1 3970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1677622389
transform 1 0 1536 0 1 3970
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1677622389
transform 1 0 1544 0 1 3970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1677622389
transform 1 0 1552 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_68
timestamp 1677622389
transform -1 0 1600 0 1 3970
box -8 -3 46 105
use FILL  FILL_1398
timestamp 1677622389
transform 1 0 1600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1677622389
transform 1 0 1608 0 1 3970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1677622389
transform 1 0 1616 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_128
timestamp 1677622389
transform -1 0 1640 0 1 3970
box -9 -3 26 105
use FILL  FILL_1401
timestamp 1677622389
transform 1 0 1640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1677622389
transform 1 0 1648 0 1 3970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1677622389
transform 1 0 1656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1677622389
transform 1 0 1664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1677622389
transform 1 0 1672 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1677622389
transform 1 0 1680 0 1 3970
box -8 -3 104 105
use FILL  FILL_1410
timestamp 1677622389
transform 1 0 1776 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_129
timestamp 1677622389
transform 1 0 1784 0 1 3970
box -9 -3 26 105
use FILL  FILL_1411
timestamp 1677622389
transform 1 0 1800 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_130
timestamp 1677622389
transform -1 0 1824 0 1 3970
box -9 -3 26 105
use FILL  FILL_1412
timestamp 1677622389
transform 1 0 1824 0 1 3970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1677622389
transform 1 0 1832 0 1 3970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1677622389
transform 1 0 1840 0 1 3970
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1677622389
transform 1 0 1848 0 1 3970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1677622389
transform 1 0 1856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1677622389
transform 1 0 1864 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1677622389
transform 1 0 1872 0 1 3970
box -9 -3 26 105
use FILL  FILL_1433
timestamp 1677622389
transform 1 0 1888 0 1 3970
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1677622389
transform 1 0 1896 0 1 3970
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1677622389
transform 1 0 1904 0 1 3970
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1677622389
transform 1 0 1912 0 1 3970
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1677622389
transform 1 0 1920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1677622389
transform 1 0 1928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1677622389
transform 1 0 1936 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_134
timestamp 1677622389
transform -1 0 1960 0 1 3970
box -9 -3 26 105
use FILL  FILL_1444
timestamp 1677622389
transform 1 0 1960 0 1 3970
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1677622389
transform 1 0 1968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1677622389
transform 1 0 1976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1677622389
transform 1 0 1984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1677622389
transform 1 0 1992 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_135
timestamp 1677622389
transform -1 0 2016 0 1 3970
box -9 -3 26 105
use FILL  FILL_1449
timestamp 1677622389
transform 1 0 2016 0 1 3970
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1677622389
transform 1 0 2024 0 1 3970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1677622389
transform 1 0 2032 0 1 3970
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1677622389
transform 1 0 2040 0 1 3970
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1677622389
transform 1 0 2048 0 1 3970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1677622389
transform 1 0 2056 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1327
timestamp 1677622389
transform 1 0 2084 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_74
timestamp 1677622389
transform -1 0 2104 0 1 3970
box -8 -3 46 105
use FILL  FILL_1459
timestamp 1677622389
transform 1 0 2104 0 1 3970
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1677622389
transform 1 0 2112 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1328
timestamp 1677622389
transform 1 0 2148 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_136
timestamp 1677622389
transform 1 0 2120 0 1 3970
box -9 -3 26 105
use FILL  FILL_1467
timestamp 1677622389
transform 1 0 2136 0 1 3970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1677622389
transform 1 0 2144 0 1 3970
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1677622389
transform 1 0 2152 0 1 3970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1677622389
transform 1 0 2160 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_76
timestamp 1677622389
transform 1 0 2168 0 1 3970
box -8 -3 46 105
use FILL  FILL_1474
timestamp 1677622389
transform 1 0 2208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1677622389
transform 1 0 2216 0 1 3970
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1677622389
transform 1 0 2224 0 1 3970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1677622389
transform 1 0 2232 0 1 3970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1677622389
transform 1 0 2240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1677622389
transform 1 0 2248 0 1 3970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1677622389
transform 1 0 2256 0 1 3970
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1677622389
transform 1 0 2264 0 1 3970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1677622389
transform 1 0 2272 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_8
timestamp 1677622389
transform 1 0 2280 0 1 3970
box -5 -3 28 105
use FILL  FILL_1494
timestamp 1677622389
transform 1 0 2304 0 1 3970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1677622389
transform 1 0 2312 0 1 3970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1677622389
transform 1 0 2320 0 1 3970
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1677622389
transform 1 0 2328 0 1 3970
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1677622389
transform 1 0 2336 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_77
timestamp 1677622389
transform 1 0 2344 0 1 3970
box -8 -3 46 105
use FILL  FILL_1506
timestamp 1677622389
transform 1 0 2384 0 1 3970
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1677622389
transform 1 0 2392 0 1 3970
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1677622389
transform 1 0 2400 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_9
timestamp 1677622389
transform 1 0 2408 0 1 3970
box -5 -3 28 105
use FILL  FILL_1513
timestamp 1677622389
transform 1 0 2432 0 1 3970
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1677622389
transform 1 0 2440 0 1 3970
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1677622389
transform 1 0 2448 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_137
timestamp 1677622389
transform 1 0 2456 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1677622389
transform -1 0 2568 0 1 3970
box -8 -3 104 105
use FILL  FILL_1516
timestamp 1677622389
transform 1 0 2568 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_138
timestamp 1677622389
transform 1 0 2576 0 1 3970
box -9 -3 26 105
use FILL  FILL_1517
timestamp 1677622389
transform 1 0 2592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1677622389
transform 1 0 2600 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1329
timestamp 1677622389
transform 1 0 2620 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_112
timestamp 1677622389
transform -1 0 2704 0 1 3970
box -8 -3 104 105
use FILL  FILL_1519
timestamp 1677622389
transform 1 0 2704 0 1 3970
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1677622389
transform 1 0 2712 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1330
timestamp 1677622389
transform 1 0 2732 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_114
timestamp 1677622389
transform 1 0 2720 0 1 3970
box -8 -3 104 105
use FILL  FILL_1534
timestamp 1677622389
transform 1 0 2816 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_39
timestamp 1677622389
transform 1 0 2824 0 1 3970
box -8 -3 34 105
use FILL  FILL_1544
timestamp 1677622389
transform 1 0 2856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1677622389
transform 1 0 2864 0 1 3970
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1677622389
transform 1 0 2872 0 1 3970
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1677622389
transform 1 0 2880 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1677622389
transform 1 0 2888 0 1 3970
box -8 -3 34 105
use FILL  FILL_1553
timestamp 1677622389
transform 1 0 2920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1677622389
transform 1 0 2928 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_41
timestamp 1677622389
transform -1 0 2968 0 1 3970
box -8 -3 34 105
use FILL  FILL_1558
timestamp 1677622389
transform 1 0 2968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1677622389
transform 1 0 2976 0 1 3970
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1677622389
transform 1 0 2984 0 1 3970
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1677622389
transform 1 0 2992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1677622389
transform 1 0 3000 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1677622389
transform 1 0 3008 0 1 3970
box -8 -3 104 105
use FILL  FILL_1568
timestamp 1677622389
transform 1 0 3104 0 1 3970
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1677622389
transform 1 0 3112 0 1 3970
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1677622389
transform 1 0 3120 0 1 3970
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1677622389
transform 1 0 3128 0 1 3970
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1677622389
transform 1 0 3136 0 1 3970
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1677622389
transform 1 0 3144 0 1 3970
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1677622389
transform 1 0 3152 0 1 3970
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1677622389
transform 1 0 3160 0 1 3970
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1677622389
transform 1 0 3168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1677622389
transform 1 0 3176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1677622389
transform 1 0 3184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1677622389
transform 1 0 3192 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1677622389
transform 1 0 3200 0 1 3970
box -8 -3 104 105
use FILL  FILL_1585
timestamp 1677622389
transform 1 0 3296 0 1 3970
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1677622389
transform 1 0 3304 0 1 3970
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1677622389
transform 1 0 3312 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_142
timestamp 1677622389
transform 1 0 3320 0 1 3970
box -9 -3 26 105
use FILL  FILL_1588
timestamp 1677622389
transform 1 0 3336 0 1 3970
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1677622389
transform 1 0 3344 0 1 3970
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1677622389
transform 1 0 3352 0 1 3970
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1677622389
transform 1 0 3360 0 1 3970
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1677622389
transform 1 0 3368 0 1 3970
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1677622389
transform 1 0 3376 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1331
timestamp 1677622389
transform 1 0 3396 0 1 3975
box -3 -3 3 3
use FILL  FILL_1598
timestamp 1677622389
transform 1 0 3384 0 1 3970
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1677622389
transform 1 0 3392 0 1 3970
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1677622389
transform 1 0 3400 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1332
timestamp 1677622389
transform 1 0 3420 0 1 3975
box -3 -3 3 3
use OAI22X1  OAI22X1_71
timestamp 1677622389
transform -1 0 3448 0 1 3970
box -8 -3 46 105
use FILL  FILL_1602
timestamp 1677622389
transform 1 0 3448 0 1 3970
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1677622389
transform 1 0 3456 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1333
timestamp 1677622389
transform 1 0 3476 0 1 3975
box -3 -3 3 3
use FILL  FILL_1609
timestamp 1677622389
transform 1 0 3464 0 1 3970
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1677622389
transform 1 0 3472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1677622389
transform 1 0 3480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1677622389
transform 1 0 3488 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_10
timestamp 1677622389
transform 1 0 3496 0 1 3970
box -5 -3 28 105
use FILL  FILL_1615
timestamp 1677622389
transform 1 0 3520 0 1 3970
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1677622389
transform 1 0 3528 0 1 3970
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1677622389
transform 1 0 3536 0 1 3970
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1677622389
transform 1 0 3544 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_72
timestamp 1677622389
transform -1 0 3592 0 1 3970
box -8 -3 46 105
use FILL  FILL_1622
timestamp 1677622389
transform 1 0 3592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1677622389
transform 1 0 3600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1677622389
transform 1 0 3608 0 1 3970
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1677622389
transform 1 0 3616 0 1 3970
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1677622389
transform 1 0 3624 0 1 3970
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1677622389
transform 1 0 3632 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1677622389
transform -1 0 3736 0 1 3970
box -8 -3 104 105
use FILL  FILL_1628
timestamp 1677622389
transform 1 0 3736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1677622389
transform 1 0 3744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1677622389
transform 1 0 3752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1677622389
transform 1 0 3760 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1334
timestamp 1677622389
transform 1 0 3788 0 1 3975
box -3 -3 3 3
use BUFX2  BUFX2_11
timestamp 1677622389
transform 1 0 3768 0 1 3970
box -5 -3 28 105
use INVX2  INVX2_144
timestamp 1677622389
transform 1 0 3792 0 1 3970
box -9 -3 26 105
use FILL  FILL_1632
timestamp 1677622389
transform 1 0 3808 0 1 3970
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1677622389
transform 1 0 3816 0 1 3970
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1677622389
transform 1 0 3824 0 1 3970
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1677622389
transform 1 0 3832 0 1 3970
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1677622389
transform 1 0 3840 0 1 3970
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1677622389
transform 1 0 3848 0 1 3970
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1677622389
transform 1 0 3856 0 1 3970
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1677622389
transform 1 0 3864 0 1 3970
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1677622389
transform 1 0 3872 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1335
timestamp 1677622389
transform 1 0 3892 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_122
timestamp 1677622389
transform 1 0 3880 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_146
timestamp 1677622389
transform 1 0 3976 0 1 3970
box -9 -3 26 105
use FILL  FILL_1652
timestamp 1677622389
transform 1 0 3992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1677622389
transform 1 0 4000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1677622389
transform 1 0 4008 0 1 3970
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1677622389
transform 1 0 4016 0 1 3970
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1677622389
transform 1 0 4024 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1677622389
transform 1 0 4032 0 1 3970
box -8 -3 104 105
use FILL  FILL_1664
timestamp 1677622389
transform 1 0 4128 0 1 3970
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1677622389
transform 1 0 4136 0 1 3970
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1677622389
transform 1 0 4144 0 1 3970
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1677622389
transform 1 0 4152 0 1 3970
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1677622389
transform 1 0 4160 0 1 3970
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1677622389
transform 1 0 4168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1677622389
transform 1 0 4176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1677622389
transform 1 0 4184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1677622389
transform 1 0 4192 0 1 3970
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1677622389
transform 1 0 4200 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_82
timestamp 1677622389
transform -1 0 4248 0 1 3970
box -8 -3 46 105
use FILL  FILL_1683
timestamp 1677622389
transform 1 0 4248 0 1 3970
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1677622389
transform 1 0 4256 0 1 3970
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1677622389
transform 1 0 4264 0 1 3970
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1677622389
transform 1 0 4272 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_76
timestamp 1677622389
transform 1 0 4280 0 1 3970
box -8 -3 46 105
use FILL  FILL_1692
timestamp 1677622389
transform 1 0 4320 0 1 3970
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1677622389
transform 1 0 4328 0 1 3970
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1677622389
transform 1 0 4336 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1677622389
transform 1 0 4344 0 1 3970
box -8 -3 104 105
use FILL  FILL_1697
timestamp 1677622389
transform 1 0 4440 0 1 3970
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1677622389
transform 1 0 4448 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_148
timestamp 1677622389
transform 1 0 4456 0 1 3970
box -9 -3 26 105
use FILL  FILL_1702
timestamp 1677622389
transform 1 0 4472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1677622389
transform 1 0 4480 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_78
timestamp 1677622389
transform 1 0 4488 0 1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1677622389
transform 1 0 4528 0 1 3970
box -8 -3 104 105
use FILL  FILL_1708
timestamp 1677622389
transform 1 0 4624 0 1 3970
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1677622389
transform 1 0 4632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1677622389
transform 1 0 4640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1677622389
transform 1 0 4648 0 1 3970
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1677622389
transform 1 0 4656 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1336
timestamp 1677622389
transform 1 0 4692 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_149
timestamp 1677622389
transform 1 0 4664 0 1 3970
box -9 -3 26 105
use FILL  FILL_1713
timestamp 1677622389
transform 1 0 4680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1677622389
transform 1 0 4688 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1337
timestamp 1677622389
transform 1 0 4724 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_128
timestamp 1677622389
transform 1 0 4696 0 1 3970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_15
timestamp 1677622389
transform 1 0 4819 0 1 3970
box -10 -3 10 3
use M2_M1  M2_M1_1576
timestamp 1677622389
transform 1 0 84 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1677622389
transform 1 0 132 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1677622389
transform 1 0 164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1677622389
transform 1 0 172 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1427
timestamp 1677622389
transform 1 0 132 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1677622389
transform 1 0 172 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1677622389
transform 1 0 164 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1577
timestamp 1677622389
transform 1 0 204 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1677622389
transform 1 0 212 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1677622389
transform 1 0 228 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1677622389
transform 1 0 196 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1512
timestamp 1677622389
transform 1 0 196 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1674
timestamp 1677622389
transform 1 0 220 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1452
timestamp 1677622389
transform 1 0 212 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1677622389
transform 1 0 260 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1677622389
transform 1 0 268 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1580
timestamp 1677622389
transform 1 0 260 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1677622389
transform 1 0 268 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1677622389
transform 1 0 284 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1677622389
transform 1 0 292 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1513
timestamp 1677622389
transform 1 0 252 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1675
timestamp 1677622389
transform 1 0 276 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1677622389
transform 1 0 292 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1677622389
transform 1 0 284 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1677
timestamp 1677622389
transform 1 0 308 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1485
timestamp 1677622389
transform 1 0 324 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1677622389
transform 1 0 356 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1677622389
transform 1 0 452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1677622389
transform 1 0 364 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1677622389
transform 1 0 372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1677622389
transform 1 0 404 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1429
timestamp 1677622389
transform 1 0 364 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1677622389
transform 1 0 404 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1677622389
transform 1 0 372 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1677622389
transform 1 0 436 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1681
timestamp 1677622389
transform 1 0 468 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1677622389
transform 1 0 468 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1682
timestamp 1677622389
transform 1 0 500 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1369
timestamp 1677622389
transform 1 0 556 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1585
timestamp 1677622389
transform 1 0 532 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1677622389
transform 1 0 540 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1677622389
transform 1 0 556 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1398
timestamp 1677622389
transform 1 0 540 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1683
timestamp 1677622389
transform 1 0 548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1677622389
transform 1 0 564 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1431
timestamp 1677622389
transform 1 0 532 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1677622389
transform 1 0 564 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1588
timestamp 1677622389
transform 1 0 588 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1399
timestamp 1677622389
transform 1 0 588 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1677622389
transform 1 0 604 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1677622389
transform 1 0 628 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1589
timestamp 1677622389
transform 1 0 628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1677622389
transform 1 0 644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1677622389
transform 1 0 620 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1677622389
transform 1 0 644 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1432
timestamp 1677622389
transform 1 0 620 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1591
timestamp 1677622389
transform 1 0 668 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1401
timestamp 1677622389
transform 1 0 668 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1677622389
transform 1 0 700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1677622389
transform 1 0 700 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1677622389
transform 1 0 708 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1370
timestamp 1677622389
transform 1 0 764 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1677622389
transform 1 0 796 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1593
timestamp 1677622389
transform 1 0 772 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1677622389
transform 1 0 780 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1677622389
transform 1 0 764 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1677622389
transform 1 0 772 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1677622389
transform 1 0 788 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1455
timestamp 1677622389
transform 1 0 780 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1677622389
transform 1 0 772 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1692
timestamp 1677622389
transform 1 0 820 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1433
timestamp 1677622389
transform 1 0 812 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1677622389
transform 1 0 804 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1677622389
transform 1 0 820 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1677622389
transform 1 0 844 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1595
timestamp 1677622389
transform 1 0 844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1677622389
transform 1 0 860 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1384
timestamp 1677622389
transform 1 0 932 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1693
timestamp 1677622389
transform 1 0 892 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1402
timestamp 1677622389
transform 1 0 932 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1677622389
transform 1 0 852 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1677622389
transform 1 0 924 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1677622389
transform 1 0 876 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1677622389
transform 1 0 948 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1573
timestamp 1677622389
transform 1 0 948 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1677622389
transform 1 0 956 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1349
timestamp 1677622389
transform 1 0 1004 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1677622389
transform 1 0 996 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1597
timestamp 1677622389
transform 1 0 980 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1677622389
transform 1 0 996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1677622389
transform 1 0 996 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1677622389
transform 1 0 1004 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1434
timestamp 1677622389
transform 1 0 1004 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1677622389
transform 1 0 996 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1677622389
transform 1 0 1036 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1599
timestamp 1677622389
transform 1 0 1028 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1385
timestamp 1677622389
transform 1 0 1036 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1697
timestamp 1677622389
transform 1 0 1036 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1494
timestamp 1677622389
transform 1 0 1028 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1677622389
transform 1 0 1068 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1779
timestamp 1677622389
transform 1 0 1060 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1677622389
transform 1 0 1084 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1600
timestamp 1677622389
transform 1 0 1076 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1339
timestamp 1677622389
transform 1 0 1100 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1677622389
transform 1 0 1108 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1571
timestamp 1677622389
transform 1 0 1116 0 1 3955
box -2 -2 2 2
use M3_M2  M3_M2_1435
timestamp 1677622389
transform 1 0 1108 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1677622389
transform 1 0 1172 0 1 3955
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1677622389
transform 1 0 1220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1677622389
transform 1 0 1220 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1677622389
transform 1 0 1244 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1403
timestamp 1677622389
transform 1 0 1244 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1780
timestamp 1677622389
transform 1 0 1284 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1677622389
transform 1 0 1316 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1495
timestamp 1677622389
transform 1 0 1300 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1677622389
transform 1 0 1316 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1603
timestamp 1677622389
transform 1 0 1348 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1458
timestamp 1677622389
transform 1 0 1348 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1604
timestamp 1677622389
transform 1 0 1364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1677622389
transform 1 0 1452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1677622389
transform 1 0 1412 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1677622389
transform 1 0 1444 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1436
timestamp 1677622389
transform 1 0 1412 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1677622389
transform 1 0 1364 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1702
timestamp 1677622389
transform 1 0 1460 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1459
timestamp 1677622389
transform 1 0 1460 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1606
timestamp 1677622389
transform 1 0 1492 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1677622389
transform 1 0 1500 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1437
timestamp 1677622389
transform 1 0 1508 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1677622389
transform 1 0 1500 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1677622389
transform 1 0 1524 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1677622389
transform 1 0 1556 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1677622389
transform 1 0 1580 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1677622389
transform 1 0 1612 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1607
timestamp 1677622389
transform 1 0 1652 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1677622389
transform 1 0 1612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1405
timestamp 1677622389
transform 1 0 1652 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1677622389
transform 1 0 1572 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1705
timestamp 1677622389
transform 1 0 1700 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1439
timestamp 1677622389
transform 1 0 1700 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1608
timestamp 1677622389
transform 1 0 1724 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1388
timestamp 1677622389
transform 1 0 1732 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1706
timestamp 1677622389
transform 1 0 1732 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1677622389
transform 1 0 1764 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1677622389
transform 1 0 1804 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1677622389
transform 1 0 1828 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1677622389
transform 1 0 1836 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1677622389
transform 1 0 1852 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1406
timestamp 1677622389
transform 1 0 1820 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1709
timestamp 1677622389
transform 1 0 1828 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1677622389
transform 1 0 1844 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1407
timestamp 1677622389
transform 1 0 1852 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1711
timestamp 1677622389
transform 1 0 1860 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1440
timestamp 1677622389
transform 1 0 1868 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1677622389
transform 1 0 1860 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1612
timestamp 1677622389
transform 1 0 1916 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1677622389
transform 1 0 1948 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1677622389
transform 1 0 1996 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1461
timestamp 1677622389
transform 1 0 1940 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1677622389
transform 1 0 1916 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1677622389
transform 1 0 1972 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1613
timestamp 1677622389
transform 1 0 2076 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1677622389
transform 1 0 2044 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1677622389
transform 1 0 2060 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1677622389
transform 1 0 2084 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1677622389
transform 1 0 2108 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1677622389
transform 1 0 2220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1677622389
transform 1 0 2244 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1516
timestamp 1677622389
transform 1 0 2244 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1616
timestamp 1677622389
transform 1 0 2292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1677622389
transform 1 0 2324 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1677622389
transform 1 0 2348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1677622389
transform 1 0 2356 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1408
timestamp 1677622389
transform 1 0 2364 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1677622389
transform 1 0 2380 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1618
timestamp 1677622389
transform 1 0 2380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1677622389
transform 1 0 2372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1677622389
transform 1 0 2396 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1409
timestamp 1677622389
transform 1 0 2396 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1677622389
transform 1 0 2500 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1677622389
transform 1 0 2484 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1677622389
transform 1 0 2452 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1677622389
transform 1 0 2500 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1677622389
transform 1 0 2532 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1677622389
transform 1 0 2444 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1677622389
transform 1 0 2452 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1677622389
transform 1 0 2500 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1462
timestamp 1677622389
transform 1 0 2444 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1677622389
transform 1 0 2500 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1677622389
transform 1 0 2532 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1724
timestamp 1677622389
transform 1 0 2556 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1464
timestamp 1677622389
transform 1 0 2564 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1677622389
transform 1 0 2580 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1621
timestamp 1677622389
transform 1 0 2580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1677622389
transform 1 0 2588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1677622389
transform 1 0 2612 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1677622389
transform 1 0 2612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1379
timestamp 1677622389
transform 1 0 2628 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1677622389
transform 1 0 2628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1677622389
transform 1 0 2620 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1465
timestamp 1677622389
transform 1 0 2612 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1624
timestamp 1677622389
transform 1 0 2668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1677622389
transform 1 0 2676 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1677622389
transform 1 0 2660 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1410
timestamp 1677622389
transform 1 0 2668 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1729
timestamp 1677622389
transform 1 0 2676 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1466
timestamp 1677622389
transform 1 0 2652 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1677622389
transform 1 0 2676 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1730
timestamp 1677622389
transform 1 0 2756 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1677622389
transform 1 0 2772 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1677622389
transform 1 0 2788 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1411
timestamp 1677622389
transform 1 0 2788 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1677622389
transform 1 0 2812 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1677622389
transform 1 0 2820 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1677622389
transform 1 0 2820 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1413
timestamp 1677622389
transform 1 0 2828 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1781
timestamp 1677622389
transform 1 0 2828 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1677622389
transform 1 0 2868 0 1 3945
box -2 -2 2 2
use M3_M2  M3_M2_1501
timestamp 1677622389
transform 1 0 2868 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1677622389
transform 1 0 2892 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1628
timestamp 1677622389
transform 1 0 2892 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1677622389
transform 1 0 2900 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1677622389
transform 1 0 2908 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1677622389
transform 1 0 2884 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1414
timestamp 1677622389
transform 1 0 2908 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1733
timestamp 1677622389
transform 1 0 2916 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1677622389
transform 1 0 2924 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1677622389
transform 1 0 2956 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1677622389
transform 1 0 2940 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1677622389
transform 1 0 3004 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1502
timestamp 1677622389
transform 1 0 3004 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1677622389
transform 1 0 3068 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1677622389
transform 1 0 3020 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1677622389
transform 1 0 3068 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1441
timestamp 1677622389
transform 1 0 3068 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1633
timestamp 1677622389
transform 1 0 3132 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1677622389
transform 1 0 3124 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1415
timestamp 1677622389
transform 1 0 3132 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1677622389
transform 1 0 3116 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1677622389
transform 1 0 3124 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1677622389
transform 1 0 3156 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1634
timestamp 1677622389
transform 1 0 3156 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1677622389
transform 1 0 3172 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1677622389
transform 1 0 3180 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1677622389
transform 1 0 3148 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1677622389
transform 1 0 3164 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1468
timestamp 1677622389
transform 1 0 3164 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1677622389
transform 1 0 3148 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1677622389
transform 1 0 3180 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1637
timestamp 1677622389
transform 1 0 3236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1677622389
transform 1 0 3228 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1677622389
transform 1 0 3244 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1469
timestamp 1677622389
transform 1 0 3244 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1677622389
transform 1 0 3260 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1638
timestamp 1677622389
transform 1 0 3260 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1355
timestamp 1677622389
transform 1 0 3324 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1639
timestamp 1677622389
transform 1 0 3276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1677622389
transform 1 0 3324 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1417
timestamp 1677622389
transform 1 0 3340 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1677622389
transform 1 0 3276 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1677622389
transform 1 0 3356 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1677622389
transform 1 0 3428 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1677622389
transform 1 0 3420 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1742
timestamp 1677622389
transform 1 0 3396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1677622389
transform 1 0 3404 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1743
timestamp 1677622389
transform 1 0 3420 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1677622389
transform 1 0 3404 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1677622389
transform 1 0 3412 0 1 3905
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1677622389
transform 1 0 3460 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1640
timestamp 1677622389
transform 1 0 3476 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1391
timestamp 1677622389
transform 1 0 3500 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1744
timestamp 1677622389
transform 1 0 3484 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1677622389
transform 1 0 3500 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1677622389
transform 1 0 3516 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1677622389
transform 1 0 3476 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1505
timestamp 1677622389
transform 1 0 3476 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1677622389
transform 1 0 3612 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1677622389
transform 1 0 3572 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1677622389
transform 1 0 3604 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1641
timestamp 1677622389
transform 1 0 3572 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1677622389
transform 1 0 3588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1677622389
transform 1 0 3564 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1419
timestamp 1677622389
transform 1 0 3588 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1748
timestamp 1677622389
transform 1 0 3612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1420
timestamp 1677622389
transform 1 0 3652 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1749
timestamp 1677622389
transform 1 0 3668 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1472
timestamp 1677622389
transform 1 0 3588 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1677622389
transform 1 0 3612 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1677622389
transform 1 0 3692 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1677622389
transform 1 0 3748 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1643
timestamp 1677622389
transform 1 0 3772 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1677622389
transform 1 0 3692 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1677622389
transform 1 0 3748 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1360
timestamp 1677622389
transform 1 0 3796 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1677622389
transform 1 0 3804 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1677622389
transform 1 0 3812 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1644
timestamp 1677622389
transform 1 0 3828 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1393
timestamp 1677622389
transform 1 0 3836 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1645
timestamp 1677622389
transform 1 0 3844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1677622389
transform 1 0 3860 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1421
timestamp 1677622389
transform 1 0 3828 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1752
timestamp 1677622389
transform 1 0 3836 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1677622389
transform 1 0 3852 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1475
timestamp 1677622389
transform 1 0 3836 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1677622389
transform 1 0 3884 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1754
timestamp 1677622389
transform 1 0 3884 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1677622389
transform 1 0 3884 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1677622389
transform 1 0 3940 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1677622389
transform 1 0 3940 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1677622389
transform 1 0 3956 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1647
timestamp 1677622389
transform 1 0 3940 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1395
timestamp 1677622389
transform 1 0 4028 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1677622389
transform 1 0 4060 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1677622389
transform 1 0 4044 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1648
timestamp 1677622389
transform 1 0 4036 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1677622389
transform 1 0 3964 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1677622389
transform 1 0 4020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1677622389
transform 1 0 4028 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1477
timestamp 1677622389
transform 1 0 3964 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1677622389
transform 1 0 4036 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1649
timestamp 1677622389
transform 1 0 4060 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1677622389
transform 1 0 4076 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1677622389
transform 1 0 4068 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1422
timestamp 1677622389
transform 1 0 4076 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1759
timestamp 1677622389
transform 1 0 4092 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1677622389
transform 1 0 4084 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1677622389
transform 1 0 4116 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1651
timestamp 1677622389
transform 1 0 4116 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1677622389
transform 1 0 4132 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1677622389
transform 1 0 4148 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1677622389
transform 1 0 4108 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1677622389
transform 1 0 4140 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1443
timestamp 1677622389
transform 1 0 4116 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1677622389
transform 1 0 4156 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1654
timestamp 1677622389
transform 1 0 4164 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1677622389
transform 1 0 4172 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1677622389
transform 1 0 4156 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1677622389
transform 1 0 4212 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1397
timestamp 1677622389
transform 1 0 4260 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1764
timestamp 1677622389
transform 1 0 4236 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1677622389
transform 1 0 4252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1677622389
transform 1 0 4260 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1480
timestamp 1677622389
transform 1 0 4236 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1677622389
transform 1 0 4292 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1656
timestamp 1677622389
transform 1 0 4284 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1677622389
transform 1 0 4292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1677622389
transform 1 0 4308 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1677622389
transform 1 0 4324 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1444
timestamp 1677622389
transform 1 0 4284 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1767
timestamp 1677622389
transform 1 0 4316 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1423
timestamp 1677622389
transform 1 0 4324 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1677622389
transform 1 0 4316 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1660
timestamp 1677622389
transform 1 0 4348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1677622389
transform 1 0 4396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1424
timestamp 1677622389
transform 1 0 4412 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1677622389
transform 1 0 4388 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1769
timestamp 1677622389
transform 1 0 4452 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1425
timestamp 1677622389
transform 1 0 4460 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1677622389
transform 1 0 4468 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1677622389
transform 1 0 4476 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1677622389
transform 1 0 4508 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1770
timestamp 1677622389
transform 1 0 4516 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1677622389
transform 1 0 4500 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1447
timestamp 1677622389
transform 1 0 4516 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1789
timestamp 1677622389
transform 1 0 4508 0 1 3905
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1677622389
transform 1 0 4532 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1426
timestamp 1677622389
transform 1 0 4532 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1787
timestamp 1677622389
transform 1 0 4532 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1481
timestamp 1677622389
transform 1 0 4532 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1677622389
transform 1 0 4588 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1677622389
transform 1 0 4588 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1662
timestamp 1677622389
transform 1 0 4572 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1677622389
transform 1 0 4588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1677622389
transform 1 0 4564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1677622389
transform 1 0 4580 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1482
timestamp 1677622389
transform 1 0 4564 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1677622389
transform 1 0 4580 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1664
timestamp 1677622389
transform 1 0 4612 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1677622389
transform 1 0 4604 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1510
timestamp 1677622389
transform 1 0 4612 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1677622389
transform 1 0 4660 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1677622389
transform 1 0 4676 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1677622389
transform 1 0 4772 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1665
timestamp 1677622389
transform 1 0 4628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1677622389
transform 1 0 4652 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1677622389
transform 1 0 4660 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1677622389
transform 1 0 4676 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1677622389
transform 1 0 4692 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1677622389
transform 1 0 4644 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1677622389
transform 1 0 4660 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1677622389
transform 1 0 4676 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1677622389
transform 1 0 4716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1677622389
transform 1 0 4772 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1448
timestamp 1677622389
transform 1 0 4636 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1677622389
transform 1 0 4652 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1677622389
transform 1 0 4676 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1677622389
transform 1 0 4628 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1677622389
transform 1 0 4652 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1677622389
transform 1 0 4644 0 1 3895
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_16
timestamp 1677622389
transform 1 0 24 0 1 3870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_98
timestamp 1677622389
transform 1 0 72 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_117
timestamp 1677622389
transform -1 0 184 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1267
timestamp 1677622389
transform 1 0 184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1677622389
transform 1 0 192 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_64
timestamp 1677622389
transform -1 0 240 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1271
timestamp 1677622389
transform 1 0 240 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1677622389
transform 1 0 248 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_65
timestamp 1677622389
transform 1 0 256 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1276
timestamp 1677622389
transform 1 0 296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1677622389
transform 1 0 304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1677622389
transform 1 0 312 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_119
timestamp 1677622389
transform 1 0 320 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1283
timestamp 1677622389
transform 1 0 336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1677622389
transform 1 0 344 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1677622389
transform 1 0 352 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1677622389
transform 1 0 360 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1677622389
transform -1 0 464 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1287
timestamp 1677622389
transform 1 0 464 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_120
timestamp 1677622389
transform -1 0 488 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1288
timestamp 1677622389
transform 1 0 488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1677622389
transform 1 0 496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1677622389
transform 1 0 504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1677622389
transform 1 0 512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1677622389
transform 1 0 520 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_68
timestamp 1677622389
transform -1 0 568 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1298
timestamp 1677622389
transform 1 0 568 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1677622389
transform 1 0 576 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1677622389
transform 1 0 584 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1677622389
transform 1 0 592 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1677622389
transform 1 0 600 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_66
timestamp 1677622389
transform -1 0 648 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1309
timestamp 1677622389
transform 1 0 648 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1677622389
transform 1 0 656 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1677622389
transform 1 0 664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1677622389
transform 1 0 672 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_121
timestamp 1677622389
transform 1 0 680 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1677622389
transform 1 0 696 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1313
timestamp 1677622389
transform 1 0 712 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1677622389
transform 1 0 720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1677622389
transform 1 0 728 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_123
timestamp 1677622389
transform -1 0 752 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1316
timestamp 1677622389
transform 1 0 752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1677622389
transform 1 0 760 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_70
timestamp 1677622389
transform 1 0 768 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1325
timestamp 1677622389
transform 1 0 808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1677622389
transform 1 0 816 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1677622389
transform 1 0 824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1677622389
transform 1 0 832 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1677622389
transform 1 0 840 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1677622389
transform 1 0 848 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1330
timestamp 1677622389
transform 1 0 944 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1677622389
transform 1 0 952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1677622389
transform 1 0 960 0 -1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_17
timestamp 1677622389
transform 1 0 968 0 -1 3970
box -8 -3 32 105
use OAI21X1  OAI21X1_35
timestamp 1677622389
transform 1 0 992 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1333
timestamp 1677622389
transform 1 0 1024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1677622389
transform 1 0 1032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1677622389
transform 1 0 1040 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1518
timestamp 1677622389
transform 1 0 1060 0 1 3875
box -3 -3 3 3
use FILL  FILL_1340
timestamp 1677622389
transform 1 0 1048 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1677622389
transform 1 0 1056 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_124
timestamp 1677622389
transform -1 0 1080 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1342
timestamp 1677622389
transform 1 0 1080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1677622389
transform 1 0 1088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1677622389
transform 1 0 1096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1677622389
transform 1 0 1104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1677622389
transform 1 0 1112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1677622389
transform 1 0 1120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1677622389
transform 1 0 1128 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1677622389
transform 1 0 1136 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1677622389
transform 1 0 1144 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1677622389
transform 1 0 1152 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1677622389
transform 1 0 1160 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1677622389
transform 1 0 1168 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1677622389
transform 1 0 1176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1677622389
transform 1 0 1184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1677622389
transform 1 0 1192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1677622389
transform 1 0 1200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1677622389
transform 1 0 1208 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_36
timestamp 1677622389
transform 1 0 1216 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1368
timestamp 1677622389
transform 1 0 1248 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1677622389
transform 1 0 1256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1677622389
transform 1 0 1264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1677622389
transform 1 0 1272 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1677622389
transform 1 0 1280 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1519
timestamp 1677622389
transform 1 0 1316 0 1 3875
box -3 -3 3 3
use OAI21X1  OAI21X1_37
timestamp 1677622389
transform -1 0 1320 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1373
timestamp 1677622389
transform 1 0 1320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1677622389
transform 1 0 1328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1677622389
transform 1 0 1336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1677622389
transform 1 0 1344 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1677622389
transform 1 0 1352 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1386
timestamp 1677622389
transform 1 0 1448 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_126
timestamp 1677622389
transform 1 0 1456 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1387
timestamp 1677622389
transform 1 0 1472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1677622389
transform 1 0 1480 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1677622389
transform 1 0 1488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1677622389
transform 1 0 1496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1677622389
transform 1 0 1504 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_127
timestamp 1677622389
transform -1 0 1528 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_1520
timestamp 1677622389
transform 1 0 1540 0 1 3875
box -3 -3 3 3
use FILL  FILL_1392
timestamp 1677622389
transform 1 0 1528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1677622389
transform 1 0 1536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1677622389
transform 1 0 1544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1677622389
transform 1 0 1552 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1677622389
transform 1 0 1560 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1521
timestamp 1677622389
transform 1 0 1628 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_108
timestamp 1677622389
transform -1 0 1664 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1407
timestamp 1677622389
transform 1 0 1664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1677622389
transform 1 0 1672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1677622389
transform 1 0 1680 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1677622389
transform 1 0 1688 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1677622389
transform 1 0 1696 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1677622389
transform 1 0 1704 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1677622389
transform 1 0 1712 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1522
timestamp 1677622389
transform 1 0 1732 0 1 3875
box -3 -3 3 3
use FILL  FILL_1423
timestamp 1677622389
transform 1 0 1720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1677622389
transform 1 0 1728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1677622389
transform 1 0 1736 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1523
timestamp 1677622389
transform 1 0 1764 0 1 3875
box -3 -3 3 3
use INVX2  INVX2_131
timestamp 1677622389
transform 1 0 1744 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1426
timestamp 1677622389
transform 1 0 1760 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_132
timestamp 1677622389
transform -1 0 1784 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_1524
timestamp 1677622389
transform 1 0 1796 0 1 3875
box -3 -3 3 3
use FILL  FILL_1427
timestamp 1677622389
transform 1 0 1784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1677622389
transform 1 0 1792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1677622389
transform 1 0 1800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1677622389
transform 1 0 1808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1677622389
transform 1 0 1816 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1525
timestamp 1677622389
transform 1 0 1836 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_73
timestamp 1677622389
transform -1 0 1864 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1432
timestamp 1677622389
transform 1 0 1864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1677622389
transform 1 0 1872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1677622389
transform 1 0 1880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1677622389
transform 1 0 1888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1677622389
transform 1 0 1896 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1526
timestamp 1677622389
transform 1 0 1916 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_110
timestamp 1677622389
transform 1 0 1904 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1450
timestamp 1677622389
transform 1 0 2000 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1677622389
transform 1 0 2008 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1677622389
transform 1 0 2016 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1677622389
transform 1 0 2024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1677622389
transform 1 0 2032 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_75
timestamp 1677622389
transform -1 0 2080 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1461
timestamp 1677622389
transform 1 0 2080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1677622389
transform 1 0 2088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1677622389
transform 1 0 2096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1677622389
transform 1 0 2104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1677622389
transform 1 0 2112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1677622389
transform 1 0 2120 0 -1 3970
box -8 -3 16 105
use BUFX2  BUFX2_6
timestamp 1677622389
transform -1 0 2152 0 -1 3970
box -5 -3 28 105
use FILL  FILL_1471
timestamp 1677622389
transform 1 0 2152 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1677622389
transform 1 0 2160 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1677622389
transform 1 0 2168 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1677622389
transform 1 0 2176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1677622389
transform 1 0 2184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1677622389
transform 1 0 2192 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1527
timestamp 1677622389
transform 1 0 2212 0 1 3875
box -3 -3 3 3
use FILL  FILL_1479
timestamp 1677622389
transform 1 0 2200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1677622389
transform 1 0 2208 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1677622389
transform 1 0 2216 0 -1 3970
box -8 -3 16 105
use BUFX2  BUFX2_7
timestamp 1677622389
transform -1 0 2248 0 -1 3970
box -5 -3 28 105
use FILL  FILL_1487
timestamp 1677622389
transform 1 0 2248 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1677622389
transform 1 0 2256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1677622389
transform 1 0 2264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1677622389
transform 1 0 2272 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1677622389
transform 1 0 2280 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1677622389
transform 1 0 2288 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1677622389
transform 1 0 2296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1677622389
transform 1 0 2304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1677622389
transform 1 0 2312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1677622389
transform 1 0 2320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1677622389
transform 1 0 2328 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_78
timestamp 1677622389
transform 1 0 2336 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1507
timestamp 1677622389
transform 1 0 2376 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1677622389
transform 1 0 2384 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1677622389
transform 1 0 2392 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1677622389
transform 1 0 2400 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1677622389
transform 1 0 2408 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1528
timestamp 1677622389
transform 1 0 2428 0 1 3875
box -3 -3 3 3
use FILL  FILL_1521
timestamp 1677622389
transform 1 0 2416 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_139
timestamp 1677622389
transform 1 0 2424 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1522
timestamp 1677622389
transform 1 0 2440 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1677622389
transform -1 0 2544 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1523
timestamp 1677622389
transform 1 0 2544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1677622389
transform 1 0 2552 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1677622389
transform 1 0 2560 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_79
timestamp 1677622389
transform 1 0 2568 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1526
timestamp 1677622389
transform 1 0 2608 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1677622389
transform 1 0 2616 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1677622389
transform 1 0 2624 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1677622389
transform 1 0 2632 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_80
timestamp 1677622389
transform 1 0 2640 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1530
timestamp 1677622389
transform 1 0 2680 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1677622389
transform 1 0 2688 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1531
timestamp 1677622389
transform 1 0 2704 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1677622389
transform 1 0 2712 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1677622389
transform 1 0 2720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1677622389
transform 1 0 2728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1677622389
transform 1 0 2736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1677622389
transform 1 0 2744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1677622389
transform 1 0 2752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1677622389
transform 1 0 2760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1677622389
transform 1 0 2768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1677622389
transform 1 0 2776 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_38
timestamp 1677622389
transform 1 0 2784 0 -1 3970
box -8 -3 34 105
use M3_M2  M3_M2_1529
timestamp 1677622389
transform 1 0 2828 0 1 3875
box -3 -3 3 3
use FILL  FILL_1543
timestamp 1677622389
transform 1 0 2816 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1677622389
transform 1 0 2824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1677622389
transform 1 0 2832 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1677622389
transform 1 0 2840 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1530
timestamp 1677622389
transform 1 0 2860 0 1 3875
box -3 -3 3 3
use NOR2X1  NOR2X1_18
timestamp 1677622389
transform 1 0 2848 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1550
timestamp 1677622389
transform 1 0 2872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1677622389
transform 1 0 2880 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1531
timestamp 1677622389
transform 1 0 2900 0 1 3875
box -3 -3 3 3
use NOR2X1  NOR2X1_19
timestamp 1677622389
transform 1 0 2888 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1554
timestamp 1677622389
transform 1 0 2912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1677622389
transform 1 0 2920 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1677622389
transform 1 0 2928 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_42
timestamp 1677622389
transform -1 0 2968 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1559
timestamp 1677622389
transform 1 0 2968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1677622389
transform 1 0 2976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1677622389
transform 1 0 2984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1677622389
transform 1 0 2992 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1677622389
transform 1 0 3000 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1677622389
transform 1 0 3008 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_141
timestamp 1677622389
transform 1 0 3104 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1571
timestamp 1677622389
transform 1 0 3120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1677622389
transform 1 0 3128 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_69
timestamp 1677622389
transform -1 0 3176 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1580
timestamp 1677622389
transform 1 0 3176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1677622389
transform 1 0 3184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1677622389
transform 1 0 3192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1677622389
transform 1 0 3200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1677622389
transform 1 0 3208 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_70
timestamp 1677622389
transform -1 0 3256 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1596
timestamp 1677622389
transform 1 0 3256 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1677622389
transform 1 0 3264 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_143
timestamp 1677622389
transform 1 0 3360 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1597
timestamp 1677622389
transform 1 0 3376 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1677622389
transform 1 0 3384 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1677622389
transform 1 0 3392 0 -1 3970
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1677622389
transform -1 0 3432 0 -1 3970
box -8 -3 40 105
use FILL  FILL_1604
timestamp 1677622389
transform 1 0 3432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1677622389
transform 1 0 3440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1677622389
transform 1 0 3448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1677622389
transform 1 0 3456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1677622389
transform 1 0 3464 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1677622389
transform 1 0 3472 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_81
timestamp 1677622389
transform 1 0 3480 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1616
timestamp 1677622389
transform 1 0 3520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1677622389
transform 1 0 3528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1677622389
transform 1 0 3536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1677622389
transform 1 0 3544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1677622389
transform 1 0 3552 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_145
timestamp 1677622389
transform -1 0 3576 0 -1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1677622389
transform 1 0 3576 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1635
timestamp 1677622389
transform 1 0 3672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1677622389
transform 1 0 3680 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1677622389
transform -1 0 3784 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1637
timestamp 1677622389
transform 1 0 3784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1677622389
transform 1 0 3792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1677622389
transform 1 0 3800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1677622389
transform 1 0 3808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1677622389
transform 1 0 3816 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_73
timestamp 1677622389
transform -1 0 3864 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1649
timestamp 1677622389
transform 1 0 3864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1677622389
transform 1 0 3872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1677622389
transform 1 0 3880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1677622389
transform 1 0 3888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1677622389
transform 1 0 3896 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1677622389
transform 1 0 3904 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1677622389
transform 1 0 3912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1677622389
transform 1 0 3920 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1677622389
transform 1 0 3928 0 -1 3970
box -8 -3 104 105
use M3_M2  M3_M2_1532
timestamp 1677622389
transform 1 0 4036 0 1 3875
box -3 -3 3 3
use FILL  FILL_1663
timestamp 1677622389
transform 1 0 4024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1677622389
transform 1 0 4032 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_74
timestamp 1677622389
transform 1 0 4040 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1669
timestamp 1677622389
transform 1 0 4080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1677622389
transform 1 0 4088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1677622389
transform 1 0 4096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1677622389
transform 1 0 4104 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_75
timestamp 1677622389
transform 1 0 4112 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1673
timestamp 1677622389
transform 1 0 4152 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1677622389
transform 1 0 4160 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_147
timestamp 1677622389
transform 1 0 4168 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1679
timestamp 1677622389
transform 1 0 4184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1677622389
transform 1 0 4192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1677622389
transform 1 0 4200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1677622389
transform 1 0 4208 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_83
timestamp 1677622389
transform -1 0 4256 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1687
timestamp 1677622389
transform 1 0 4256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1677622389
transform 1 0 4264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1677622389
transform 1 0 4272 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1677622389
transform 1 0 4280 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_77
timestamp 1677622389
transform 1 0 4288 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1695
timestamp 1677622389
transform 1 0 4328 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1677622389
transform 1 0 4336 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1698
timestamp 1677622389
transform 1 0 4432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1677622389
transform 1 0 4440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1677622389
transform 1 0 4448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1677622389
transform 1 0 4456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1677622389
transform 1 0 4464 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1677622389
transform 1 0 4472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1677622389
transform 1 0 4480 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1677622389
transform 1 0 4488 0 -1 3970
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1677622389
transform -1 0 4528 0 -1 3970
box -8 -3 40 105
use FILL  FILL_1716
timestamp 1677622389
transform 1 0 4528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1677622389
transform 1 0 4536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1677622389
transform 1 0 4544 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_79
timestamp 1677622389
transform -1 0 4592 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1719
timestamp 1677622389
transform 1 0 4592 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1677622389
transform 1 0 4600 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1677622389
transform 1 0 4608 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1533
timestamp 1677622389
transform 1 0 4628 0 1 3875
box -3 -3 3 3
use FILL  FILL_1722
timestamp 1677622389
transform 1 0 4616 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1534
timestamp 1677622389
transform 1 0 4660 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_84
timestamp 1677622389
transform -1 0 4664 0 -1 3970
box -8 -3 46 105
use M3_M2  M3_M2_1535
timestamp 1677622389
transform 1 0 4676 0 1 3875
box -3 -3 3 3
use INVX2  INVX2_150
timestamp 1677622389
transform -1 0 4680 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_1536
timestamp 1677622389
transform 1 0 4716 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_129
timestamp 1677622389
transform 1 0 4680 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1723
timestamp 1677622389
transform 1 0 4776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1677622389
transform 1 0 4784 0 -1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_17
timestamp 1677622389
transform 1 0 4843 0 1 3870
box -10 -3 10 3
use M2_M1  M2_M1_1800
timestamp 1677622389
transform 1 0 108 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1677622389
transform 1 0 140 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1637
timestamp 1677622389
transform 1 0 140 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1677622389
transform 1 0 172 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1911
timestamp 1677622389
transform 1 0 172 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1677
timestamp 1677622389
transform 1 0 172 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1677622389
transform 1 0 204 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1677622389
transform 1 0 244 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1677622389
transform 1 0 220 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1677622389
transform 1 0 260 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1677622389
transform 1 0 276 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1801
timestamp 1677622389
transform 1 0 212 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1677622389
transform 1 0 220 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1677622389
transform 1 0 236 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1677622389
transform 1 0 252 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1677622389
transform 1 0 260 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1677622389
transform 1 0 276 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1677622389
transform 1 0 292 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1677622389
transform 1 0 220 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1677622389
transform 1 0 228 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1677622389
transform 1 0 244 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1638
timestamp 1677622389
transform 1 0 236 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1677622389
transform 1 0 244 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1915
timestamp 1677622389
transform 1 0 268 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1619
timestamp 1677622389
transform 1 0 276 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1916
timestamp 1677622389
transform 1 0 284 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1677622389
transform 1 0 308 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1620
timestamp 1677622389
transform 1 0 300 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1677622389
transform 1 0 292 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1917
timestamp 1677622389
transform 1 0 324 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1677622389
transform 1 0 356 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1621
timestamp 1677622389
transform 1 0 340 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1918
timestamp 1677622389
transform 1 0 348 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1677622389
transform 1 0 372 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1677622389
transform 1 0 436 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1677622389
transform 1 0 404 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1677622389
transform 1 0 540 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1677622389
transform 1 0 548 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1677622389
transform 1 0 604 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1677622389
transform 1 0 620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1677622389
transform 1 0 596 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1580
timestamp 1677622389
transform 1 0 644 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1677622389
transform 1 0 756 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1815
timestamp 1677622389
transform 1 0 668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1677622389
transform 1 0 700 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1677622389
transform 1 0 748 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1639
timestamp 1677622389
transform 1 0 668 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1677622389
transform 1 0 764 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1817
timestamp 1677622389
transform 1 0 764 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1556
timestamp 1677622389
transform 1 0 788 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1923
timestamp 1677622389
transform 1 0 780 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1640
timestamp 1677622389
transform 1 0 780 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1677622389
transform 1 0 828 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1677622389
transform 1 0 820 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1677622389
transform 1 0 812 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1818
timestamp 1677622389
transform 1 0 812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1677622389
transform 1 0 804 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1677622389
transform 1 0 828 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1677622389
transform 1 0 836 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1539
timestamp 1677622389
transform 1 0 876 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1677622389
transform 1 0 860 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1821
timestamp 1677622389
transform 1 0 860 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1677622389
transform 1 0 876 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1677622389
transform 1 0 844 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1677622389
transform 1 0 852 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1641
timestamp 1677622389
transform 1 0 860 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1823
timestamp 1677622389
transform 1 0 892 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1677622389
transform 1 0 892 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1680
timestamp 1677622389
transform 1 0 892 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1928
timestamp 1677622389
transform 1 0 908 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1622
timestamp 1677622389
transform 1 0 916 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1677622389
transform 1 0 932 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1677622389
transform 1 0 940 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1677622389
transform 1 0 924 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1642
timestamp 1677622389
transform 1 0 908 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2005
timestamp 1677622389
transform 1 0 916 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1643
timestamp 1677622389
transform 1 0 940 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1930
timestamp 1677622389
transform 1 0 956 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1681
timestamp 1677622389
transform 1 0 956 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1931
timestamp 1677622389
transform 1 0 1012 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1548
timestamp 1677622389
transform 1 0 1028 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1793
timestamp 1677622389
transform 1 0 1028 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1559
timestamp 1677622389
transform 1 0 1044 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1677622389
transform 1 0 1124 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1677622389
transform 1 0 1092 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1677622389
transform 1 0 1132 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1826
timestamp 1677622389
transform 1 0 1092 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1677622389
transform 1 0 1124 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1677622389
transform 1 0 1132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1677622389
transform 1 0 1044 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1540
timestamp 1677622389
transform 1 0 1148 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1677622389
transform 1 0 1156 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1829
timestamp 1677622389
transform 1 0 1148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1677622389
transform 1 0 1164 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1677622389
transform 1 0 1180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1677622389
transform 1 0 1148 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1677622389
transform 1 0 1156 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1677622389
transform 1 0 1172 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1549
timestamp 1677622389
transform 1 0 1196 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1936
timestamp 1677622389
transform 1 0 1196 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1677622389
transform 1 0 1220 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1794
timestamp 1677622389
transform 1 0 1212 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1644
timestamp 1677622389
transform 1 0 1220 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1677622389
transform 1 0 1212 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1832
timestamp 1677622389
transform 1 0 1244 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1677622389
transform 1 0 1252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1677622389
transform 1 0 1260 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1677622389
transform 1 0 1284 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1677622389
transform 1 0 1300 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1645
timestamp 1677622389
transform 1 0 1284 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1677622389
transform 1 0 1284 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1796
timestamp 1677622389
transform 1 0 1324 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1677622389
transform 1 0 1316 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1677622389
transform 1 0 1332 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1646
timestamp 1677622389
transform 1 0 1324 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1835
timestamp 1677622389
transform 1 0 1356 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1647
timestamp 1677622389
transform 1 0 1340 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1677622389
transform 1 0 1332 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1836
timestamp 1677622389
transform 1 0 1380 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1677622389
transform 1 0 1364 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1677622389
transform 1 0 1372 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1648
timestamp 1677622389
transform 1 0 1372 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1837
timestamp 1677622389
transform 1 0 1412 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1685
timestamp 1677622389
transform 1 0 1412 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1942
timestamp 1677622389
transform 1 0 1444 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1677622389
transform 1 0 1468 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1677622389
transform 1 0 1484 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1677622389
transform 1 0 1500 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1677622389
transform 1 0 1516 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1677622389
transform 1 0 1508 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1649
timestamp 1677622389
transform 1 0 1500 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1945
timestamp 1677622389
transform 1 0 1532 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1650
timestamp 1677622389
transform 1 0 1540 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1841
timestamp 1677622389
transform 1 0 1580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1677622389
transform 1 0 1556 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1651
timestamp 1677622389
transform 1 0 1556 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1677622389
transform 1 0 1580 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1842
timestamp 1677622389
transform 1 0 1668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1677622389
transform 1 0 1732 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1677622389
transform 1 0 1692 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1653
timestamp 1677622389
transform 1 0 1692 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1677622389
transform 1 0 1716 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1677622389
transform 1 0 1732 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1844
timestamp 1677622389
transform 1 0 1796 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1677622389
transform 1 0 1804 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1677622389
transform 1 0 1820 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1677622389
transform 1 0 1836 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1677622389
transform 1 0 1844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1677622389
transform 1 0 1812 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1677622389
transform 1 0 1828 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1655
timestamp 1677622389
transform 1 0 1820 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1677622389
transform 1 0 1844 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1950
timestamp 1677622389
transform 1 0 1892 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1656
timestamp 1677622389
transform 1 0 1884 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1677622389
transform 1 0 1940 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1677622389
transform 1 0 1948 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1849
timestamp 1677622389
transform 1 0 1924 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1607
timestamp 1677622389
transform 1 0 1932 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1850
timestamp 1677622389
transform 1 0 1940 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1677622389
transform 1 0 1916 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1677622389
transform 1 0 1932 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1623
timestamp 1677622389
transform 1 0 1940 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1677622389
transform 1 0 1964 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1677622389
transform 1 0 1964 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1677622389
transform 1 0 1972 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1953
timestamp 1677622389
transform 1 0 1988 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1567
timestamp 1677622389
transform 1 0 2076 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1851
timestamp 1677622389
transform 1 0 2028 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1677622389
transform 1 0 2004 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1658
timestamp 1677622389
transform 1 0 2004 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1677622389
transform 1 0 2020 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1677622389
transform 1 0 2036 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1852
timestamp 1677622389
transform 1 0 2092 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1568
timestamp 1677622389
transform 1 0 2156 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1677622389
transform 1 0 2204 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1677622389
transform 1 0 2180 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1853
timestamp 1677622389
transform 1 0 2156 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1677622389
transform 1 0 2188 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1677622389
transform 1 0 2204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1677622389
transform 1 0 2108 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1609
timestamp 1677622389
transform 1 0 2212 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1956
timestamp 1677622389
transform 1 0 2228 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1689
timestamp 1677622389
transform 1 0 2236 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1677622389
transform 1 0 2260 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1856
timestamp 1677622389
transform 1 0 2260 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1610
timestamp 1677622389
transform 1 0 2268 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1857
timestamp 1677622389
transform 1 0 2284 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1677622389
transform 1 0 2252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1677622389
transform 1 0 2268 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1570
timestamp 1677622389
transform 1 0 2308 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1677622389
transform 1 0 2324 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1858
timestamp 1677622389
transform 1 0 2372 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1677622389
transform 1 0 2380 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1541
timestamp 1677622389
transform 1 0 2484 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1677622389
transform 1 0 2476 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1677622389
transform 1 0 2476 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1859
timestamp 1677622389
transform 1 0 2444 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1677622389
transform 1 0 2476 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1677622389
transform 1 0 2492 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1677622389
transform 1 0 2508 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1611
timestamp 1677622389
transform 1 0 2532 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1861
timestamp 1677622389
transform 1 0 2540 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1612
timestamp 1677622389
transform 1 0 2548 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1862
timestamp 1677622389
transform 1 0 2564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1677622389
transform 1 0 2548 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1677622389
transform 1 0 2556 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1590
timestamp 1677622389
transform 1 0 2596 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1677622389
transform 1 0 2588 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1677622389
transform 1 0 2644 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1863
timestamp 1677622389
transform 1 0 2644 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1592
timestamp 1677622389
transform 1 0 2684 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1864
timestamp 1677622389
transform 1 0 2684 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1613
timestamp 1677622389
transform 1 0 2732 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1865
timestamp 1677622389
transform 1 0 2740 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1677622389
transform 1 0 2660 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1624
timestamp 1677622389
transform 1 0 2740 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1677622389
transform 1 0 2660 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1677622389
transform 1 0 2724 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1677622389
transform 1 0 2692 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_2006
timestamp 1677622389
transform 1 0 2748 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1542
timestamp 1677622389
transform 1 0 2772 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1677622389
transform 1 0 2804 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1677622389
transform 1 0 2812 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1866
timestamp 1677622389
transform 1 0 2820 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1677622389
transform 1 0 2804 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1677622389
transform 1 0 2812 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1677622389
transform 1 0 2804 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1677622389
transform 1 0 2852 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1867
timestamp 1677622389
transform 1 0 2852 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1677622389
transform 1 0 2884 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1677622389
transform 1 0 2924 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1677622389
transform 1 0 2948 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1593
timestamp 1677622389
transform 1 0 2972 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1968
timestamp 1677622389
transform 1 0 2972 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1677622389
transform 1 0 3036 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1677622389
transform 1 0 2988 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1664
timestamp 1677622389
transform 1 0 2988 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1677622389
transform 1 0 3084 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1870
timestamp 1677622389
transform 1 0 3084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1677622389
transform 1 0 3100 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1595
timestamp 1677622389
transform 1 0 3132 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1871
timestamp 1677622389
transform 1 0 3132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1677622389
transform 1 0 3124 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1677622389
transform 1 0 3140 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1625
timestamp 1677622389
transform 1 0 3148 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1872
timestamp 1677622389
transform 1 0 3164 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1665
timestamp 1677622389
transform 1 0 3172 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1973
timestamp 1677622389
transform 1 0 3188 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1677622389
transform 1 0 3228 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1677622389
transform 1 0 3204 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1626
timestamp 1677622389
transform 1 0 3228 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1677622389
transform 1 0 3204 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1677622389
transform 1 0 3316 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1874
timestamp 1677622389
transform 1 0 3316 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1544
timestamp 1677622389
transform 1 0 3412 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1677622389
transform 1 0 3436 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1875
timestamp 1677622389
transform 1 0 3396 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1615
timestamp 1677622389
transform 1 0 3420 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1975
timestamp 1677622389
transform 1 0 3356 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1677622389
transform 1 0 3396 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1677622389
transform 1 0 3460 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1677622389
transform 1 0 3452 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1677622389
transform 1 0 3492 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1876
timestamp 1677622389
transform 1 0 3452 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1677622389
transform 1 0 3460 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1677622389
transform 1 0 3476 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1616
timestamp 1677622389
transform 1 0 3484 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1976
timestamp 1677622389
transform 1 0 3452 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1677622389
transform 1 0 3468 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1627
timestamp 1677622389
transform 1 0 3476 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1978
timestamp 1677622389
transform 1 0 3484 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1677622389
transform 1 0 3492 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1668
timestamp 1677622389
transform 1 0 3468 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1879
timestamp 1677622389
transform 1 0 3508 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1628
timestamp 1677622389
transform 1 0 3508 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1677622389
transform 1 0 3540 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1677622389
transform 1 0 3540 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1880
timestamp 1677622389
transform 1 0 3564 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1630
timestamp 1677622389
transform 1 0 3580 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1677622389
transform 1 0 3572 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1790
timestamp 1677622389
transform 1 0 3644 0 1 3845
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1677622389
transform 1 0 3660 0 1 3845
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1677622389
transform 1 0 3660 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1677622389
transform 1 0 3724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1677622389
transform 1 0 3756 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1677622389
transform 1 0 3676 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1670
timestamp 1677622389
transform 1 0 3724 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1677622389
transform 1 0 3676 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1883
timestamp 1677622389
transform 1 0 3772 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1677622389
transform 1 0 3788 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1677622389
transform 1 0 3812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1677622389
transform 1 0 3828 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1677622389
transform 1 0 3836 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1677622389
transform 1 0 3804 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1671
timestamp 1677622389
transform 1 0 3804 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1677622389
transform 1 0 3820 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1677622389
transform 1 0 3860 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1677622389
transform 1 0 3876 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1677622389
transform 1 0 3892 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1888
timestamp 1677622389
transform 1 0 3876 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1677622389
transform 1 0 3892 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1601
timestamp 1677622389
transform 1 0 3908 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1890
timestamp 1677622389
transform 1 0 3908 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1677622389
transform 1 0 3860 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1677622389
transform 1 0 3868 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1677622389
transform 1 0 3884 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1677622389
transform 1 0 3900 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1631
timestamp 1677622389
transform 1 0 3908 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1677622389
transform 1 0 3908 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1798
timestamp 1677622389
transform 1 0 4012 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1677622389
transform 1 0 4020 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1677622389
transform 1 0 4036 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1677622389
transform 1 0 4044 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1573
timestamp 1677622389
transform 1 0 4060 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1677622389
transform 1 0 4084 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1677622389
transform 1 0 4076 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1799
timestamp 1677622389
transform 1 0 4076 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1677622389
transform 1 0 4060 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1617
timestamp 1677622389
transform 1 0 4068 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1677622389
transform 1 0 4108 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1892
timestamp 1677622389
transform 1 0 4092 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1677622389
transform 1 0 4108 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1677622389
transform 1 0 4084 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1677622389
transform 1 0 4100 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1632
timestamp 1677622389
transform 1 0 4108 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1677622389
transform 1 0 4124 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1991
timestamp 1677622389
transform 1 0 4116 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1677622389
transform 1 0 4124 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1673
timestamp 1677622389
transform 1 0 4100 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1677622389
transform 1 0 4172 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1677622389
transform 1 0 4180 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1894
timestamp 1677622389
transform 1 0 4156 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1677622389
transform 1 0 4172 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1633
timestamp 1677622389
transform 1 0 4148 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1677622389
transform 1 0 4164 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1993
timestamp 1677622389
transform 1 0 4180 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1677622389
transform 1 0 4212 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1576
timestamp 1677622389
transform 1 0 4252 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1677622389
transform 1 0 4268 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1897
timestamp 1677622389
transform 1 0 4252 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1677622389
transform 1 0 4228 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1674
timestamp 1677622389
transform 1 0 4252 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1677622389
transform 1 0 4332 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1677622389
transform 1 0 4324 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1898
timestamp 1677622389
transform 1 0 4324 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1677622389
transform 1 0 4332 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1677622389
transform 1 0 4356 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1677622389
transform 1 0 4364 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1677622389
transform 1 0 4364 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1677622389
transform 1 0 4404 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1900
timestamp 1677622389
transform 1 0 4388 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1677622389
transform 1 0 4404 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1677622389
transform 1 0 4396 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1677622389
transform 1 0 4412 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1606
timestamp 1677622389
transform 1 0 4436 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1902
timestamp 1677622389
transform 1 0 4436 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1677622389
transform 1 0 4452 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1677622389
transform 1 0 4532 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1677622389
transform 1 0 4580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1677622389
transform 1 0 4556 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1551
timestamp 1677622389
transform 1 0 4692 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1677622389
transform 1 0 4724 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1677622389
transform 1 0 4652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1677622389
transform 1 0 4668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1677622389
transform 1 0 4684 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1677622389
transform 1 0 4660 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1677622389
transform 1 0 4676 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1676
timestamp 1677622389
transform 1 0 4636 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1677622389
transform 1 0 4684 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1677622389
transform 1 0 4732 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1677622389
transform 1 0 4788 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1677622389
transform 1 0 4692 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1677622389
transform 1 0 4708 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1636
timestamp 1677622389
transform 1 0 4732 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1677622389
transform 1 0 4756 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1677622389
transform 1 0 4788 0 1 3785
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_18
timestamp 1677622389
transform 1 0 48 0 1 3770
box -10 -3 10 3
use FILL  FILL_1725
timestamp 1677622389
transform 1 0 72 0 1 3770
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1677622389
transform 1 0 80 0 1 3770
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1677622389
transform 1 0 88 0 1 3770
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1677622389
transform 1 0 96 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_151
timestamp 1677622389
transform -1 0 120 0 1 3770
box -9 -3 26 105
use FILL  FILL_1729
timestamp 1677622389
transform 1 0 120 0 1 3770
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1677622389
transform 1 0 128 0 1 3770
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1677622389
transform 1 0 136 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_152
timestamp 1677622389
transform -1 0 160 0 1 3770
box -9 -3 26 105
use FILL  FILL_1732
timestamp 1677622389
transform 1 0 160 0 1 3770
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1677622389
transform 1 0 168 0 1 3770
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1677622389
transform 1 0 176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1677622389
transform 1 0 184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1677622389
transform 1 0 192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1677622389
transform 1 0 200 0 1 3770
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1677622389
transform 1 0 208 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_85
timestamp 1677622389
transform 1 0 216 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1677622389
transform 1 0 256 0 1 3770
box -8 -3 46 105
use FILL  FILL_1740
timestamp 1677622389
transform 1 0 296 0 1 3770
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1677622389
transform 1 0 304 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1696
timestamp 1677622389
transform 1 0 324 0 1 3775
box -3 -3 3 3
use FILL  FILL_1742
timestamp 1677622389
transform 1 0 312 0 1 3770
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1677622389
transform 1 0 320 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1697
timestamp 1677622389
transform 1 0 356 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_80
timestamp 1677622389
transform 1 0 328 0 1 3770
box -8 -3 46 105
use FILL  FILL_1744
timestamp 1677622389
transform 1 0 368 0 1 3770
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1677622389
transform 1 0 376 0 1 3770
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1677622389
transform 1 0 384 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1677622389
transform 1 0 392 0 1 3770
box -8 -3 104 105
use FILL  FILL_1747
timestamp 1677622389
transform 1 0 488 0 1 3770
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1677622389
transform 1 0 496 0 1 3770
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1677622389
transform 1 0 504 0 1 3770
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1677622389
transform 1 0 512 0 1 3770
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1677622389
transform 1 0 520 0 1 3770
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1677622389
transform 1 0 528 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1698
timestamp 1677622389
transform 1 0 548 0 1 3775
box -3 -3 3 3
use FILL  FILL_1762
timestamp 1677622389
transform 1 0 536 0 1 3770
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1677622389
transform 1 0 544 0 1 3770
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1677622389
transform 1 0 552 0 1 3770
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1677622389
transform 1 0 560 0 1 3770
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1677622389
transform 1 0 568 0 1 3770
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1677622389
transform 1 0 576 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_88
timestamp 1677622389
transform 1 0 584 0 1 3770
box -8 -3 46 105
use FILL  FILL_1774
timestamp 1677622389
transform 1 0 624 0 1 3770
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1677622389
transform 1 0 632 0 1 3770
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1677622389
transform 1 0 640 0 1 3770
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1677622389
transform 1 0 648 0 1 3770
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1677622389
transform 1 0 656 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1677622389
transform -1 0 760 0 1 3770
box -8 -3 104 105
use FILL  FILL_1788
timestamp 1677622389
transform 1 0 760 0 1 3770
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1677622389
transform 1 0 768 0 1 3770
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1677622389
transform 1 0 776 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_82
timestamp 1677622389
transform 1 0 784 0 1 3770
box -8 -3 46 105
use FILL  FILL_1795
timestamp 1677622389
transform 1 0 824 0 1 3770
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1677622389
transform 1 0 832 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_89
timestamp 1677622389
transform 1 0 840 0 1 3770
box -8 -3 46 105
use FILL  FILL_1797
timestamp 1677622389
transform 1 0 880 0 1 3770
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1677622389
transform 1 0 888 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_154
timestamp 1677622389
transform -1 0 912 0 1 3770
box -9 -3 26 105
use NOR2X1  NOR2X1_20
timestamp 1677622389
transform 1 0 912 0 1 3770
box -8 -3 32 105
use FILL  FILL_1799
timestamp 1677622389
transform 1 0 936 0 1 3770
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1677622389
transform 1 0 944 0 1 3770
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1677622389
transform 1 0 952 0 1 3770
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1677622389
transform 1 0 960 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_43
timestamp 1677622389
transform 1 0 968 0 1 3770
box -8 -3 34 105
use FILL  FILL_1812
timestamp 1677622389
transform 1 0 1000 0 1 3770
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1677622389
transform 1 0 1008 0 1 3770
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1677622389
transform 1 0 1016 0 1 3770
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1677622389
transform 1 0 1024 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1677622389
transform 1 0 1032 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_156
timestamp 1677622389
transform -1 0 1144 0 1 3770
box -9 -3 26 105
use M3_M2  M3_M2_1699
timestamp 1677622389
transform 1 0 1180 0 1 3775
box -3 -3 3 3
use AOI22X1  AOI22X1_90
timestamp 1677622389
transform -1 0 1184 0 1 3770
box -8 -3 46 105
use FILL  FILL_1821
timestamp 1677622389
transform 1 0 1184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1677622389
transform 1 0 1192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1677622389
transform 1 0 1200 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_45
timestamp 1677622389
transform -1 0 1240 0 1 3770
box -8 -3 34 105
use FILL  FILL_1837
timestamp 1677622389
transform 1 0 1240 0 1 3770
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1677622389
transform 1 0 1248 0 1 3770
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1677622389
transform 1 0 1256 0 1 3770
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1677622389
transform 1 0 1264 0 1 3770
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1677622389
transform 1 0 1272 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_47
timestamp 1677622389
transform -1 0 1312 0 1 3770
box -8 -3 34 105
use FILL  FILL_1848
timestamp 1677622389
transform 1 0 1312 0 1 3770
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1677622389
transform 1 0 1320 0 1 3770
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1677622389
transform 1 0 1328 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_48
timestamp 1677622389
transform -1 0 1368 0 1 3770
box -8 -3 34 105
use FILL  FILL_1854
timestamp 1677622389
transform 1 0 1368 0 1 3770
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1677622389
transform 1 0 1376 0 1 3770
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1677622389
transform 1 0 1384 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_159
timestamp 1677622389
transform 1 0 1392 0 1 3770
box -9 -3 26 105
use FILL  FILL_1857
timestamp 1677622389
transform 1 0 1408 0 1 3770
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1677622389
transform 1 0 1416 0 1 3770
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1677622389
transform 1 0 1424 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_160
timestamp 1677622389
transform -1 0 1448 0 1 3770
box -9 -3 26 105
use FILL  FILL_1860
timestamp 1677622389
transform 1 0 1448 0 1 3770
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1677622389
transform 1 0 1456 0 1 3770
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1677622389
transform 1 0 1464 0 1 3770
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1677622389
transform 1 0 1472 0 1 3770
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1677622389
transform 1 0 1480 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_83
timestamp 1677622389
transform -1 0 1528 0 1 3770
box -8 -3 46 105
use FILL  FILL_1869
timestamp 1677622389
transform 1 0 1528 0 1 3770
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1677622389
transform 1 0 1536 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1677622389
transform 1 0 1544 0 1 3770
box -8 -3 104 105
use FILL  FILL_1871
timestamp 1677622389
transform 1 0 1640 0 1 3770
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1677622389
transform 1 0 1648 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_161
timestamp 1677622389
transform 1 0 1656 0 1 3770
box -9 -3 26 105
use FILL  FILL_1885
timestamp 1677622389
transform 1 0 1672 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1677622389
transform 1 0 1680 0 1 3770
box -8 -3 104 105
use FILL  FILL_1889
timestamp 1677622389
transform 1 0 1776 0 1 3770
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1677622389
transform 1 0 1784 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1700
timestamp 1677622389
transform 1 0 1804 0 1 3775
box -3 -3 3 3
use FILL  FILL_1891
timestamp 1677622389
transform 1 0 1792 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_91
timestamp 1677622389
transform 1 0 1800 0 1 3770
box -8 -3 46 105
use FILL  FILL_1893
timestamp 1677622389
transform 1 0 1840 0 1 3770
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1677622389
transform 1 0 1848 0 1 3770
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1677622389
transform 1 0 1856 0 1 3770
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1677622389
transform 1 0 1864 0 1 3770
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1677622389
transform 1 0 1872 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_163
timestamp 1677622389
transform -1 0 1896 0 1 3770
box -9 -3 26 105
use FILL  FILL_1907
timestamp 1677622389
transform 1 0 1896 0 1 3770
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1677622389
transform 1 0 1904 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_86
timestamp 1677622389
transform 1 0 1912 0 1 3770
box -8 -3 46 105
use FILL  FILL_1914
timestamp 1677622389
transform 1 0 1952 0 1 3770
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1677622389
transform 1 0 1960 0 1 3770
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1677622389
transform 1 0 1968 0 1 3770
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1677622389
transform 1 0 1976 0 1 3770
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1677622389
transform 1 0 1984 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1677622389
transform 1 0 1992 0 1 3770
box -8 -3 104 105
use FILL  FILL_1925
timestamp 1677622389
transform 1 0 2088 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1701
timestamp 1677622389
transform 1 0 2132 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_143
timestamp 1677622389
transform 1 0 2096 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_166
timestamp 1677622389
transform -1 0 2208 0 1 3770
box -9 -3 26 105
use FILL  FILL_1926
timestamp 1677622389
transform 1 0 2208 0 1 3770
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1677622389
transform 1 0 2216 0 1 3770
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1677622389
transform 1 0 2224 0 1 3770
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1677622389
transform 1 0 2232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1677622389
transform 1 0 2240 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_88
timestamp 1677622389
transform -1 0 2288 0 1 3770
box -8 -3 46 105
use FILL  FILL_1947
timestamp 1677622389
transform 1 0 2288 0 1 3770
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1677622389
transform 1 0 2296 0 1 3770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1677622389
transform 1 0 2304 0 1 3770
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1677622389
transform 1 0 2312 0 1 3770
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1677622389
transform 1 0 2320 0 1 3770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1677622389
transform 1 0 2328 0 1 3770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1677622389
transform 1 0 2336 0 1 3770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1677622389
transform 1 0 2344 0 1 3770
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1677622389
transform 1 0 2352 0 1 3770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1677622389
transform 1 0 2360 0 1 3770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1677622389
transform 1 0 2368 0 1 3770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1677622389
transform 1 0 2376 0 1 3770
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1677622389
transform 1 0 2384 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1702
timestamp 1677622389
transform 1 0 2420 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_144
timestamp 1677622389
transform -1 0 2488 0 1 3770
box -8 -3 104 105
use FILL  FILL_1967
timestamp 1677622389
transform 1 0 2488 0 1 3770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1677622389
transform 1 0 2496 0 1 3770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1677622389
transform 1 0 2504 0 1 3770
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1677622389
transform 1 0 2512 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_95
timestamp 1677622389
transform 1 0 2520 0 1 3770
box -8 -3 46 105
use FILL  FILL_1982
timestamp 1677622389
transform 1 0 2560 0 1 3770
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1677622389
transform 1 0 2568 0 1 3770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1677622389
transform 1 0 2576 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_169
timestamp 1677622389
transform 1 0 2584 0 1 3770
box -9 -3 26 105
use FILL  FILL_1991
timestamp 1677622389
transform 1 0 2600 0 1 3770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1677622389
transform 1 0 2608 0 1 3770
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1677622389
transform 1 0 2616 0 1 3770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1677622389
transform 1 0 2624 0 1 3770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1677622389
transform 1 0 2632 0 1 3770
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1677622389
transform 1 0 2640 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1677622389
transform 1 0 2648 0 1 3770
box -8 -3 104 105
use FILL  FILL_2000
timestamp 1677622389
transform 1 0 2744 0 1 3770
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1677622389
transform 1 0 2752 0 1 3770
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1677622389
transform 1 0 2760 0 1 3770
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1677622389
transform 1 0 2768 0 1 3770
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1677622389
transform 1 0 2776 0 1 3770
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1677622389
transform 1 0 2784 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_23
timestamp 1677622389
transform 1 0 2792 0 1 3770
box -8 -3 32 105
use FILL  FILL_2006
timestamp 1677622389
transform 1 0 2816 0 1 3770
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1677622389
transform 1 0 2824 0 1 3770
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1677622389
transform 1 0 2832 0 1 3770
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1677622389
transform 1 0 2840 0 1 3770
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1677622389
transform 1 0 2848 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_49
timestamp 1677622389
transform 1 0 2856 0 1 3770
box -8 -3 34 105
use FILL  FILL_2017
timestamp 1677622389
transform 1 0 2888 0 1 3770
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1677622389
transform 1 0 2896 0 1 3770
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1677622389
transform 1 0 2904 0 1 3770
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1677622389
transform 1 0 2912 0 1 3770
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1677622389
transform 1 0 2920 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_50
timestamp 1677622389
transform -1 0 2960 0 1 3770
box -8 -3 34 105
use FILL  FILL_2022
timestamp 1677622389
transform 1 0 2960 0 1 3770
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1677622389
transform 1 0 2968 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1677622389
transform 1 0 2976 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_172
timestamp 1677622389
transform 1 0 3072 0 1 3770
box -9 -3 26 105
use FILL  FILL_2034
timestamp 1677622389
transform 1 0 3088 0 1 3770
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1677622389
transform 1 0 3096 0 1 3770
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1677622389
transform 1 0 3104 0 1 3770
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1677622389
transform 1 0 3112 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_90
timestamp 1677622389
transform -1 0 3160 0 1 3770
box -8 -3 46 105
use FILL  FILL_2038
timestamp 1677622389
transform 1 0 3160 0 1 3770
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1677622389
transform 1 0 3168 0 1 3770
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1677622389
transform 1 0 3176 0 1 3770
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1677622389
transform 1 0 3184 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1677622389
transform 1 0 3192 0 1 3770
box -8 -3 104 105
use FILL  FILL_2042
timestamp 1677622389
transform 1 0 3288 0 1 3770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1677622389
transform 1 0 3296 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_174
timestamp 1677622389
transform 1 0 3304 0 1 3770
box -9 -3 26 105
use FILL  FILL_2062
timestamp 1677622389
transform 1 0 3320 0 1 3770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1677622389
transform 1 0 3328 0 1 3770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1677622389
transform 1 0 3336 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1677622389
transform 1 0 3344 0 1 3770
box -8 -3 104 105
use FILL  FILL_2065
timestamp 1677622389
transform 1 0 3440 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_92
timestamp 1677622389
transform 1 0 3448 0 1 3770
box -8 -3 46 105
use FILL  FILL_2072
timestamp 1677622389
transform 1 0 3488 0 1 3770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1677622389
transform 1 0 3496 0 1 3770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1677622389
transform 1 0 3504 0 1 3770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1677622389
transform 1 0 3512 0 1 3770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1677622389
transform 1 0 3520 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_175
timestamp 1677622389
transform 1 0 3528 0 1 3770
box -9 -3 26 105
use FILL  FILL_2077
timestamp 1677622389
transform 1 0 3544 0 1 3770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1677622389
transform 1 0 3552 0 1 3770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1677622389
transform 1 0 3560 0 1 3770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1677622389
transform 1 0 3568 0 1 3770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1677622389
transform 1 0 3576 0 1 3770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1677622389
transform 1 0 3584 0 1 3770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1677622389
transform 1 0 3592 0 1 3770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1677622389
transform 1 0 3600 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_176
timestamp 1677622389
transform -1 0 3624 0 1 3770
box -9 -3 26 105
use M3_M2  M3_M2_1703
timestamp 1677622389
transform 1 0 3636 0 1 3775
box -3 -3 3 3
use FILL  FILL_2095
timestamp 1677622389
transform 1 0 3624 0 1 3770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1677622389
transform 1 0 3632 0 1 3770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1677622389
transform 1 0 3640 0 1 3770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1677622389
transform 1 0 3648 0 1 3770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1677622389
transform 1 0 3656 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1677622389
transform 1 0 3664 0 1 3770
box -8 -3 104 105
use FILL  FILL_2106
timestamp 1677622389
transform 1 0 3760 0 1 3770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1677622389
transform 1 0 3768 0 1 3770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1677622389
transform 1 0 3776 0 1 3770
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1677622389
transform 1 0 3784 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_99
timestamp 1677622389
transform 1 0 3792 0 1 3770
box -8 -3 46 105
use FILL  FILL_2121
timestamp 1677622389
transform 1 0 3832 0 1 3770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1677622389
transform 1 0 3840 0 1 3770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1677622389
transform 1 0 3848 0 1 3770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1677622389
transform 1 0 3856 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_95
timestamp 1677622389
transform 1 0 3864 0 1 3770
box -8 -3 46 105
use FILL  FILL_2130
timestamp 1677622389
transform 1 0 3904 0 1 3770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1677622389
transform 1 0 3912 0 1 3770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1677622389
transform 1 0 3920 0 1 3770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1677622389
transform 1 0 3928 0 1 3770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1677622389
transform 1 0 3936 0 1 3770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1677622389
transform 1 0 3944 0 1 3770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1677622389
transform 1 0 3952 0 1 3770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1677622389
transform 1 0 3960 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_179
timestamp 1677622389
transform -1 0 3984 0 1 3770
box -9 -3 26 105
use FILL  FILL_2139
timestamp 1677622389
transform 1 0 3984 0 1 3770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1677622389
transform 1 0 3992 0 1 3770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1677622389
transform 1 0 4000 0 1 3770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1677622389
transform 1 0 4008 0 1 3770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1677622389
transform 1 0 4016 0 1 3770
box -8 -3 16 105
use NAND3X1  NAND3X1_10
timestamp 1677622389
transform -1 0 4056 0 1 3770
box -8 -3 40 105
use FILL  FILL_2144
timestamp 1677622389
transform 1 0 4056 0 1 3770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1677622389
transform 1 0 4064 0 1 3770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1677622389
transform 1 0 4072 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_96
timestamp 1677622389
transform 1 0 4080 0 1 3770
box -8 -3 46 105
use FILL  FILL_2150
timestamp 1677622389
transform 1 0 4120 0 1 3770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1677622389
transform 1 0 4128 0 1 3770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1677622389
transform 1 0 4136 0 1 3770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1677622389
transform 1 0 4144 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_100
timestamp 1677622389
transform 1 0 4152 0 1 3770
box -8 -3 46 105
use FILL  FILL_2154
timestamp 1677622389
transform 1 0 4192 0 1 3770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1677622389
transform 1 0 4200 0 1 3770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1677622389
transform 1 0 4208 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1677622389
transform 1 0 4216 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_180
timestamp 1677622389
transform 1 0 4312 0 1 3770
box -9 -3 26 105
use FILL  FILL_2157
timestamp 1677622389
transform 1 0 4328 0 1 3770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1677622389
transform 1 0 4336 0 1 3770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1677622389
transform 1 0 4344 0 1 3770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1677622389
transform 1 0 4352 0 1 3770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1677622389
transform 1 0 4360 0 1 3770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1677622389
transform 1 0 4368 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1704
timestamp 1677622389
transform 1 0 4412 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_99
timestamp 1677622389
transform 1 0 4376 0 1 3770
box -8 -3 46 105
use FILL  FILL_2180
timestamp 1677622389
transform 1 0 4416 0 1 3770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1677622389
transform 1 0 4424 0 1 3770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1677622389
transform 1 0 4432 0 1 3770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1677622389
transform 1 0 4440 0 1 3770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1677622389
transform 1 0 4448 0 1 3770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1677622389
transform 1 0 4456 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_183
timestamp 1677622389
transform 1 0 4464 0 1 3770
box -9 -3 26 105
use FILL  FILL_2186
timestamp 1677622389
transform 1 0 4480 0 1 3770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1677622389
transform 1 0 4488 0 1 3770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1677622389
transform 1 0 4496 0 1 3770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1677622389
transform 1 0 4504 0 1 3770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1677622389
transform 1 0 4512 0 1 3770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1677622389
transform 1 0 4520 0 1 3770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1677622389
transform 1 0 4528 0 1 3770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1677622389
transform 1 0 4536 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1677622389
transform 1 0 4544 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_184
timestamp 1677622389
transform 1 0 4640 0 1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_100
timestamp 1677622389
transform 1 0 4656 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1677622389
transform 1 0 4696 0 1 3770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_19
timestamp 1677622389
transform 1 0 4819 0 1 3770
box -10 -3 10 3
use M3_M2  M3_M2_1740
timestamp 1677622389
transform 1 0 156 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2010
timestamp 1677622389
transform 1 0 84 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1677622389
transform 1 0 108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1677622389
transform 1 0 172 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1705
timestamp 1677622389
transform 1 0 204 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1677622389
transform 1 0 236 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1677622389
transform 1 0 188 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2011
timestamp 1677622389
transform 1 0 188 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1677622389
transform 1 0 212 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1742
timestamp 1677622389
transform 1 0 284 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2012
timestamp 1677622389
transform 1 0 292 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1677622389
transform 1 0 284 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1728
timestamp 1677622389
transform 1 0 316 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1677622389
transform 1 0 332 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2013
timestamp 1677622389
transform 1 0 316 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1677622389
transform 1 0 332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1677622389
transform 1 0 308 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1677622389
transform 1 0 324 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1744
timestamp 1677622389
transform 1 0 364 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1677622389
transform 1 0 404 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2015
timestamp 1677622389
transform 1 0 364 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1677622389
transform 1 0 412 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1677622389
transform 1 0 444 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1824
timestamp 1677622389
transform 1 0 412 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1677622389
transform 1 0 444 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2111
timestamp 1677622389
transform 1 0 460 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1825
timestamp 1677622389
transform 1 0 460 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2016
timestamp 1677622389
transform 1 0 508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1677622389
transform 1 0 516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1677622389
transform 1 0 500 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1677622389
transform 1 0 524 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1842
timestamp 1677622389
transform 1 0 516 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2018
timestamp 1677622389
transform 1 0 556 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1677622389
transform 1 0 548 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1677622389
transform 1 0 596 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1746
timestamp 1677622389
transform 1 0 684 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2020
timestamp 1677622389
transform 1 0 684 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1677622389
transform 1 0 708 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1677622389
transform 1 0 772 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1707
timestamp 1677622389
transform 1 0 804 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2021
timestamp 1677622389
transform 1 0 812 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1791
timestamp 1677622389
transform 1 0 836 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2117
timestamp 1677622389
transform 1 0 836 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1677622389
transform 1 0 892 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1843
timestamp 1677622389
transform 1 0 844 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1677622389
transform 1 0 884 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1677622389
transform 1 0 916 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2022
timestamp 1677622389
transform 1 0 948 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1729
timestamp 1677622389
transform 1 0 964 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2007
timestamp 1677622389
transform 1 0 964 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1677622389
transform 1 0 956 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1677622389
transform 1 0 1004 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1677622389
transform 1 0 1012 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1708
timestamp 1677622389
transform 1 0 1028 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2008
timestamp 1677622389
transform 1 0 1028 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1677622389
transform 1 0 1076 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1747
timestamp 1677622389
transform 1 0 1092 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2121
timestamp 1677622389
transform 1 0 1092 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1677622389
transform 1 0 1108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1677622389
transform 1 0 1124 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1748
timestamp 1677622389
transform 1 0 1148 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2026
timestamp 1677622389
transform 1 0 1148 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1709
timestamp 1677622389
transform 1 0 1196 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2207
timestamp 1677622389
transform 1 0 1196 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1710
timestamp 1677622389
transform 1 0 1212 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1677622389
transform 1 0 1220 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1711
timestamp 1677622389
transform 1 0 1252 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1677622389
transform 1 0 1244 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1677622389
transform 1 0 1252 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2027
timestamp 1677622389
transform 1 0 1252 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1677622389
transform 1 0 1244 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1864
timestamp 1677622389
transform 1 0 1268 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2125
timestamp 1677622389
transform 1 0 1292 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1677622389
transform 1 0 1300 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1731
timestamp 1677622389
transform 1 0 1356 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1677622389
transform 1 0 1380 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1677622389
transform 1 0 1396 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2028
timestamp 1677622389
transform 1 0 1420 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1677622389
transform 1 0 1340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1812
timestamp 1677622389
transform 1 0 1380 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2128
timestamp 1677622389
transform 1 0 1396 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1826
timestamp 1677622389
transform 1 0 1420 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1677622389
transform 1 0 1396 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1677622389
transform 1 0 1436 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1677622389
transform 1 0 1468 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1677622389
transform 1 0 1484 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2029
timestamp 1677622389
transform 1 0 1468 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1677622389
transform 1 0 1484 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1813
timestamp 1677622389
transform 1 0 1468 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2129
timestamp 1677622389
transform 1 0 1476 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1827
timestamp 1677622389
transform 1 0 1500 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2130
timestamp 1677622389
transform 1 0 1516 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1828
timestamp 1677622389
transform 1 0 1516 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1677622389
transform 1 0 1548 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1677622389
transform 1 0 1540 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1677622389
transform 1 0 1532 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1677622389
transform 1 0 1572 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2031
timestamp 1677622389
transform 1 0 1532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1677622389
transform 1 0 1540 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1677622389
transform 1 0 1556 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1814
timestamp 1677622389
transform 1 0 1532 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2131
timestamp 1677622389
transform 1 0 1548 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1677622389
transform 1 0 1564 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1829
timestamp 1677622389
transform 1 0 1564 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2034
timestamp 1677622389
transform 1 0 1612 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1677622389
transform 1 0 1620 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1830
timestamp 1677622389
transform 1 0 1612 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2133
timestamp 1677622389
transform 1 0 1652 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1865
timestamp 1677622389
transform 1 0 1652 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1677622389
transform 1 0 1668 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1677622389
transform 1 0 1780 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1677622389
transform 1 0 1692 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1677622389
transform 1 0 1716 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1677622389
transform 1 0 1788 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2036
timestamp 1677622389
transform 1 0 1692 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1792
timestamp 1677622389
transform 1 0 1772 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2037
timestamp 1677622389
transform 1 0 1788 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1677622389
transform 1 0 1732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1677622389
transform 1 0 1772 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1677622389
transform 1 0 1780 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1831
timestamp 1677622389
transform 1 0 1780 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1677622389
transform 1 0 1828 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1677622389
transform 1 0 1820 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1677622389
transform 1 0 1828 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2137
timestamp 1677622389
transform 1 0 1908 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1794
timestamp 1677622389
transform 1 0 1924 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1677622389
transform 1 0 1964 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2038
timestamp 1677622389
transform 1 0 1964 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1715
timestamp 1677622389
transform 1 0 1988 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2138
timestamp 1677622389
transform 1 0 1988 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1677622389
transform 1 0 1996 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1846
timestamp 1677622389
transform 1 0 1996 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2139
timestamp 1677622389
transform 1 0 2012 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1832
timestamp 1677622389
transform 1 0 2012 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1677622389
transform 1 0 2028 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1677622389
transform 1 0 2044 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2040
timestamp 1677622389
transform 1 0 2036 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1718
timestamp 1677622389
transform 1 0 2100 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1677622389
transform 1 0 2092 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2041
timestamp 1677622389
transform 1 0 2068 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1677622389
transform 1 0 2092 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1677622389
transform 1 0 2100 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1815
timestamp 1677622389
transform 1 0 2076 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2140
timestamp 1677622389
transform 1 0 2084 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1795
timestamp 1677622389
transform 1 0 2108 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2141
timestamp 1677622389
transform 1 0 2108 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1847
timestamp 1677622389
transform 1 0 2084 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1677622389
transform 1 0 2100 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1677622389
transform 1 0 2084 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2044
timestamp 1677622389
transform 1 0 2132 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1761
timestamp 1677622389
transform 1 0 2172 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2045
timestamp 1677622389
transform 1 0 2156 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1796
timestamp 1677622389
transform 1 0 2164 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2046
timestamp 1677622389
transform 1 0 2172 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1816
timestamp 1677622389
transform 1 0 2156 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2142
timestamp 1677622389
transform 1 0 2164 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1719
timestamp 1677622389
transform 1 0 2188 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2143
timestamp 1677622389
transform 1 0 2212 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1859
timestamp 1677622389
transform 1 0 2212 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1677622389
transform 1 0 2244 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1677622389
transform 1 0 2228 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2047
timestamp 1677622389
transform 1 0 2228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1677622389
transform 1 0 2244 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1677622389
transform 1 0 2236 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1677622389
transform 1 0 2252 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1763
timestamp 1677622389
transform 1 0 2292 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2146
timestamp 1677622389
transform 1 0 2284 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1721
timestamp 1677622389
transform 1 0 2316 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2049
timestamp 1677622389
transform 1 0 2316 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1817
timestamp 1677622389
transform 1 0 2316 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2147
timestamp 1677622389
transform 1 0 2324 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1677622389
transform 1 0 2340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1849
timestamp 1677622389
transform 1 0 2340 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1677622389
transform 1 0 2380 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2050
timestamp 1677622389
transform 1 0 2372 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1677622389
transform 1 0 2388 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1677622389
transform 1 0 2380 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1860
timestamp 1677622389
transform 1 0 2372 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1677622389
transform 1 0 2404 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2052
timestamp 1677622389
transform 1 0 2404 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1797
timestamp 1677622389
transform 1 0 2412 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1677622389
transform 1 0 2428 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2150
timestamp 1677622389
transform 1 0 2428 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1850
timestamp 1677622389
transform 1 0 2428 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2151
timestamp 1677622389
transform 1 0 2444 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1677622389
transform 1 0 2460 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1851
timestamp 1677622389
transform 1 0 2460 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1677622389
transform 1 0 2492 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1677622389
transform 1 0 2508 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1677622389
transform 1 0 2524 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2053
timestamp 1677622389
transform 1 0 2508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1677622389
transform 1 0 2516 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1800
timestamp 1677622389
transform 1 0 2564 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2154
timestamp 1677622389
transform 1 0 2564 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1768
timestamp 1677622389
transform 1 0 2580 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1677622389
transform 1 0 2604 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1677622389
transform 1 0 2620 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2054
timestamp 1677622389
transform 1 0 2596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1677622389
transform 1 0 2604 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1677622389
transform 1 0 2588 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1818
timestamp 1677622389
transform 1 0 2596 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1677622389
transform 1 0 2636 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2056
timestamp 1677622389
transform 1 0 2644 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1677622389
transform 1 0 2604 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1677622389
transform 1 0 2620 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1677622389
transform 1 0 2636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1861
timestamp 1677622389
transform 1 0 2588 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2159
timestamp 1677622389
transform 1 0 2652 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1852
timestamp 1677622389
transform 1 0 2644 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1677622389
transform 1 0 2684 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2057
timestamp 1677622389
transform 1 0 2676 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1677622389
transform 1 0 2684 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1819
timestamp 1677622389
transform 1 0 2668 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1677622389
transform 1 0 2660 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1677622389
transform 1 0 2652 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1677622389
transform 1 0 2716 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1677622389
transform 1 0 2756 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2059
timestamp 1677622389
transform 1 0 2804 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1677622389
transform 1 0 2716 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1677622389
transform 1 0 2724 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1820
timestamp 1677622389
transform 1 0 2732 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2162
timestamp 1677622389
transform 1 0 2756 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1853
timestamp 1677622389
transform 1 0 2724 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1677622389
transform 1 0 2740 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1677622389
transform 1 0 2820 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2009
timestamp 1677622389
transform 1 0 2820 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1677622389
transform 1 0 2836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1677622389
transform 1 0 2868 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1677622389
transform 1 0 2884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1677622389
transform 1 0 2916 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1677622389
transform 1 0 2924 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1855
timestamp 1677622389
transform 1 0 2924 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2063
timestamp 1677622389
transform 1 0 2956 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1821
timestamp 1677622389
transform 1 0 2956 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2164
timestamp 1677622389
transform 1 0 2964 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1677622389
transform 1 0 2972 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1856
timestamp 1677622389
transform 1 0 2972 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2165
timestamp 1677622389
transform 1 0 3004 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1677622389
transform 1 0 3020 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1804
timestamp 1677622389
transform 1 0 3036 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1677622389
transform 1 0 3076 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2064
timestamp 1677622389
transform 1 0 3076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1677622389
transform 1 0 3084 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1735
timestamp 1677622389
transform 1 0 3124 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1677622389
transform 1 0 3132 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2066
timestamp 1677622389
transform 1 0 3100 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1805
timestamp 1677622389
transform 1 0 3108 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2067
timestamp 1677622389
transform 1 0 3116 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1677622389
transform 1 0 3132 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1677622389
transform 1 0 3108 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1833
timestamp 1677622389
transform 1 0 3124 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2168
timestamp 1677622389
transform 1 0 3148 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1677622389
transform 1 0 3172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1677622389
transform 1 0 3196 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1677622389
transform 1 0 3284 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1774
timestamp 1677622389
transform 1 0 3316 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1677622389
transform 1 0 3356 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2070
timestamp 1677622389
transform 1 0 3316 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1677622389
transform 1 0 3364 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1677622389
transform 1 0 3396 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1834
timestamp 1677622389
transform 1 0 3364 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2173
timestamp 1677622389
transform 1 0 3412 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1723
timestamp 1677622389
transform 1 0 3452 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2071
timestamp 1677622389
transform 1 0 3476 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1835
timestamp 1677622389
transform 1 0 3468 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1677622389
transform 1 0 3508 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1677622389
transform 1 0 3524 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1724
timestamp 1677622389
transform 1 0 3572 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1677622389
transform 1 0 3564 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1677622389
transform 1 0 3596 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1677622389
transform 1 0 3564 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1677622389
transform 1 0 3572 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1677622389
transform 1 0 3588 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1677622389
transform 1 0 3556 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1677622389
transform 1 0 3572 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1677622389
transform 1 0 3596 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1677622389
transform 1 0 3612 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1677622389
transform 1 0 3620 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1725
timestamp 1677622389
transform 1 0 3676 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1677622389
transform 1 0 3724 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2076
timestamp 1677622389
transform 1 0 3716 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1677622389
transform 1 0 3724 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1779
timestamp 1677622389
transform 1 0 3756 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1677622389
transform 1 0 3788 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1677622389
transform 1 0 3828 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2078
timestamp 1677622389
transform 1 0 3788 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1677622389
transform 1 0 3804 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1677622389
transform 1 0 3820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1677622389
transform 1 0 3780 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1677622389
transform 1 0 3796 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1677622389
transform 1 0 3820 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1677622389
transform 1 0 3836 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1726
timestamp 1677622389
transform 1 0 3940 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1677622389
transform 1 0 3900 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2081
timestamp 1677622389
transform 1 0 3868 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1677622389
transform 1 0 3892 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1677622389
transform 1 0 3948 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1727
timestamp 1677622389
transform 1 0 3972 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1677622389
transform 1 0 4020 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2082
timestamp 1677622389
transform 1 0 3972 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1677622389
transform 1 0 4020 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1822
timestamp 1677622389
transform 1 0 4044 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1677622389
transform 1 0 4092 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1677622389
transform 1 0 4116 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1677622389
transform 1 0 4132 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2083
timestamp 1677622389
transform 1 0 4116 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1807
timestamp 1677622389
transform 1 0 4124 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2084
timestamp 1677622389
transform 1 0 4132 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1677622389
transform 1 0 4148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1677622389
transform 1 0 4116 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1677622389
transform 1 0 4124 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1677622389
transform 1 0 4140 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1836
timestamp 1677622389
transform 1 0 4116 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1677622389
transform 1 0 4140 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2190
timestamp 1677622389
transform 1 0 4156 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1677622389
transform 1 0 4196 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1808
timestamp 1677622389
transform 1 0 4204 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1677622389
transform 1 0 4228 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2087
timestamp 1677622389
transform 1 0 4212 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1677622389
transform 1 0 4220 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1677622389
transform 1 0 4228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1677622389
transform 1 0 4204 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1838
timestamp 1677622389
transform 1 0 4212 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1677622389
transform 1 0 4244 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1677622389
transform 1 0 4268 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1677622389
transform 1 0 4284 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2090
timestamp 1677622389
transform 1 0 4268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1677622389
transform 1 0 4284 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1677622389
transform 1 0 4260 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1809
timestamp 1677622389
transform 1 0 4292 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2193
timestamp 1677622389
transform 1 0 4292 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1839
timestamp 1677622389
transform 1 0 4268 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2092
timestamp 1677622389
transform 1 0 4316 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1677622389
transform 1 0 4308 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1840
timestamp 1677622389
transform 1 0 4324 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1677622389
transform 1 0 4364 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2093
timestamp 1677622389
transform 1 0 4364 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1739
timestamp 1677622389
transform 1 0 4460 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1677622389
transform 1 0 4404 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2094
timestamp 1677622389
transform 1 0 4380 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1677622389
transform 1 0 4404 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1677622389
transform 1 0 4460 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1677622389
transform 1 0 4476 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1677622389
transform 1 0 4508 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1810
timestamp 1677622389
transform 1 0 4516 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2096
timestamp 1677622389
transform 1 0 4532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1677622389
transform 1 0 4548 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1823
timestamp 1677622389
transform 1 0 4508 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2198
timestamp 1677622389
transform 1 0 4516 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1677622389
transform 1 0 4532 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1677622389
transform 1 0 4572 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1677622389
transform 1 0 4636 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1677622389
transform 1 0 4636 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1677622389
transform 1 0 4652 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1789
timestamp 1677622389
transform 1 0 4676 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1677622389
transform 1 0 4700 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2099
timestamp 1677622389
transform 1 0 4684 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1811
timestamp 1677622389
transform 1 0 4692 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2100
timestamp 1677622389
transform 1 0 4700 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1677622389
transform 1 0 4668 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1677622389
transform 1 0 4692 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1677622389
transform 1 0 4708 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1677622389
transform 1 0 4740 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1677622389
transform 1 0 4756 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1677622389
transform 1 0 4780 0 1 3735
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_20
timestamp 1677622389
transform 1 0 24 0 1 3670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_130
timestamp 1677622389
transform 1 0 72 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1734
timestamp 1677622389
transform 1 0 168 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1867
timestamp 1677622389
transform 1 0 196 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_132
timestamp 1677622389
transform 1 0 176 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1748
timestamp 1677622389
transform 1 0 272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1677622389
transform 1 0 280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1677622389
transform 1 0 288 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_81
timestamp 1677622389
transform 1 0 296 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1751
timestamp 1677622389
transform 1 0 336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1677622389
transform 1 0 344 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1677622389
transform 1 0 352 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1753
timestamp 1677622389
transform 1 0 448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1677622389
transform 1 0 456 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_153
timestamp 1677622389
transform -1 0 480 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1755
timestamp 1677622389
transform 1 0 480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1677622389
transform 1 0 488 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1677622389
transform 1 0 496 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_87
timestamp 1677622389
transform -1 0 544 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1765
timestamp 1677622389
transform 1 0 544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1677622389
transform 1 0 552 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1677622389
transform 1 0 560 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1677622389
transform 1 0 568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1677622389
transform 1 0 576 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1677622389
transform 1 0 584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1677622389
transform 1 0 592 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1677622389
transform 1 0 600 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1677622389
transform 1 0 608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1677622389
transform 1 0 616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1677622389
transform 1 0 624 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1677622389
transform 1 0 632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1677622389
transform 1 0 640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1677622389
transform 1 0 648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1677622389
transform 1 0 656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1677622389
transform 1 0 664 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1677622389
transform 1 0 672 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1792
timestamp 1677622389
transform 1 0 768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1677622389
transform 1 0 776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1677622389
transform 1 0 784 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1677622389
transform 1 0 792 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1868
timestamp 1677622389
transform 1 0 844 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_136
timestamp 1677622389
transform 1 0 800 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1802
timestamp 1677622389
transform 1 0 896 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1677622389
transform 1 0 904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1677622389
transform 1 0 912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1677622389
transform 1 0 920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1677622389
transform 1 0 928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1677622389
transform 1 0 936 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_155
timestamp 1677622389
transform 1 0 944 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1811
timestamp 1677622389
transform 1 0 960 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1677622389
transform 1 0 968 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1677622389
transform 1 0 976 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1677622389
transform 1 0 984 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_21
timestamp 1677622389
transform 1 0 992 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1818
timestamp 1677622389
transform 1 0 1016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1677622389
transform 1 0 1024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1677622389
transform 1 0 1032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1677622389
transform 1 0 1040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1677622389
transform 1 0 1048 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_22
timestamp 1677622389
transform 1 0 1056 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1825
timestamp 1677622389
transform 1 0 1080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1677622389
transform 1 0 1088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1677622389
transform 1 0 1096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1677622389
transform 1 0 1104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1677622389
transform 1 0 1112 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_44
timestamp 1677622389
transform 1 0 1120 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1830
timestamp 1677622389
transform 1 0 1152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1677622389
transform 1 0 1160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1677622389
transform 1 0 1168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1677622389
transform 1 0 1176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1677622389
transform 1 0 1184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1677622389
transform 1 0 1192 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_46
timestamp 1677622389
transform -1 0 1232 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1839
timestamp 1677622389
transform 1 0 1232 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1677622389
transform 1 0 1240 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1677622389
transform 1 0 1248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1677622389
transform 1 0 1256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1677622389
transform 1 0 1264 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_157
timestamp 1677622389
transform 1 0 1272 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1677622389
transform 1 0 1288 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1849
timestamp 1677622389
transform 1 0 1304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1677622389
transform 1 0 1312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1677622389
transform 1 0 1320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1677622389
transform 1 0 1328 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_138
timestamp 1677622389
transform -1 0 1432 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1862
timestamp 1677622389
transform 1 0 1432 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1677622389
transform 1 0 1440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1677622389
transform 1 0 1448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1677622389
transform 1 0 1456 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_84
timestamp 1677622389
transform -1 0 1504 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1873
timestamp 1677622389
transform 1 0 1504 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1677622389
transform 1 0 1512 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1677622389
transform 1 0 1520 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1677622389
transform 1 0 1528 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_85
timestamp 1677622389
transform -1 0 1576 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1877
timestamp 1677622389
transform 1 0 1576 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1677622389
transform 1 0 1584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1677622389
transform 1 0 1592 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1677622389
transform 1 0 1600 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1677622389
transform 1 0 1608 0 -1 3770
box -8 -3 16 105
use BUFX2  BUFX2_12
timestamp 1677622389
transform -1 0 1640 0 -1 3770
box -5 -3 28 105
use FILL  FILL_1882
timestamp 1677622389
transform 1 0 1640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1677622389
transform 1 0 1648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1677622389
transform 1 0 1656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1677622389
transform 1 0 1664 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1677622389
transform 1 0 1672 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1869
timestamp 1677622389
transform 1 0 1740 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_141
timestamp 1677622389
transform 1 0 1680 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_162
timestamp 1677622389
transform -1 0 1792 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1892
timestamp 1677622389
transform 1 0 1792 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1677622389
transform 1 0 1800 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1677622389
transform 1 0 1808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1677622389
transform 1 0 1816 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1677622389
transform 1 0 1824 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1677622389
transform 1 0 1832 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1677622389
transform 1 0 1840 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1677622389
transform 1 0 1848 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1677622389
transform 1 0 1856 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1677622389
transform 1 0 1864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1677622389
transform 1 0 1872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1677622389
transform 1 0 1880 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1677622389
transform 1 0 1888 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1677622389
transform 1 0 1896 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1677622389
transform 1 0 1904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1677622389
transform 1 0 1912 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_164
timestamp 1677622389
transform -1 0 1936 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1916
timestamp 1677622389
transform 1 0 1936 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1677622389
transform 1 0 1944 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1870
timestamp 1677622389
transform 1 0 1964 0 1 3675
box -3 -3 3 3
use FILL  FILL_1918
timestamp 1677622389
transform 1 0 1952 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1677622389
transform 1 0 1960 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_165
timestamp 1677622389
transform -1 0 1984 0 -1 3770
box -9 -3 26 105
use M3_M2  M3_M2_1871
timestamp 1677622389
transform 1 0 1996 0 1 3675
box -3 -3 3 3
use FILL  FILL_1924
timestamp 1677622389
transform 1 0 1984 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1677622389
transform 1 0 1992 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1677622389
transform 1 0 2000 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_167
timestamp 1677622389
transform -1 0 2024 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1929
timestamp 1677622389
transform 1 0 2024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1677622389
transform 1 0 2032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1677622389
transform 1 0 2040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1677622389
transform 1 0 2048 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1677622389
transform 1 0 2056 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_92
timestamp 1677622389
transform 1 0 2064 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1934
timestamp 1677622389
transform 1 0 2104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1677622389
transform 1 0 2112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1677622389
transform 1 0 2120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1677622389
transform 1 0 2128 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_87
timestamp 1677622389
transform 1 0 2136 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1938
timestamp 1677622389
transform 1 0 2176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1677622389
transform 1 0 2184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1677622389
transform 1 0 2192 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1677622389
transform 1 0 2200 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1677622389
transform 1 0 2208 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1872
timestamp 1677622389
transform 1 0 2244 0 1 3675
box -3 -3 3 3
use AOI22X1  AOI22X1_93
timestamp 1677622389
transform 1 0 2216 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1948
timestamp 1677622389
transform 1 0 2256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1677622389
transform 1 0 2264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1677622389
transform 1 0 2272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1677622389
transform 1 0 2280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1677622389
transform 1 0 2288 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_89
timestamp 1677622389
transform 1 0 2296 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1959
timestamp 1677622389
transform 1 0 2336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1677622389
transform 1 0 2344 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1873
timestamp 1677622389
transform 1 0 2364 0 1 3675
box -3 -3 3 3
use FILL  FILL_1968
timestamp 1677622389
transform 1 0 2352 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_94
timestamp 1677622389
transform -1 0 2400 0 -1 3770
box -8 -3 46 105
use M3_M2  M3_M2_1874
timestamp 1677622389
transform 1 0 2412 0 1 3675
box -3 -3 3 3
use FILL  FILL_1969
timestamp 1677622389
transform 1 0 2400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1677622389
transform 1 0 2408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1677622389
transform 1 0 2416 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_168
timestamp 1677622389
transform 1 0 2424 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1972
timestamp 1677622389
transform 1 0 2440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1677622389
transform 1 0 2448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1677622389
transform 1 0 2456 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1677622389
transform 1 0 2464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1677622389
transform 1 0 2472 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1677622389
transform 1 0 2480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1677622389
transform 1 0 2488 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_96
timestamp 1677622389
transform 1 0 2496 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1983
timestamp 1677622389
transform 1 0 2536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1677622389
transform 1 0 2544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1677622389
transform 1 0 2552 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1677622389
transform 1 0 2560 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1677622389
transform 1 0 2568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1677622389
transform 1 0 2576 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1677622389
transform 1 0 2584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1677622389
transform 1 0 2592 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_97
timestamp 1677622389
transform 1 0 2600 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1999
timestamp 1677622389
transform 1 0 2640 0 -1 3770
box -8 -3 16 105
use BUFX2  BUFX2_13
timestamp 1677622389
transform 1 0 2648 0 -1 3770
box -5 -3 28 105
use FILL  FILL_2007
timestamp 1677622389
transform 1 0 2672 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1677622389
transform 1 0 2680 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_170
timestamp 1677622389
transform 1 0 2688 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2009
timestamp 1677622389
transform 1 0 2704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1677622389
transform 1 0 2712 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1875
timestamp 1677622389
transform 1 0 2748 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_146
timestamp 1677622389
transform -1 0 2816 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2011
timestamp 1677622389
transform 1 0 2816 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_24
timestamp 1677622389
transform 1 0 2824 0 -1 3770
box -8 -3 32 105
use FILL  FILL_2016
timestamp 1677622389
transform 1 0 2848 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1677622389
transform 1 0 2856 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1677622389
transform 1 0 2864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1677622389
transform 1 0 2872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1677622389
transform 1 0 2880 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1677622389
transform 1 0 2888 0 -1 3770
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1677622389
transform -1 0 2920 0 -1 3770
box -8 -3 32 105
use FILL  FILL_2028
timestamp 1677622389
transform 1 0 2920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1677622389
transform 1 0 2928 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1876
timestamp 1677622389
transform 1 0 2964 0 1 3675
box -3 -3 3 3
use INVX2  INVX2_171
timestamp 1677622389
transform 1 0 2936 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2030
timestamp 1677622389
transform 1 0 2952 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1677622389
transform 1 0 2960 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1677622389
transform 1 0 2968 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1677622389
transform 1 0 2976 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1677622389
transform 1 0 2984 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1677622389
transform 1 0 2992 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1877
timestamp 1677622389
transform 1 0 3028 0 1 3675
box -3 -3 3 3
use OAI21X1  OAI21X1_51
timestamp 1677622389
transform -1 0 3032 0 -1 3770
box -8 -3 34 105
use FILL  FILL_2046
timestamp 1677622389
transform 1 0 3032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1677622389
transform 1 0 3040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1677622389
transform 1 0 3048 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1677622389
transform 1 0 3056 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1677622389
transform 1 0 3064 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1677622389
transform 1 0 3072 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1677622389
transform 1 0 3080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1677622389
transform 1 0 3088 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_91
timestamp 1677622389
transform -1 0 3136 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2054
timestamp 1677622389
transform 1 0 3136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1677622389
transform 1 0 3144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1677622389
transform 1 0 3152 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1878
timestamp 1677622389
transform 1 0 3180 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_149
timestamp 1677622389
transform 1 0 3160 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2057
timestamp 1677622389
transform 1 0 3256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1677622389
transform 1 0 3264 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1879
timestamp 1677622389
transform 1 0 3284 0 1 3675
box -3 -3 3 3
use INVX2  INVX2_173
timestamp 1677622389
transform 1 0 3272 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2059
timestamp 1677622389
transform 1 0 3288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1677622389
transform 1 0 3296 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_151
timestamp 1677622389
transform 1 0 3304 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2066
timestamp 1677622389
transform 1 0 3400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1677622389
transform 1 0 3408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1677622389
transform 1 0 3416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1677622389
transform 1 0 3424 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1677622389
transform 1 0 3432 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1677622389
transform 1 0 3440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1677622389
transform 1 0 3448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1677622389
transform 1 0 3456 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1677622389
transform 1 0 3464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1677622389
transform 1 0 3472 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1677622389
transform 1 0 3480 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_98
timestamp 1677622389
transform 1 0 3488 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2083
timestamp 1677622389
transform 1 0 3528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1677622389
transform 1 0 3536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1677622389
transform 1 0 3544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1677622389
transform 1 0 3552 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1677622389
transform 1 0 3560 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_93
timestamp 1677622389
transform 1 0 3568 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2096
timestamp 1677622389
transform 1 0 3608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1677622389
transform 1 0 3616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1677622389
transform 1 0 3624 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1677622389
transform 1 0 3632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1677622389
transform 1 0 3640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1677622389
transform 1 0 3648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1677622389
transform 1 0 3656 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_177
timestamp 1677622389
transform -1 0 3680 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2108
timestamp 1677622389
transform 1 0 3680 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1677622389
transform 1 0 3688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1677622389
transform 1 0 3696 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1677622389
transform 1 0 3704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1677622389
transform 1 0 3712 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_178
timestamp 1677622389
transform 1 0 3720 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2113
timestamp 1677622389
transform 1 0 3736 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1677622389
transform 1 0 3744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1677622389
transform 1 0 3752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1677622389
transform 1 0 3760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1677622389
transform 1 0 3768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1677622389
transform 1 0 3776 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_94
timestamp 1677622389
transform -1 0 3824 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2123
timestamp 1677622389
transform 1 0 3824 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1677622389
transform 1 0 3832 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1677622389
transform 1 0 3840 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1677622389
transform 1 0 3848 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_153
timestamp 1677622389
transform 1 0 3856 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2137
timestamp 1677622389
transform 1 0 3952 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_154
timestamp 1677622389
transform 1 0 3960 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2145
timestamp 1677622389
transform 1 0 4056 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1677622389
transform 1 0 4064 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1677622389
transform 1 0 4072 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_181
timestamp 1677622389
transform 1 0 4080 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2159
timestamp 1677622389
transform 1 0 4096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1677622389
transform 1 0 4104 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_97
timestamp 1677622389
transform 1 0 4112 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2161
timestamp 1677622389
transform 1 0 4152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1677622389
transform 1 0 4160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1677622389
transform 1 0 4168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1677622389
transform 1 0 4176 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_101
timestamp 1677622389
transform 1 0 4184 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2165
timestamp 1677622389
transform 1 0 4224 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1677622389
transform 1 0 4232 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1677622389
transform 1 0 4240 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1677622389
transform 1 0 4248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1677622389
transform 1 0 4256 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_98
timestamp 1677622389
transform 1 0 4264 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2170
timestamp 1677622389
transform 1 0 4304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1677622389
transform 1 0 4312 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_182
timestamp 1677622389
transform -1 0 4336 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2172
timestamp 1677622389
transform 1 0 4336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1677622389
transform 1 0 4344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1677622389
transform 1 0 4352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1677622389
transform 1 0 4360 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1677622389
transform 1 0 4368 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2187
timestamp 1677622389
transform 1 0 4464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1677622389
transform 1 0 4472 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1677622389
transform 1 0 4480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1677622389
transform 1 0 4488 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_102
timestamp 1677622389
transform 1 0 4496 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_159
timestamp 1677622389
transform 1 0 4536 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2198
timestamp 1677622389
transform 1 0 4632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1677622389
transform 1 0 4640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1677622389
transform 1 0 4648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1677622389
transform 1 0 4656 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_101
timestamp 1677622389
transform 1 0 4664 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2202
timestamp 1677622389
transform 1 0 4704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1677622389
transform 1 0 4712 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1677622389
transform 1 0 4720 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_185
timestamp 1677622389
transform -1 0 4744 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2205
timestamp 1677622389
transform 1 0 4744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1677622389
transform 1 0 4752 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_186
timestamp 1677622389
transform -1 0 4776 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2207
timestamp 1677622389
transform 1 0 4776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1677622389
transform 1 0 4784 0 -1 3770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_21
timestamp 1677622389
transform 1 0 4843 0 1 3670
box -10 -3 10 3
use M3_M2  M3_M2_1951
timestamp 1677622389
transform 1 0 140 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1677622389
transform 1 0 180 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1677622389
transform 1 0 92 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2228
timestamp 1677622389
transform 1 0 140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1677622389
transform 1 0 172 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1677622389
transform 1 0 180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1677622389
transform 1 0 92 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2035
timestamp 1677622389
transform 1 0 172 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2231
timestamp 1677622389
transform 1 0 196 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1900
timestamp 1677622389
transform 1 0 220 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2232
timestamp 1677622389
transform 1 0 228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1677622389
transform 1 0 212 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1677622389
transform 1 0 220 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1677622389
transform 1 0 236 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2036
timestamp 1677622389
transform 1 0 236 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1677622389
transform 1 0 252 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2233
timestamp 1677622389
transform 1 0 260 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2017
timestamp 1677622389
transform 1 0 260 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1677622389
transform 1 0 356 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1677622389
transform 1 0 276 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1677622389
transform 1 0 300 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1677622389
transform 1 0 364 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1677622389
transform 1 0 276 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2234
timestamp 1677622389
transform 1 0 300 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1677622389
transform 1 0 356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1677622389
transform 1 0 364 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1677622389
transform 1 0 372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1677622389
transform 1 0 276 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2037
timestamp 1677622389
transform 1 0 300 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1677622389
transform 1 0 372 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1677622389
transform 1 0 428 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1677622389
transform 1 0 412 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2238
timestamp 1677622389
transform 1 0 420 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1677622389
transform 1 0 404 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1677622389
transform 1 0 412 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1677622389
transform 1 0 428 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1957
timestamp 1677622389
transform 1 0 444 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2239
timestamp 1677622389
transform 1 0 444 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1888
timestamp 1677622389
transform 1 0 556 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1677622389
transform 1 0 540 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1677622389
transform 1 0 532 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1677622389
transform 1 0 508 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1677622389
transform 1 0 548 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1677622389
transform 1 0 460 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2240
timestamp 1677622389
transform 1 0 508 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1677622389
transform 1 0 540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1677622389
transform 1 0 548 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1677622389
transform 1 0 460 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2038
timestamp 1677622389
transform 1 0 460 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1677622389
transform 1 0 508 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2243
timestamp 1677622389
transform 1 0 588 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2040
timestamp 1677622389
transform 1 0 580 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1677622389
transform 1 0 612 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1677622389
transform 1 0 628 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2244
timestamp 1677622389
transform 1 0 620 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1677622389
transform 1 0 636 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1677622389
transform 1 0 604 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1677622389
transform 1 0 612 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1677622389
transform 1 0 628 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2041
timestamp 1677622389
transform 1 0 628 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2354
timestamp 1677622389
transform 1 0 668 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1677622389
transform 1 0 708 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1677622389
transform 1 0 748 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1904
timestamp 1677622389
transform 1 0 780 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2212
timestamp 1677622389
transform 1 0 764 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2019
timestamp 1677622389
transform 1 0 764 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2356
timestamp 1677622389
transform 1 0 804 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2061
timestamp 1677622389
transform 1 0 804 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1677622389
transform 1 0 828 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2247
timestamp 1677622389
transform 1 0 828 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1677622389
transform 1 0 836 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1677622389
transform 1 0 844 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1905
timestamp 1677622389
transform 1 0 876 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1677622389
transform 1 0 892 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1677622389
transform 1 0 868 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2250
timestamp 1677622389
transform 1 0 876 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1677622389
transform 1 0 892 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1677622389
transform 1 0 860 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1677622389
transform 1 0 868 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1677622389
transform 1 0 884 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2062
timestamp 1677622389
transform 1 0 884 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1677622389
transform 1 0 916 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1677622389
transform 1 0 908 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2252
timestamp 1677622389
transform 1 0 916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1677622389
transform 1 0 908 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1881
timestamp 1677622389
transform 1 0 940 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1677622389
transform 1 0 964 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2253
timestamp 1677622389
transform 1 0 948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1677622389
transform 1 0 964 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1882
timestamp 1677622389
transform 1 0 980 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2213
timestamp 1677622389
transform 1 0 980 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1677622389
transform 1 0 996 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1677622389
transform 1 0 1012 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1890
timestamp 1677622389
transform 1 0 1044 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1677622389
transform 1 0 1028 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2255
timestamp 1677622389
transform 1 0 1028 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1677622389
transform 1 0 1044 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1677622389
transform 1 0 1068 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1997
timestamp 1677622389
transform 1 0 1068 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1677622389
transform 1 0 1060 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1677622389
transform 1 0 1060 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1677622389
transform 1 0 1100 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1677622389
transform 1 0 1092 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2363
timestamp 1677622389
transform 1 0 1092 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1929
timestamp 1677622389
transform 1 0 1108 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1677622389
transform 1 0 1156 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1677622389
transform 1 0 1132 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2256
timestamp 1677622389
transform 1 0 1116 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1677622389
transform 1 0 1124 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1677622389
transform 1 0 1140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1677622389
transform 1 0 1156 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2021
timestamp 1677622389
transform 1 0 1124 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2364
timestamp 1677622389
transform 1 0 1132 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2022
timestamp 1677622389
transform 1 0 1140 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1677622389
transform 1 0 1140 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1677622389
transform 1 0 1172 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2365
timestamp 1677622389
transform 1 0 1180 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1930
timestamp 1677622389
transform 1 0 1196 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2216
timestamp 1677622389
transform 1 0 1196 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1677622389
transform 1 0 1196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2064
timestamp 1677622389
transform 1 0 1196 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2260
timestamp 1677622389
transform 1 0 1220 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1677622389
transform 1 0 1228 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1931
timestamp 1677622389
transform 1 0 1244 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2217
timestamp 1677622389
transform 1 0 1244 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1998
timestamp 1677622389
transform 1 0 1252 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2368
timestamp 1677622389
transform 1 0 1252 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1677622389
transform 1 0 1276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1677622389
transform 1 0 1292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1677622389
transform 1 0 1300 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1677622389
transform 1 0 1300 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1932
timestamp 1677622389
transform 1 0 1316 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2264
timestamp 1677622389
transform 1 0 1316 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2024
timestamp 1677622389
transform 1 0 1332 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2265
timestamp 1677622389
transform 1 0 1356 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2025
timestamp 1677622389
transform 1 0 1356 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1677622389
transform 1 0 1388 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2218
timestamp 1677622389
transform 1 0 1412 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1883
timestamp 1677622389
transform 1 0 1452 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2266
timestamp 1677622389
transform 1 0 1460 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2000
timestamp 1677622389
transform 1 0 1500 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1677622389
transform 1 0 1428 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1677622389
transform 1 0 1460 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2370
timestamp 1677622389
transform 1 0 1500 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2001
timestamp 1677622389
transform 1 0 1532 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2267
timestamp 1677622389
transform 1 0 1556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1677622389
transform 1 0 1612 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1677622389
transform 1 0 1532 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2043
timestamp 1677622389
transform 1 0 1580 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1677622389
transform 1 0 1524 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1677622389
transform 1 0 1556 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1677622389
transform 1 0 1636 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1677622389
transform 1 0 1628 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1677622389
transform 1 0 1684 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1677622389
transform 1 0 1732 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2269
timestamp 1677622389
transform 1 0 1636 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1677622389
transform 1 0 1684 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2003
timestamp 1677622389
transform 1 0 1716 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2271
timestamp 1677622389
transform 1 0 1732 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1677622389
transform 1 0 1716 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1934
timestamp 1677622389
transform 1 0 1780 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1677622389
transform 1 0 1796 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1677622389
transform 1 0 1788 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2272
timestamp 1677622389
transform 1 0 1788 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1677622389
transform 1 0 1804 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1677622389
transform 1 0 1788 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1677622389
transform 1 0 1796 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1677622389
transform 1 0 1812 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2067
timestamp 1677622389
transform 1 0 1812 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1677622389
transform 1 0 1836 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1677622389
transform 1 0 1836 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1677622389
transform 1 0 1828 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2044
timestamp 1677622389
transform 1 0 1828 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1677622389
transform 1 0 1844 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1677622389
transform 1 0 1892 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1677622389
transform 1 0 1940 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1677622389
transform 1 0 1924 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1677622389
transform 1 0 1956 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1677622389
transform 1 0 2060 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1677622389
transform 1 0 2004 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1677622389
transform 1 0 2052 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1677622389
transform 1 0 1996 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1677622389
transform 1 0 1876 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1677622389
transform 1 0 1900 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1677622389
transform 1 0 1956 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1677622389
transform 1 0 1988 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1677622389
transform 1 0 1876 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2275
timestamp 1677622389
transform 1 0 1908 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1677622389
transform 1 0 1956 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1677622389
transform 1 0 1964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1677622389
transform 1 0 1980 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1677622389
transform 1 0 1996 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1677622389
transform 1 0 1876 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1677622389
transform 1 0 1964 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1677622389
transform 1 0 1988 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2046
timestamp 1677622389
transform 1 0 1948 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1677622389
transform 1 0 1988 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1677622389
transform 1 0 1964 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1677622389
transform 1 0 2164 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1677622389
transform 1 0 2108 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1677622389
transform 1 0 2092 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1677622389
transform 1 0 2156 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2280
timestamp 1677622389
transform 1 0 2044 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1677622389
transform 1 0 2100 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1677622389
transform 1 0 2020 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2005
timestamp 1677622389
transform 1 0 2116 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2282
timestamp 1677622389
transform 1 0 2156 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1677622389
transform 1 0 2116 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1973
timestamp 1677622389
transform 1 0 2252 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2283
timestamp 1677622389
transform 1 0 2204 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1677622389
transform 1 0 2212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1677622389
transform 1 0 2228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1677622389
transform 1 0 2244 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1677622389
transform 1 0 2252 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1677622389
transform 1 0 2212 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1677622389
transform 1 0 2220 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1677622389
transform 1 0 2236 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2048
timestamp 1677622389
transform 1 0 2212 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1677622389
transform 1 0 2228 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1677622389
transform 1 0 2204 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1677622389
transform 1 0 2236 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1677622389
transform 1 0 2284 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1677622389
transform 1 0 2276 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2384
timestamp 1677622389
transform 1 0 2292 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2050
timestamp 1677622389
transform 1 0 2292 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2288
timestamp 1677622389
transform 1 0 2340 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1677622389
transform 1 0 2356 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2006
timestamp 1677622389
transform 1 0 2364 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2290
timestamp 1677622389
transform 1 0 2372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1677622389
transform 1 0 2348 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1885
timestamp 1677622389
transform 1 0 2388 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1677622389
transform 1 0 2388 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2386
timestamp 1677622389
transform 1 0 2380 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1677622389
transform 1 0 2388 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2071
timestamp 1677622389
transform 1 0 2388 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2291
timestamp 1677622389
transform 1 0 2436 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1677622389
transform 1 0 2516 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1940
timestamp 1677622389
transform 1 0 2540 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1677622389
transform 1 0 2572 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1677622389
transform 1 0 2572 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2292
timestamp 1677622389
transform 1 0 2572 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1975
timestamp 1677622389
transform 1 0 2620 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2293
timestamp 1677622389
transform 1 0 2620 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1677622389
transform 1 0 2668 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1677622389
transform 1 0 2588 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1677622389
transform 1 0 2708 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1677622389
transform 1 0 2732 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1677622389
transform 1 0 2732 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1677622389
transform 1 0 2748 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_1942
timestamp 1677622389
transform 1 0 2764 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2391
timestamp 1677622389
transform 1 0 2764 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1677622389
transform 1 0 2796 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1677622389
transform 1 0 2812 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1886
timestamp 1677622389
transform 1 0 2836 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1677622389
transform 1 0 2844 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2220
timestamp 1677622389
transform 1 0 2844 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2072
timestamp 1677622389
transform 1 0 2868 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1677622389
transform 1 0 2892 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1677622389
transform 1 0 2900 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1677622389
transform 1 0 2924 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2221
timestamp 1677622389
transform 1 0 2924 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1677622389
transform 1 0 2916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1677622389
transform 1 0 2900 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1677622389
transform 1 0 2908 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2051
timestamp 1677622389
transform 1 0 2908 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1677622389
transform 1 0 2948 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2297
timestamp 1677622389
transform 1 0 2940 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1677622389
transform 1 0 2924 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1677622389
transform 1 0 3012 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2009
timestamp 1677622389
transform 1 0 3052 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2299
timestamp 1677622389
transform 1 0 3060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1677622389
transform 1 0 2948 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1677622389
transform 1 0 2964 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2052
timestamp 1677622389
transform 1 0 2940 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1677622389
transform 1 0 2916 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1677622389
transform 1 0 2932 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1677622389
transform 1 0 3012 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2399
timestamp 1677622389
transform 1 0 3068 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1677622389
transform 1 0 3084 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1677622389
transform 1 0 3092 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1677622389
transform 1 0 3132 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2300
timestamp 1677622389
transform 1 0 3100 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1677622389
transform 1 0 3084 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2011
timestamp 1677622389
transform 1 0 3124 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1677622389
transform 1 0 3100 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2401
timestamp 1677622389
transform 1 0 3108 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1677622389
transform 1 0 3124 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1677622389
transform 1 0 3132 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1677622389
transform 1 0 3108 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1677622389
transform 1 0 3148 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2301
timestamp 1677622389
transform 1 0 3148 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1896
timestamp 1677622389
transform 1 0 3204 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1677622389
transform 1 0 3196 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1677622389
transform 1 0 3180 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2302
timestamp 1677622389
transform 1 0 3180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1677622389
transform 1 0 3196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1677622389
transform 1 0 3188 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1677622389
transform 1 0 3260 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2210
timestamp 1677622389
transform 1 0 3260 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1677622389
transform 1 0 3244 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1677622389
transform 1 0 3236 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2055
timestamp 1677622389
transform 1 0 3236 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1677622389
transform 1 0 3260 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2304
timestamp 1677622389
transform 1 0 3260 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1917
timestamp 1677622389
transform 1 0 3276 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2223
timestamp 1677622389
transform 1 0 3276 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1677622389
transform 1 0 3276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1677622389
transform 1 0 3340 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2056
timestamp 1677622389
transform 1 0 3364 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2406
timestamp 1677622389
transform 1 0 3396 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1677622389
transform 1 0 3420 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2029
timestamp 1677622389
transform 1 0 3420 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2407
timestamp 1677622389
transform 1 0 3428 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2012
timestamp 1677622389
transform 1 0 3452 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2308
timestamp 1677622389
transform 1 0 3460 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1677622389
transform 1 0 3476 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2030
timestamp 1677622389
transform 1 0 3460 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2408
timestamp 1677622389
transform 1 0 3468 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1677622389
transform 1 0 3492 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1979
timestamp 1677622389
transform 1 0 3508 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1677622389
transform 1 0 3508 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1677622389
transform 1 0 3524 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1677622389
transform 1 0 3572 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1677622389
transform 1 0 3588 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2310
timestamp 1677622389
transform 1 0 3572 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1677622389
transform 1 0 3596 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1677622389
transform 1 0 3588 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1677622389
transform 1 0 3604 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2076
timestamp 1677622389
transform 1 0 3604 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2412
timestamp 1677622389
transform 1 0 3620 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1981
timestamp 1677622389
transform 1 0 3676 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2312
timestamp 1677622389
transform 1 0 3676 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1677622389
transform 1 0 3732 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1677622389
transform 1 0 3652 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1677622389
transform 1 0 3748 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1918
timestamp 1677622389
transform 1 0 3788 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1677622389
transform 1 0 3788 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2315
timestamp 1677622389
transform 1 0 3796 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1677622389
transform 1 0 3812 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1677622389
transform 1 0 3788 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1677622389
transform 1 0 3804 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1677622389
transform 1 0 3812 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1677622389
transform 1 0 3836 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1677622389
transform 1 0 3844 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1983
timestamp 1677622389
transform 1 0 3868 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1677622389
transform 1 0 3892 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2318
timestamp 1677622389
transform 1 0 3868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1677622389
transform 1 0 3884 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1677622389
transform 1 0 3892 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1677622389
transform 1 0 3876 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1677622389
transform 1 0 3908 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1677622389
transform 1 0 3948 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1985
timestamp 1677622389
transform 1 0 4036 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2321
timestamp 1677622389
transform 1 0 4036 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1677622389
transform 1 0 3988 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1897
timestamp 1677622389
transform 1 0 4108 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1677622389
transform 1 0 4116 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1677622389
transform 1 0 4140 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1677622389
transform 1 0 4132 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2322
timestamp 1677622389
transform 1 0 4116 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1677622389
transform 1 0 4124 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1677622389
transform 1 0 4140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1677622389
transform 1 0 4116 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1677622389
transform 1 0 4132 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1677622389
transform 1 0 4148 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2077
timestamp 1677622389
transform 1 0 4116 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2224
timestamp 1677622389
transform 1 0 4172 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1887
timestamp 1677622389
transform 1 0 4196 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2211
timestamp 1677622389
transform 1 0 4196 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1677622389
transform 1 0 4204 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1987
timestamp 1677622389
transform 1 0 4212 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2325
timestamp 1677622389
transform 1 0 4204 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1677622389
transform 1 0 4228 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2078
timestamp 1677622389
transform 1 0 4228 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2326
timestamp 1677622389
transform 1 0 4260 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1677622389
transform 1 0 4284 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1677622389
transform 1 0 4276 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1948
timestamp 1677622389
transform 1 0 4300 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2328
timestamp 1677622389
transform 1 0 4300 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1677622389
transform 1 0 4316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1677622389
transform 1 0 4324 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1677622389
transform 1 0 4356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1677622389
transform 1 0 4348 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1898
timestamp 1677622389
transform 1 0 4380 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2330
timestamp 1677622389
transform 1 0 4388 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2013
timestamp 1677622389
transform 1 0 4396 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2430
timestamp 1677622389
transform 1 0 4380 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2032
timestamp 1677622389
transform 1 0 4404 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2331
timestamp 1677622389
transform 1 0 4420 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1677622389
transform 1 0 4412 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2033
timestamp 1677622389
transform 1 0 4420 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1677622389
transform 1 0 4428 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1677622389
transform 1 0 4444 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1677622389
transform 1 0 4460 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2332
timestamp 1677622389
transform 1 0 4444 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1677622389
transform 1 0 4436 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2079
timestamp 1677622389
transform 1 0 4436 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1677622389
transform 1 0 4452 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1677622389
transform 1 0 4484 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1677622389
transform 1 0 4484 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2333
timestamp 1677622389
transform 1 0 4460 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1677622389
transform 1 0 4476 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1677622389
transform 1 0 4452 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2058
timestamp 1677622389
transform 1 0 4468 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2434
timestamp 1677622389
transform 1 0 4484 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1677622389
transform 1 0 4492 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2080
timestamp 1677622389
transform 1 0 4516 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1677622389
transform 1 0 4532 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1677622389
transform 1 0 4524 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2336
timestamp 1677622389
transform 1 0 4532 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2034
timestamp 1677622389
transform 1 0 4532 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2435
timestamp 1677622389
transform 1 0 4540 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1899
timestamp 1677622389
transform 1 0 4572 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2226
timestamp 1677622389
transform 1 0 4612 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2015
timestamp 1677622389
transform 1 0 4612 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2227
timestamp 1677622389
transform 1 0 4628 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1923
timestamp 1677622389
transform 1 0 4660 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1677622389
transform 1 0 4660 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2337
timestamp 1677622389
transform 1 0 4636 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1677622389
transform 1 0 4644 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2016
timestamp 1677622389
transform 1 0 4652 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2339
timestamp 1677622389
transform 1 0 4660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1677622389
transform 1 0 4636 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1677622389
transform 1 0 4652 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1677622389
transform 1 0 4668 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2059
timestamp 1677622389
transform 1 0 4652 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1677622389
transform 1 0 4740 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1677622389
transform 1 0 4796 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1677622389
transform 1 0 4724 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1677622389
transform 1 0 4780 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1677622389
transform 1 0 4700 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2060
timestamp 1677622389
transform 1 0 4724 0 1 3595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_22
timestamp 1677622389
transform 1 0 48 0 1 3570
box -10 -3 10 3
use FILL  FILL_2209
timestamp 1677622389
transform 1 0 72 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1677622389
transform 1 0 80 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_2081
timestamp 1677622389
transform 1 0 188 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_187
timestamp 1677622389
transform -1 0 192 0 1 3570
box -9 -3 26 105
use FILL  FILL_2210
timestamp 1677622389
transform 1 0 192 0 1 3570
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1677622389
transform 1 0 200 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_103
timestamp 1677622389
transform 1 0 208 0 1 3570
box -8 -3 46 105
use FILL  FILL_2214
timestamp 1677622389
transform 1 0 248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1677622389
transform 1 0 256 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2082
timestamp 1677622389
transform 1 0 332 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1677622389
transform 1 0 348 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_162
timestamp 1677622389
transform 1 0 264 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_189
timestamp 1677622389
transform -1 0 376 0 1 3570
box -9 -3 26 105
use FILL  FILL_2218
timestamp 1677622389
transform 1 0 376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1677622389
transform 1 0 384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1677622389
transform 1 0 392 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_105
timestamp 1677622389
transform -1 0 440 0 1 3570
box -8 -3 46 105
use FILL  FILL_2221
timestamp 1677622389
transform 1 0 440 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1677622389
transform 1 0 448 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_2084
timestamp 1677622389
transform 1 0 556 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_190
timestamp 1677622389
transform -1 0 560 0 1 3570
box -9 -3 26 105
use FILL  FILL_2222
timestamp 1677622389
transform 1 0 560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1677622389
transform 1 0 568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1677622389
transform 1 0 576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1677622389
transform 1 0 584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1677622389
transform 1 0 592 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2085
timestamp 1677622389
transform 1 0 644 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_106
timestamp 1677622389
transform 1 0 600 0 1 3570
box -8 -3 46 105
use FILL  FILL_2227
timestamp 1677622389
transform 1 0 640 0 1 3570
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1677622389
transform 1 0 648 0 1 3570
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1677622389
transform 1 0 656 0 1 3570
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1677622389
transform 1 0 664 0 1 3570
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1677622389
transform 1 0 672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1677622389
transform 1 0 680 0 1 3570
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1677622389
transform 1 0 688 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_192
timestamp 1677622389
transform 1 0 696 0 1 3570
box -9 -3 26 105
use FILL  FILL_2245
timestamp 1677622389
transform 1 0 712 0 1 3570
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1677622389
transform 1 0 720 0 1 3570
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1677622389
transform 1 0 728 0 1 3570
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1677622389
transform 1 0 736 0 1 3570
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1677622389
transform 1 0 744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1677622389
transform 1 0 752 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_52
timestamp 1677622389
transform -1 0 792 0 1 3570
box -8 -3 34 105
use FILL  FILL_2255
timestamp 1677622389
transform 1 0 792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1677622389
transform 1 0 800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1677622389
transform 1 0 808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1677622389
transform 1 0 816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1677622389
transform 1 0 824 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_193
timestamp 1677622389
transform -1 0 848 0 1 3570
box -9 -3 26 105
use FILL  FILL_2260
timestamp 1677622389
transform 1 0 848 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2086
timestamp 1677622389
transform 1 0 892 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_109
timestamp 1677622389
transform 1 0 856 0 1 3570
box -8 -3 46 105
use FILL  FILL_2269
timestamp 1677622389
transform 1 0 896 0 1 3570
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1677622389
transform 1 0 904 0 1 3570
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1677622389
transform 1 0 912 0 1 3570
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1677622389
transform 1 0 920 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_110
timestamp 1677622389
transform 1 0 928 0 1 3570
box -8 -3 46 105
use FILL  FILL_2277
timestamp 1677622389
transform 1 0 968 0 1 3570
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1677622389
transform 1 0 976 0 1 3570
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1677622389
transform 1 0 984 0 1 3570
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1677622389
transform 1 0 992 0 1 3570
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1677622389
transform 1 0 1000 0 1 3570
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1677622389
transform 1 0 1008 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2087
timestamp 1677622389
transform 1 0 1044 0 1 3575
box -3 -3 3 3
use OAI21X1  OAI21X1_53
timestamp 1677622389
transform 1 0 1016 0 1 3570
box -8 -3 34 105
use FILL  FILL_2284
timestamp 1677622389
transform 1 0 1048 0 1 3570
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1677622389
transform 1 0 1056 0 1 3570
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1677622389
transform 1 0 1064 0 1 3570
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1677622389
transform 1 0 1072 0 1 3570
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1677622389
transform 1 0 1080 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_194
timestamp 1677622389
transform 1 0 1088 0 1 3570
box -9 -3 26 105
use FILL  FILL_2295
timestamp 1677622389
transform 1 0 1104 0 1 3570
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1677622389
transform 1 0 1112 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_111
timestamp 1677622389
transform 1 0 1120 0 1 3570
box -8 -3 46 105
use FILL  FILL_2297
timestamp 1677622389
transform 1 0 1160 0 1 3570
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1677622389
transform 1 0 1168 0 1 3570
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1677622389
transform 1 0 1176 0 1 3570
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1677622389
transform 1 0 1184 0 1 3570
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1677622389
transform 1 0 1192 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1677622389
transform -1 0 1232 0 1 3570
box -8 -3 34 105
use FILL  FILL_2303
timestamp 1677622389
transform 1 0 1232 0 1 3570
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1677622389
transform 1 0 1240 0 1 3570
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1677622389
transform 1 0 1248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1677622389
transform 1 0 1256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1677622389
transform 1 0 1264 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_56
timestamp 1677622389
transform -1 0 1304 0 1 3570
box -8 -3 34 105
use FILL  FILL_2313
timestamp 1677622389
transform 1 0 1304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1677622389
transform 1 0 1312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1677622389
transform 1 0 1320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1677622389
transform 1 0 1328 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1677622389
transform 1 0 1336 0 1 3570
box -8 -3 32 105
use FILL  FILL_2320
timestamp 1677622389
transform 1 0 1360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1677622389
transform 1 0 1368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1677622389
transform 1 0 1376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1677622389
transform 1 0 1384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1677622389
transform 1 0 1392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1677622389
transform 1 0 1400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1677622389
transform 1 0 1408 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_167
timestamp 1677622389
transform -1 0 1512 0 1 3570
box -8 -3 104 105
use FILL  FILL_2333
timestamp 1677622389
transform 1 0 1512 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_168
timestamp 1677622389
transform 1 0 1520 0 1 3570
box -8 -3 104 105
use FILL  FILL_2334
timestamp 1677622389
transform 1 0 1616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1677622389
transform 1 0 1624 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2088
timestamp 1677622389
transform 1 0 1676 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1677622389
transform 1 0 1708 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1677622389
transform 1 0 1732 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_169
timestamp 1677622389
transform -1 0 1728 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_198
timestamp 1677622389
transform -1 0 1744 0 1 3570
box -9 -3 26 105
use FILL  FILL_2354
timestamp 1677622389
transform 1 0 1744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1677622389
transform 1 0 1752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1677622389
transform 1 0 1760 0 1 3570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1677622389
transform 1 0 1768 0 1 3570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1677622389
transform 1 0 1776 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_112
timestamp 1677622389
transform -1 0 1824 0 1 3570
box -8 -3 46 105
use FILL  FILL_2367
timestamp 1677622389
transform 1 0 1824 0 1 3570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1677622389
transform 1 0 1832 0 1 3570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1677622389
transform 1 0 1840 0 1 3570
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1677622389
transform 1 0 1848 0 1 3570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1677622389
transform 1 0 1856 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1677622389
transform 1 0 1864 0 1 3570
box -8 -3 104 105
use AOI22X1  AOI22X1_113
timestamp 1677622389
transform 1 0 1960 0 1 3570
box -8 -3 46 105
use FILL  FILL_2372
timestamp 1677622389
transform 1 0 2000 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1677622389
transform 1 0 2008 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1677622389
transform 1 0 2104 0 1 3570
box -8 -3 104 105
use FILL  FILL_2385
timestamp 1677622389
transform 1 0 2200 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_114
timestamp 1677622389
transform 1 0 2208 0 1 3570
box -8 -3 46 105
use FILL  FILL_2404
timestamp 1677622389
transform 1 0 2248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1677622389
transform 1 0 2256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1677622389
transform 1 0 2264 0 1 3570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1677622389
transform 1 0 2272 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_201
timestamp 1677622389
transform -1 0 2296 0 1 3570
box -9 -3 26 105
use FILL  FILL_2413
timestamp 1677622389
transform 1 0 2296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1677622389
transform 1 0 2304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1677622389
transform 1 0 2312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1677622389
transform 1 0 2320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1677622389
transform 1 0 2328 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_115
timestamp 1677622389
transform -1 0 2376 0 1 3570
box -8 -3 46 105
use FILL  FILL_2418
timestamp 1677622389
transform 1 0 2376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1677622389
transform 1 0 2384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1677622389
transform 1 0 2392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1677622389
transform 1 0 2400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1677622389
transform 1 0 2408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1677622389
transform 1 0 2416 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_202
timestamp 1677622389
transform 1 0 2424 0 1 3570
box -9 -3 26 105
use FILL  FILL_2424
timestamp 1677622389
transform 1 0 2440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1677622389
transform 1 0 2448 0 1 3570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1677622389
transform 1 0 2456 0 1 3570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1677622389
transform 1 0 2464 0 1 3570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1677622389
transform 1 0 2472 0 1 3570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1677622389
transform 1 0 2480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1677622389
transform 1 0 2488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1677622389
transform 1 0 2496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1677622389
transform 1 0 2504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1677622389
transform 1 0 2512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1677622389
transform 1 0 2520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1677622389
transform 1 0 2528 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_203
timestamp 1677622389
transform 1 0 2536 0 1 3570
box -9 -3 26 105
use FILL  FILL_2445
timestamp 1677622389
transform 1 0 2552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1677622389
transform 1 0 2560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1677622389
transform 1 0 2568 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1677622389
transform 1 0 2576 0 1 3570
box -8 -3 104 105
use FILL  FILL_2452
timestamp 1677622389
transform 1 0 2672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1677622389
transform 1 0 2680 0 1 3570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1677622389
transform 1 0 2688 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1677622389
transform 1 0 2696 0 1 3570
box -8 -3 34 105
use FILL  FILL_2455
timestamp 1677622389
transform 1 0 2728 0 1 3570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1677622389
transform 1 0 2736 0 1 3570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1677622389
transform 1 0 2744 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_30
timestamp 1677622389
transform 1 0 2752 0 1 3570
box -8 -3 32 105
use FILL  FILL_2469
timestamp 1677622389
transform 1 0 2776 0 1 3570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1677622389
transform 1 0 2784 0 1 3570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1677622389
transform 1 0 2792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1677622389
transform 1 0 2800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1677622389
transform 1 0 2808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1677622389
transform 1 0 2816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1677622389
transform 1 0 2824 0 1 3570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1677622389
transform 1 0 2832 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_58
timestamp 1677622389
transform -1 0 2872 0 1 3570
box -8 -3 34 105
use FILL  FILL_2477
timestamp 1677622389
transform 1 0 2872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1677622389
transform 1 0 2880 0 1 3570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1677622389
transform 1 0 2888 0 1 3570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1677622389
transform 1 0 2896 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_204
timestamp 1677622389
transform 1 0 2904 0 1 3570
box -9 -3 26 105
use OAI21X1  OAI21X1_61
timestamp 1677622389
transform -1 0 2952 0 1 3570
box -8 -3 34 105
use M3_M2  M3_M2_2091
timestamp 1677622389
transform 1 0 3020 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_176
timestamp 1677622389
transform 1 0 2952 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_205
timestamp 1677622389
transform 1 0 3048 0 1 3570
box -9 -3 26 105
use FILL  FILL_2489
timestamp 1677622389
transform 1 0 3064 0 1 3570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1677622389
transform 1 0 3072 0 1 3570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1677622389
transform 1 0 3080 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_110
timestamp 1677622389
transform -1 0 3128 0 1 3570
box -8 -3 46 105
use FILL  FILL_2502
timestamp 1677622389
transform 1 0 3128 0 1 3570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1677622389
transform 1 0 3136 0 1 3570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1677622389
transform 1 0 3144 0 1 3570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1677622389
transform 1 0 3152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1677622389
transform 1 0 3160 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_111
timestamp 1677622389
transform -1 0 3208 0 1 3570
box -8 -3 46 105
use FILL  FILL_2513
timestamp 1677622389
transform 1 0 3208 0 1 3570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1677622389
transform 1 0 3216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1677622389
transform 1 0 3224 0 1 3570
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1677622389
transform 1 0 3232 0 1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1677622389
transform -1 0 3272 0 1 3570
box -8 -3 40 105
use FILL  FILL_2517
timestamp 1677622389
transform 1 0 3272 0 1 3570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1677622389
transform 1 0 3280 0 1 3570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1677622389
transform 1 0 3288 0 1 3570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1677622389
transform 1 0 3296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1677622389
transform 1 0 3304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1677622389
transform 1 0 3312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1677622389
transform 1 0 3320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1677622389
transform 1 0 3328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1677622389
transform 1 0 3336 0 1 3570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1677622389
transform 1 0 3344 0 1 3570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1677622389
transform 1 0 3352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1677622389
transform 1 0 3360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1677622389
transform 1 0 3368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1677622389
transform 1 0 3376 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_207
timestamp 1677622389
transform -1 0 3400 0 1 3570
box -9 -3 26 105
use FILL  FILL_2542
timestamp 1677622389
transform 1 0 3400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1677622389
transform 1 0 3408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1677622389
transform 1 0 3416 0 1 3570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1677622389
transform 1 0 3424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1677622389
transform 1 0 3432 0 1 3570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1677622389
transform 1 0 3440 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2092
timestamp 1677622389
transform 1 0 3492 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_113
timestamp 1677622389
transform -1 0 3488 0 1 3570
box -8 -3 46 105
use FILL  FILL_2552
timestamp 1677622389
transform 1 0 3488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1677622389
transform 1 0 3496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1677622389
transform 1 0 3504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1677622389
transform 1 0 3512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1677622389
transform 1 0 3520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1677622389
transform 1 0 3528 0 1 3570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1677622389
transform 1 0 3536 0 1 3570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1677622389
transform 1 0 3544 0 1 3570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1677622389
transform 1 0 3552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1677622389
transform 1 0 3560 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_114
timestamp 1677622389
transform 1 0 3568 0 1 3570
box -8 -3 46 105
use FILL  FILL_2571
timestamp 1677622389
transform 1 0 3608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1677622389
transform 1 0 3616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1677622389
transform 1 0 3624 0 1 3570
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1677622389
transform 1 0 3632 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2093
timestamp 1677622389
transform 1 0 3708 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_177
timestamp 1677622389
transform 1 0 3640 0 1 3570
box -8 -3 104 105
use FILL  FILL_2575
timestamp 1677622389
transform 1 0 3736 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2094
timestamp 1677622389
transform 1 0 3756 0 1 3575
box -3 -3 3 3
use FILL  FILL_2576
timestamp 1677622389
transform 1 0 3744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1677622389
transform 1 0 3752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1677622389
transform 1 0 3760 0 1 3570
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1677622389
transform 1 0 3768 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2095
timestamp 1677622389
transform 1 0 3796 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1677622389
transform 1 0 3820 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_118
timestamp 1677622389
transform 1 0 3776 0 1 3570
box -8 -3 46 105
use FILL  FILL_2587
timestamp 1677622389
transform 1 0 3816 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2097
timestamp 1677622389
transform 1 0 3836 0 1 3575
box -3 -3 3 3
use FILL  FILL_2588
timestamp 1677622389
transform 1 0 3824 0 1 3570
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1677622389
transform 1 0 3832 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2098
timestamp 1677622389
transform 1 0 3860 0 1 3575
box -3 -3 3 3
use FILL  FILL_2590
timestamp 1677622389
transform 1 0 3840 0 1 3570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1677622389
transform 1 0 3848 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_117
timestamp 1677622389
transform -1 0 3896 0 1 3570
box -8 -3 46 105
use FILL  FILL_2592
timestamp 1677622389
transform 1 0 3896 0 1 3570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1677622389
transform 1 0 3904 0 1 3570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1677622389
transform 1 0 3912 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_208
timestamp 1677622389
transform -1 0 3936 0 1 3570
box -9 -3 26 105
use FILL  FILL_2595
timestamp 1677622389
transform 1 0 3936 0 1 3570
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1677622389
transform 1 0 3944 0 1 3570
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1677622389
transform 1 0 3952 0 1 3570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1677622389
transform 1 0 3960 0 1 3570
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1677622389
transform 1 0 3968 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1677622389
transform 1 0 3976 0 1 3570
box -8 -3 104 105
use FILL  FILL_2607
timestamp 1677622389
transform 1 0 4072 0 1 3570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1677622389
transform 1 0 4080 0 1 3570
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1677622389
transform 1 0 4088 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_210
timestamp 1677622389
transform 1 0 4096 0 1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_119
timestamp 1677622389
transform 1 0 4112 0 1 3570
box -8 -3 46 105
use FILL  FILL_2615
timestamp 1677622389
transform 1 0 4152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1677622389
transform 1 0 4160 0 1 3570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1677622389
transform 1 0 4168 0 1 3570
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1677622389
transform 1 0 4176 0 1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1677622389
transform -1 0 4216 0 1 3570
box -8 -3 40 105
use FILL  FILL_2619
timestamp 1677622389
transform 1 0 4216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1677622389
transform 1 0 4224 0 1 3570
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1677622389
transform 1 0 4232 0 1 3570
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1677622389
transform 1 0 4240 0 1 3570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1677622389
transform 1 0 4248 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_120
timestamp 1677622389
transform 1 0 4256 0 1 3570
box -8 -3 46 105
use FILL  FILL_2624
timestamp 1677622389
transform 1 0 4296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1677622389
transform 1 0 4304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1677622389
transform 1 0 4312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1677622389
transform 1 0 4320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1677622389
transform 1 0 4328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1677622389
transform 1 0 4336 0 1 3570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1677622389
transform 1 0 4344 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2099
timestamp 1677622389
transform 1 0 4364 0 1 3575
box -3 -3 3 3
use FILL  FILL_2631
timestamp 1677622389
transform 1 0 4352 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_121
timestamp 1677622389
transform 1 0 4360 0 1 3570
box -8 -3 46 105
use FILL  FILL_2632
timestamp 1677622389
transform 1 0 4400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1677622389
transform 1 0 4408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1677622389
transform 1 0 4416 0 1 3570
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1677622389
transform 1 0 4424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1677622389
transform 1 0 4432 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2100
timestamp 1677622389
transform 1 0 4452 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_120
timestamp 1677622389
transform -1 0 4480 0 1 3570
box -8 -3 46 105
use FILL  FILL_2652
timestamp 1677622389
transform 1 0 4480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1677622389
transform 1 0 4488 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_211
timestamp 1677622389
transform -1 0 4512 0 1 3570
box -9 -3 26 105
use FILL  FILL_2654
timestamp 1677622389
transform 1 0 4512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1677622389
transform 1 0 4520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1677622389
transform 1 0 4528 0 1 3570
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1677622389
transform 1 0 4536 0 1 3570
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1677622389
transform 1 0 4544 0 1 3570
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1677622389
transform 1 0 4552 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_212
timestamp 1677622389
transform -1 0 4576 0 1 3570
box -9 -3 26 105
use FILL  FILL_2660
timestamp 1677622389
transform 1 0 4576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1677622389
transform 1 0 4584 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2101
timestamp 1677622389
transform 1 0 4604 0 1 3575
box -3 -3 3 3
use FILL  FILL_2662
timestamp 1677622389
transform 1 0 4592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1677622389
transform 1 0 4600 0 1 3570
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1677622389
transform 1 0 4608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1677622389
transform 1 0 4616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1677622389
transform 1 0 4624 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_122
timestamp 1677622389
transform 1 0 4632 0 1 3570
box -8 -3 46 105
use FILL  FILL_2667
timestamp 1677622389
transform 1 0 4672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1677622389
transform 1 0 4680 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1677622389
transform 1 0 4688 0 1 3570
box -8 -3 104 105
use FILL  FILL_2669
timestamp 1677622389
transform 1 0 4784 0 1 3570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_23
timestamp 1677622389
transform 1 0 4819 0 1 3570
box -10 -3 10 3
use M3_M2  M3_M2_2126
timestamp 1677622389
transform 1 0 84 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1677622389
transform 1 0 164 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2449
timestamp 1677622389
transform 1 0 84 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1677622389
transform 1 0 132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1677622389
transform 1 0 164 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1677622389
transform 1 0 172 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2232
timestamp 1677622389
transform 1 0 132 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1677622389
transform 1 0 172 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1677622389
transform 1 0 188 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1677622389
transform 1 0 228 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2450
timestamp 1677622389
transform 1 0 204 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1677622389
transform 1 0 212 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1677622389
transform 1 0 228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1677622389
transform 1 0 196 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2209
timestamp 1677622389
transform 1 0 212 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2559
timestamp 1677622389
transform 1 0 220 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1677622389
transform 1 0 236 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2266
timestamp 1677622389
transform 1 0 236 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1677622389
transform 1 0 276 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2441
timestamp 1677622389
transform 1 0 308 0 1 3555
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1677622389
transform 1 0 284 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1677622389
transform 1 0 300 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1677622389
transform 1 0 276 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1677622389
transform 1 0 300 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2280
timestamp 1677622389
transform 1 0 292 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1677622389
transform 1 0 340 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1677622389
transform 1 0 324 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1677622389
transform 1 0 316 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1677622389
transform 1 0 412 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2455
timestamp 1677622389
transform 1 0 332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1677622389
transform 1 0 380 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1677622389
transform 1 0 412 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1677622389
transform 1 0 420 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1677622389
transform 1 0 380 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1677622389
transform 1 0 420 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1677622389
transform 1 0 452 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2566
timestamp 1677622389
transform 1 0 444 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2131
timestamp 1677622389
transform 1 0 484 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1677622389
transform 1 0 492 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2456
timestamp 1677622389
transform 1 0 468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1677622389
transform 1 0 476 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1677622389
transform 1 0 492 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1677622389
transform 1 0 508 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2210
timestamp 1677622389
transform 1 0 476 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2567
timestamp 1677622389
transform 1 0 484 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1677622389
transform 1 0 500 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2267
timestamp 1677622389
transform 1 0 500 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2460
timestamp 1677622389
transform 1 0 532 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2236
timestamp 1677622389
transform 1 0 524 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1677622389
transform 1 0 612 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1677622389
transform 1 0 604 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1677622389
transform 1 0 580 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1677622389
transform 1 0 596 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1677622389
transform 1 0 620 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2461
timestamp 1677622389
transform 1 0 564 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2191
timestamp 1677622389
transform 1 0 572 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2462
timestamp 1677622389
transform 1 0 580 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1677622389
transform 1 0 596 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1677622389
transform 1 0 612 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1677622389
transform 1 0 620 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1677622389
transform 1 0 548 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1677622389
transform 1 0 556 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1677622389
transform 1 0 572 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1677622389
transform 1 0 588 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2237
timestamp 1677622389
transform 1 0 572 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1677622389
transform 1 0 548 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1677622389
transform 1 0 596 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2573
timestamp 1677622389
transform 1 0 604 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1677622389
transform 1 0 620 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2268
timestamp 1677622389
transform 1 0 612 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1677622389
transform 1 0 668 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2466
timestamp 1677622389
transform 1 0 660 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1677622389
transform 1 0 652 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1677622389
transform 1 0 668 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2238
timestamp 1677622389
transform 1 0 644 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1677622389
transform 1 0 668 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2443
timestamp 1677622389
transform 1 0 692 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1677622389
transform 1 0 684 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2281
timestamp 1677622389
transform 1 0 692 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1677622389
transform 1 0 684 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2468
timestamp 1677622389
transform 1 0 724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1677622389
transform 1 0 732 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2282
timestamp 1677622389
transform 1 0 724 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1677622389
transform 1 0 716 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2577
timestamp 1677622389
transform 1 0 748 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1677622389
transform 1 0 756 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2283
timestamp 1677622389
transform 1 0 740 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1677622389
transform 1 0 772 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2470
timestamp 1677622389
transform 1 0 780 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2105
timestamp 1677622389
transform 1 0 820 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1677622389
transform 1 0 804 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2444
timestamp 1677622389
transform 1 0 828 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1677622389
transform 1 0 804 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1677622389
transform 1 0 820 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1677622389
transform 1 0 812 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2192
timestamp 1677622389
transform 1 0 828 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2473
timestamp 1677622389
transform 1 0 852 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2307
timestamp 1677622389
transform 1 0 868 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2580
timestamp 1677622389
transform 1 0 892 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2166
timestamp 1677622389
transform 1 0 924 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1677622389
transform 1 0 948 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2474
timestamp 1677622389
transform 1 0 924 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1677622389
transform 1 0 956 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2284
timestamp 1677622389
transform 1 0 924 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2582
timestamp 1677622389
transform 1 0 1012 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2135
timestamp 1677622389
transform 1 0 1028 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2445
timestamp 1677622389
transform 1 0 1028 0 1 3545
box -2 -2 2 2
use M3_M2  M3_M2_2136
timestamp 1677622389
transform 1 0 1076 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1677622389
transform 1 0 1076 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2475
timestamp 1677622389
transform 1 0 1068 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1677622389
transform 1 0 1076 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2308
timestamp 1677622389
transform 1 0 1068 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1677622389
transform 1 0 1100 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1677622389
transform 1 0 1132 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2476
timestamp 1677622389
transform 1 0 1100 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1677622389
transform 1 0 1124 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1677622389
transform 1 0 1180 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2285
timestamp 1677622389
transform 1 0 1100 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1677622389
transform 1 0 1108 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1677622389
transform 1 0 1252 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1677622389
transform 1 0 1244 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1677622389
transform 1 0 1228 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2477
timestamp 1677622389
transform 1 0 1244 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1677622389
transform 1 0 1228 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2286
timestamp 1677622389
transform 1 0 1228 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2478
timestamp 1677622389
transform 1 0 1252 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1677622389
transform 1 0 1260 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2287
timestamp 1677622389
transform 1 0 1260 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1677622389
transform 1 0 1292 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2479
timestamp 1677622389
transform 1 0 1300 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1677622389
transform 1 0 1292 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1677622389
transform 1 0 1332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1677622389
transform 1 0 1340 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1677622389
transform 1 0 1324 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2288
timestamp 1677622389
transform 1 0 1324 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1677622389
transform 1 0 1340 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2589
timestamp 1677622389
transform 1 0 1388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2170
timestamp 1677622389
transform 1 0 1412 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2590
timestamp 1677622389
transform 1 0 1412 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2289
timestamp 1677622389
transform 1 0 1420 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1677622389
transform 1 0 1436 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1677622389
transform 1 0 1444 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2482
timestamp 1677622389
transform 1 0 1468 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2310
timestamp 1677622389
transform 1 0 1460 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1677622389
transform 1 0 1516 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2483
timestamp 1677622389
transform 1 0 1524 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1677622389
transform 1 0 1516 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1677622389
transform 1 0 1532 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2311
timestamp 1677622389
transform 1 0 1532 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2484
timestamp 1677622389
transform 1 0 1548 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2290
timestamp 1677622389
transform 1 0 1548 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2593
timestamp 1677622389
transform 1 0 1564 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1677622389
transform 1 0 1572 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1677622389
transform 1 0 1580 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2195
timestamp 1677622389
transform 1 0 1588 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2595
timestamp 1677622389
transform 1 0 1588 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2269
timestamp 1677622389
transform 1 0 1572 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2486
timestamp 1677622389
transform 1 0 1612 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1677622389
transform 1 0 1628 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1677622389
transform 1 0 1660 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1677622389
transform 1 0 1684 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1677622389
transform 1 0 1652 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1677622389
transform 1 0 1676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1677622389
transform 1 0 1740 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1677622389
transform 1 0 1724 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1677622389
transform 1 0 1732 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2240
timestamp 1677622389
transform 1 0 1724 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1677622389
transform 1 0 1732 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1677622389
transform 1 0 1788 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2491
timestamp 1677622389
transform 1 0 1780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1677622389
transform 1 0 1796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1677622389
transform 1 0 1772 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2196
timestamp 1677622389
transform 1 0 1804 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2601
timestamp 1677622389
transform 1 0 1804 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2109
timestamp 1677622389
transform 1 0 1860 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1677622389
transform 1 0 1908 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2493
timestamp 1677622389
transform 1 0 1908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1677622389
transform 1 0 1828 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1677622389
transform 1 0 1868 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2292
timestamp 1677622389
transform 1 0 1884 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1677622389
transform 1 0 1844 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1677622389
transform 1 0 1916 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1677622389
transform 1 0 1972 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1677622389
transform 1 0 1996 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1677622389
transform 1 0 2020 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2494
timestamp 1677622389
transform 1 0 2028 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2212
timestamp 1677622389
transform 1 0 2028 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2604
timestamp 1677622389
transform 1 0 2044 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2294
timestamp 1677622389
transform 1 0 2036 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1677622389
transform 1 0 2100 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2495
timestamp 1677622389
transform 1 0 2092 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2213
timestamp 1677622389
transform 1 0 2092 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1677622389
transform 1 0 2188 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2496
timestamp 1677622389
transform 1 0 2172 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1677622389
transform 1 0 2188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1677622389
transform 1 0 2164 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2214
timestamp 1677622389
transform 1 0 2172 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2606
timestamp 1677622389
transform 1 0 2180 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1677622389
transform 1 0 2204 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1677622389
transform 1 0 2204 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1677622389
transform 1 0 2228 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2498
timestamp 1677622389
transform 1 0 2228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1677622389
transform 1 0 2236 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2111
timestamp 1677622389
transform 1 0 2260 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1677622389
transform 1 0 2260 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2608
timestamp 1677622389
transform 1 0 2276 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2144
timestamp 1677622389
transform 1 0 2316 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2500
timestamp 1677622389
transform 1 0 2316 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1677622389
transform 1 0 2324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1677622389
transform 1 0 2348 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2215
timestamp 1677622389
transform 1 0 2348 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1677622389
transform 1 0 2380 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1677622389
transform 1 0 2372 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1677622389
transform 1 0 2388 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2502
timestamp 1677622389
transform 1 0 2460 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2216
timestamp 1677622389
transform 1 0 2412 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2610
timestamp 1677622389
transform 1 0 2436 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2243
timestamp 1677622389
transform 1 0 2436 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1677622389
transform 1 0 2404 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1677622389
transform 1 0 2452 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1677622389
transform 1 0 2476 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2611
timestamp 1677622389
transform 1 0 2476 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2173
timestamp 1677622389
transform 1 0 2516 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2503
timestamp 1677622389
transform 1 0 2516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1677622389
transform 1 0 2508 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2217
timestamp 1677622389
transform 1 0 2516 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2613
timestamp 1677622389
transform 1 0 2524 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2244
timestamp 1677622389
transform 1 0 2524 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1677622389
transform 1 0 2548 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2504
timestamp 1677622389
transform 1 0 2556 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1677622389
transform 1 0 2548 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1677622389
transform 1 0 2572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1677622389
transform 1 0 2564 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2245
timestamp 1677622389
transform 1 0 2572 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1677622389
transform 1 0 2564 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2446
timestamp 1677622389
transform 1 0 2644 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1677622389
transform 1 0 2620 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1677622389
transform 1 0 2636 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2218
timestamp 1677622389
transform 1 0 2660 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2506
timestamp 1677622389
transform 1 0 2676 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2246
timestamp 1677622389
transform 1 0 2676 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2447
timestamp 1677622389
transform 1 0 2692 0 1 3545
box -2 -2 2 2
use M3_M2  M3_M2_2197
timestamp 1677622389
transform 1 0 2692 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2618
timestamp 1677622389
transform 1 0 2700 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1677622389
transform 1 0 2716 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1677622389
transform 1 0 2724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1677622389
transform 1 0 2740 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1677622389
transform 1 0 2732 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2318
timestamp 1677622389
transform 1 0 2724 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2510
timestamp 1677622389
transform 1 0 2796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1677622389
transform 1 0 2804 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1677622389
transform 1 0 2780 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1677622389
transform 1 0 2796 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2219
timestamp 1677622389
transform 1 0 2804 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2669
timestamp 1677622389
transform 1 0 2796 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2145
timestamp 1677622389
transform 1 0 2836 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2448
timestamp 1677622389
transform 1 0 2836 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1677622389
transform 1 0 2844 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2220
timestamp 1677622389
transform 1 0 2836 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1677622389
transform 1 0 2828 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2670
timestamp 1677622389
transform 1 0 2836 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2248
timestamp 1677622389
transform 1 0 2844 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1677622389
transform 1 0 2884 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2513
timestamp 1677622389
transform 1 0 2884 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1677622389
transform 1 0 2892 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1677622389
transform 1 0 2884 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2221
timestamp 1677622389
transform 1 0 2892 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1677622389
transform 1 0 2884 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2671
timestamp 1677622389
transform 1 0 2900 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1677622389
transform 1 0 2932 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2222
timestamp 1677622389
transform 1 0 2964 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2515
timestamp 1677622389
transform 1 0 2980 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2115
timestamp 1677622389
transform 1 0 3004 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1677622389
transform 1 0 3004 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1677622389
transform 1 0 3028 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2516
timestamp 1677622389
transform 1 0 3020 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1677622389
transform 1 0 3036 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1677622389
transform 1 0 3020 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1677622389
transform 1 0 3028 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1677622389
transform 1 0 3044 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2250
timestamp 1677622389
transform 1 0 3020 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1677622389
transform 1 0 3044 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1677622389
transform 1 0 3012 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2518
timestamp 1677622389
transform 1 0 3068 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2223
timestamp 1677622389
transform 1 0 3060 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1677622389
transform 1 0 3108 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2519
timestamp 1677622389
transform 1 0 3108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1677622389
transform 1 0 3100 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2252
timestamp 1677622389
transform 1 0 3084 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1677622389
transform 1 0 3100 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1677622389
transform 1 0 3148 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1677622389
transform 1 0 3164 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2628
timestamp 1677622389
transform 1 0 3164 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1677622389
transform 1 0 3204 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1677622389
transform 1 0 3196 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2270
timestamp 1677622389
transform 1 0 3188 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1677622389
transform 1 0 3204 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1677622389
transform 1 0 3220 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2630
timestamp 1677622389
transform 1 0 3228 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2224
timestamp 1677622389
transform 1 0 3236 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2676
timestamp 1677622389
transform 1 0 3220 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1677622389
transform 1 0 3260 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1677622389
transform 1 0 3292 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1677622389
transform 1 0 3284 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2254
timestamp 1677622389
transform 1 0 3292 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1677622389
transform 1 0 3284 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1677622389
transform 1 0 3332 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1677622389
transform 1 0 3364 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2521
timestamp 1677622389
transform 1 0 3332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1677622389
transform 1 0 3348 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2200
timestamp 1677622389
transform 1 0 3356 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2523
timestamp 1677622389
transform 1 0 3364 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1677622389
transform 1 0 3340 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1677622389
transform 1 0 3356 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1677622389
transform 1 0 3364 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2255
timestamp 1677622389
transform 1 0 3340 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1677622389
transform 1 0 3428 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2524
timestamp 1677622389
transform 1 0 3412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1677622389
transform 1 0 3420 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2225
timestamp 1677622389
transform 1 0 3420 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2635
timestamp 1677622389
transform 1 0 3428 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2256
timestamp 1677622389
transform 1 0 3436 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1677622389
transform 1 0 3452 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2526
timestamp 1677622389
transform 1 0 3452 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1677622389
transform 1 0 3460 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1677622389
transform 1 0 3476 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2527
timestamp 1677622389
transform 1 0 3484 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2272
timestamp 1677622389
transform 1 0 3484 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2528
timestamp 1677622389
transform 1 0 3508 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2226
timestamp 1677622389
transform 1 0 3508 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2442
timestamp 1677622389
transform 1 0 3524 0 1 3555
box -2 -2 2 2
use M3_M2  M3_M2_2119
timestamp 1677622389
transform 1 0 3564 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1677622389
transform 1 0 3548 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2529
timestamp 1677622389
transform 1 0 3548 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1677622389
transform 1 0 3564 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1677622389
transform 1 0 3540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1677622389
transform 1 0 3572 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2149
timestamp 1677622389
transform 1 0 3596 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1677622389
transform 1 0 3644 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1677622389
transform 1 0 3628 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2531
timestamp 1677622389
transform 1 0 3676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1677622389
transform 1 0 3596 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1677622389
transform 1 0 3628 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2120
timestamp 1677622389
transform 1 0 3692 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2532
timestamp 1677622389
transform 1 0 3692 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2179
timestamp 1677622389
transform 1 0 3724 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2533
timestamp 1677622389
transform 1 0 3724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1677622389
transform 1 0 3740 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1677622389
transform 1 0 3716 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1677622389
transform 1 0 3732 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1677622389
transform 1 0 3740 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1677622389
transform 1 0 3716 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1677622389
transform 1 0 3732 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1677622389
transform 1 0 3764 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1677622389
transform 1 0 3772 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2535
timestamp 1677622389
transform 1 0 3756 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1677622389
transform 1 0 3772 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1677622389
transform 1 0 3788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1677622389
transform 1 0 3756 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1677622389
transform 1 0 3764 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1677622389
transform 1 0 3780 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2228
timestamp 1677622389
transform 1 0 3788 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1677622389
transform 1 0 3756 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1677622389
transform 1 0 3772 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1677622389
transform 1 0 3748 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1677622389
transform 1 0 3780 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2538
timestamp 1677622389
transform 1 0 3804 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2122
timestamp 1677622389
transform 1 0 3852 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1677622389
transform 1 0 3884 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1677622389
transform 1 0 3828 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1677622389
transform 1 0 3868 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1677622389
transform 1 0 3852 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2539
timestamp 1677622389
transform 1 0 3828 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2202
timestamp 1677622389
transform 1 0 3876 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1677622389
transform 1 0 3908 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2646
timestamp 1677622389
transform 1 0 3852 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1677622389
transform 1 0 3908 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2274
timestamp 1677622389
transform 1 0 3828 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1677622389
transform 1 0 3956 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2540
timestamp 1677622389
transform 1 0 3956 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1677622389
transform 1 0 3980 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2260
timestamp 1677622389
transform 1 0 3980 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2649
timestamp 1677622389
transform 1 0 4076 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1677622389
transform 1 0 4084 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2300
timestamp 1677622389
transform 1 0 4076 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1677622389
transform 1 0 4140 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2541
timestamp 1677622389
transform 1 0 4148 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1677622389
transform 1 0 4132 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2229
timestamp 1677622389
transform 1 0 4140 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2677
timestamp 1677622389
transform 1 0 4124 0 1 3505
box -2 -2 2 2
use M3_M2  M3_M2_2319
timestamp 1677622389
transform 1 0 4124 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2675
timestamp 1677622389
transform 1 0 4156 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2275
timestamp 1677622389
transform 1 0 4156 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1677622389
transform 1 0 4188 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2542
timestamp 1677622389
transform 1 0 4188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1677622389
transform 1 0 4180 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1677622389
transform 1 0 4196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1677622389
transform 1 0 4236 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1677622389
transform 1 0 4252 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2276
timestamp 1677622389
transform 1 0 4236 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1677622389
transform 1 0 4276 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2543
timestamp 1677622389
transform 1 0 4284 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2124
timestamp 1677622389
transform 1 0 4348 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1677622389
transform 1 0 4356 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1677622389
transform 1 0 4372 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1677622389
transform 1 0 4388 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1677622389
transform 1 0 4340 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2544
timestamp 1677622389
transform 1 0 4388 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1677622389
transform 1 0 4308 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1677622389
transform 1 0 4340 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2185
timestamp 1677622389
transform 1 0 4428 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1677622389
transform 1 0 4460 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2545
timestamp 1677622389
transform 1 0 4428 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1677622389
transform 1 0 4444 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1677622389
transform 1 0 4452 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1677622389
transform 1 0 4420 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1677622389
transform 1 0 4436 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1677622389
transform 1 0 4452 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1677622389
transform 1 0 4460 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2261
timestamp 1677622389
transform 1 0 4436 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1677622389
transform 1 0 4444 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1677622389
transform 1 0 4500 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1677622389
transform 1 0 4492 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1677622389
transform 1 0 4596 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1677622389
transform 1 0 4548 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1677622389
transform 1 0 4588 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2548
timestamp 1677622389
transform 1 0 4484 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1677622389
transform 1 0 4500 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2206
timestamp 1677622389
transform 1 0 4540 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1677622389
transform 1 0 4556 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1677622389
transform 1 0 4636 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1677622389
transform 1 0 4636 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2550
timestamp 1677622389
transform 1 0 4588 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1677622389
transform 1 0 4604 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1677622389
transform 1 0 4620 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1677622389
transform 1 0 4492 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2230
timestamp 1677622389
transform 1 0 4500 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1677622389
transform 1 0 4628 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2662
timestamp 1677622389
transform 1 0 4508 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1677622389
transform 1 0 4540 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2262
timestamp 1677622389
transform 1 0 4484 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1677622389
transform 1 0 4604 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2664
timestamp 1677622389
transform 1 0 4612 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1677622389
transform 1 0 4628 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2263
timestamp 1677622389
transform 1 0 4540 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1677622389
transform 1 0 4508 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1677622389
transform 1 0 4556 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1677622389
transform 1 0 4620 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1677622389
transform 1 0 4628 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2553
timestamp 1677622389
transform 1 0 4668 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1677622389
transform 1 0 4684 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1677622389
transform 1 0 4708 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2265
timestamp 1677622389
transform 1 0 4708 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2667
timestamp 1677622389
transform 1 0 4780 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2279
timestamp 1677622389
transform 1 0 4780 0 1 3505
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_24
timestamp 1677622389
transform 1 0 24 0 1 3470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_161
timestamp 1677622389
transform 1 0 72 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_188
timestamp 1677622389
transform -1 0 184 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2211
timestamp 1677622389
transform 1 0 184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1677622389
transform 1 0 192 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_104
timestamp 1677622389
transform 1 0 200 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2215
timestamp 1677622389
transform 1 0 240 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1677622389
transform 1 0 248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1677622389
transform 1 0 256 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_102
timestamp 1677622389
transform -1 0 304 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2235
timestamp 1677622389
transform 1 0 304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1677622389
transform 1 0 312 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1677622389
transform 1 0 320 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2237
timestamp 1677622389
transform 1 0 416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1677622389
transform 1 0 424 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_191
timestamp 1677622389
transform -1 0 448 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2239
timestamp 1677622389
transform 1 0 448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1677622389
transform 1 0 456 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_107
timestamp 1677622389
transform 1 0 464 0 -1 3570
box -8 -3 46 105
use BUFX2  BUFX2_14
timestamp 1677622389
transform -1 0 528 0 -1 3570
box -5 -3 28 105
use M3_M2  M3_M2_2320
timestamp 1677622389
transform 1 0 540 0 1 3475
box -3 -3 3 3
use FILL  FILL_2241
timestamp 1677622389
transform 1 0 528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1677622389
transform 1 0 536 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2321
timestamp 1677622389
transform 1 0 580 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_103
timestamp 1677622389
transform 1 0 544 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1677622389
transform 1 0 584 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2243
timestamp 1677622389
transform 1 0 624 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1677622389
transform -1 0 664 0 -1 3570
box -8 -3 40 105
use BUFX2  BUFX2_15
timestamp 1677622389
transform 1 0 664 0 -1 3570
box -5 -3 28 105
use FILL  FILL_2244
timestamp 1677622389
transform 1 0 688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1677622389
transform 1 0 696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1677622389
transform 1 0 704 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2322
timestamp 1677622389
transform 1 0 724 0 1 3475
box -3 -3 3 3
use FILL  FILL_2248
timestamp 1677622389
transform 1 0 712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1677622389
transform 1 0 720 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_25
timestamp 1677622389
transform 1 0 728 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2261
timestamp 1677622389
transform 1 0 752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1677622389
transform 1 0 760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1677622389
transform 1 0 768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1677622389
transform 1 0 776 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2323
timestamp 1677622389
transform 1 0 812 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_104
timestamp 1677622389
transform 1 0 784 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2265
timestamp 1677622389
transform 1 0 824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1677622389
transform 1 0 832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1677622389
transform 1 0 840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1677622389
transform 1 0 848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1677622389
transform 1 0 856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1677622389
transform 1 0 864 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_26
timestamp 1677622389
transform 1 0 872 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2272
timestamp 1677622389
transform 1 0 896 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1677622389
transform 1 0 904 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1677622389
transform 1 0 912 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2283
timestamp 1677622389
transform 1 0 1008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1677622389
transform 1 0 1016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1677622389
transform 1 0 1024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1677622389
transform 1 0 1032 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_27
timestamp 1677622389
transform 1 0 1040 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2290
timestamp 1677622389
transform 1 0 1064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1677622389
transform 1 0 1072 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2324
timestamp 1677622389
transform 1 0 1092 0 1 3475
box -3 -3 3 3
use FILL  FILL_2294
timestamp 1677622389
transform 1 0 1080 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1677622389
transform 1 0 1088 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2301
timestamp 1677622389
transform 1 0 1184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1677622389
transform 1 0 1192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1677622389
transform 1 0 1200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1677622389
transform 1 0 1208 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1677622389
transform 1 0 1216 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2309
timestamp 1677622389
transform 1 0 1248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1677622389
transform 1 0 1256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1677622389
transform 1 0 1264 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_16
timestamp 1677622389
transform -1 0 1296 0 -1 3570
box -5 -3 28 105
use FILL  FILL_2315
timestamp 1677622389
transform 1 0 1296 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1677622389
transform 1 0 1304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1677622389
transform 1 0 1312 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_195
timestamp 1677622389
transform -1 0 1336 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2322
timestamp 1677622389
transform 1 0 1336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1677622389
transform 1 0 1344 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1677622389
transform 1 0 1352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1677622389
transform 1 0 1360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1677622389
transform 1 0 1368 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1677622389
transform 1 0 1376 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2335
timestamp 1677622389
transform 1 0 1408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1677622389
transform 1 0 1416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1677622389
transform 1 0 1424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1677622389
transform 1 0 1432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1677622389
transform 1 0 1440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1677622389
transform 1 0 1448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1677622389
transform 1 0 1456 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1677622389
transform 1 0 1464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1677622389
transform 1 0 1472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1677622389
transform 1 0 1480 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1677622389
transform 1 0 1488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1677622389
transform 1 0 1496 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_105
timestamp 1677622389
transform -1 0 1544 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2347
timestamp 1677622389
transform 1 0 1544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1677622389
transform 1 0 1552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1677622389
transform 1 0 1560 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_196
timestamp 1677622389
transform -1 0 1584 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1677622389
transform -1 0 1600 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2350
timestamp 1677622389
transform 1 0 1600 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1677622389
transform 1 0 1608 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1677622389
transform 1 0 1616 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1677622389
transform 1 0 1624 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_17
timestamp 1677622389
transform -1 0 1656 0 -1 3570
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1677622389
transform -1 0 1680 0 -1 3570
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1677622389
transform -1 0 1704 0 -1 3570
box -5 -3 28 105
use FILL  FILL_2356
timestamp 1677622389
transform 1 0 1704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1677622389
transform 1 0 1712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1677622389
transform 1 0 1720 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_199
timestamp 1677622389
transform -1 0 1744 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2359
timestamp 1677622389
transform 1 0 1744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1677622389
transform 1 0 1752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1677622389
transform 1 0 1760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1677622389
transform 1 0 1768 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_106
timestamp 1677622389
transform 1 0 1776 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2373
timestamp 1677622389
transform 1 0 1816 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1677622389
transform -1 0 1920 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2374
timestamp 1677622389
transform 1 0 1920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1677622389
transform 1 0 1928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1677622389
transform 1 0 1936 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1677622389
transform 1 0 1944 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1677622389
transform 1 0 1952 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1677622389
transform 1 0 1960 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1677622389
transform 1 0 1968 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1677622389
transform 1 0 1976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1677622389
transform 1 0 1984 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1677622389
transform 1 0 1992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1677622389
transform 1 0 2000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1677622389
transform 1 0 2008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1677622389
transform 1 0 2016 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_200
timestamp 1677622389
transform 1 0 2024 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2388
timestamp 1677622389
transform 1 0 2040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1677622389
transform 1 0 2048 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1677622389
transform 1 0 2056 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1677622389
transform 1 0 2064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1677622389
transform 1 0 2072 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1677622389
transform 1 0 2080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1677622389
transform 1 0 2088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1677622389
transform 1 0 2096 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1677622389
transform 1 0 2104 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1677622389
transform 1 0 2112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1677622389
transform 1 0 2120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1677622389
transform 1 0 2128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1677622389
transform 1 0 2136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1677622389
transform 1 0 2144 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_107
timestamp 1677622389
transform 1 0 2152 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2402
timestamp 1677622389
transform 1 0 2192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1677622389
transform 1 0 2200 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_20
timestamp 1677622389
transform 1 0 2208 0 -1 3570
box -5 -3 28 105
use FILL  FILL_2405
timestamp 1677622389
transform 1 0 2232 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1677622389
transform 1 0 2240 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1677622389
transform 1 0 2248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1677622389
transform 1 0 2256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1677622389
transform 1 0 2264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1677622389
transform 1 0 2272 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1677622389
transform 1 0 2280 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1677622389
transform 1 0 2288 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_108
timestamp 1677622389
transform 1 0 2296 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2432
timestamp 1677622389
transform 1 0 2336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1677622389
transform 1 0 2344 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1677622389
transform 1 0 2352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1677622389
transform 1 0 2360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1677622389
transform 1 0 2368 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1677622389
transform -1 0 2472 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2437
timestamp 1677622389
transform 1 0 2472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1677622389
transform 1 0 2480 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1677622389
transform -1 0 2520 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2448
timestamp 1677622389
transform 1 0 2520 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_3
timestamp 1677622389
transform -1 0 2560 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2449
timestamp 1677622389
transform 1 0 2560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1677622389
transform 1 0 2568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1677622389
transform 1 0 2576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1677622389
transform 1 0 2584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1677622389
transform 1 0 2592 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_116
timestamp 1677622389
transform 1 0 2600 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2460
timestamp 1677622389
transform 1 0 2640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1677622389
transform 1 0 2648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1677622389
transform 1 0 2656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1677622389
transform 1 0 2664 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_28
timestamp 1677622389
transform 1 0 2672 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2464
timestamp 1677622389
transform 1 0 2696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1677622389
transform 1 0 2704 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_29
timestamp 1677622389
transform 1 0 2712 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2466
timestamp 1677622389
transform 1 0 2736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1677622389
transform 1 0 2744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1677622389
transform 1 0 2752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1677622389
transform 1 0 2760 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_59
timestamp 1677622389
transform 1 0 2768 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1677622389
transform 1 0 2800 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2482
timestamp 1677622389
transform 1 0 2832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1677622389
transform 1 0 2840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1677622389
transform 1 0 2848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1677622389
transform 1 0 2856 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_31
timestamp 1677622389
transform 1 0 2864 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2486
timestamp 1677622389
transform 1 0 2888 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1677622389
transform 1 0 2896 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1677622389
transform 1 0 2904 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1677622389
transform -1 0 2944 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2491
timestamp 1677622389
transform 1 0 2944 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1677622389
transform 1 0 2952 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1677622389
transform 1 0 2960 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1677622389
transform 1 0 2968 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_206
timestamp 1677622389
transform 1 0 2976 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2495
timestamp 1677622389
transform 1 0 2992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1677622389
transform 1 0 3000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1677622389
transform 1 0 3008 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_109
timestamp 1677622389
transform 1 0 3016 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2498
timestamp 1677622389
transform 1 0 3056 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1677622389
transform 1 0 3064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1677622389
transform 1 0 3072 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_4
timestamp 1677622389
transform -1 0 3112 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2504
timestamp 1677622389
transform 1 0 3112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1677622389
transform 1 0 3120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1677622389
transform 1 0 3128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1677622389
transform 1 0 3136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1677622389
transform 1 0 3144 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_5
timestamp 1677622389
transform 1 0 3152 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2518
timestamp 1677622389
transform 1 0 3184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1677622389
transform 1 0 3192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1677622389
transform 1 0 3200 0 -1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1677622389
transform -1 0 3240 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2521
timestamp 1677622389
transform 1 0 3240 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1677622389
transform 1 0 3248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1677622389
transform 1 0 3256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1677622389
transform 1 0 3264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1677622389
transform 1 0 3272 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_6
timestamp 1677622389
transform 1 0 3280 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2531
timestamp 1677622389
transform 1 0 3312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1677622389
transform 1 0 3320 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_112
timestamp 1677622389
transform -1 0 3368 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2540
timestamp 1677622389
transform 1 0 3368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1677622389
transform 1 0 3376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1677622389
transform 1 0 3384 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1677622389
transform 1 0 3392 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1677622389
transform 1 0 3400 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_117
timestamp 1677622389
transform 1 0 3408 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2553
timestamp 1677622389
transform 1 0 3448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1677622389
transform 1 0 3456 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1677622389
transform 1 0 3464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1677622389
transform 1 0 3472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1677622389
transform 1 0 3480 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1677622389
transform 1 0 3488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1677622389
transform 1 0 3496 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1677622389
transform 1 0 3504 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1677622389
transform 1 0 3512 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1677622389
transform 1 0 3520 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_115
timestamp 1677622389
transform -1 0 3568 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2578
timestamp 1677622389
transform 1 0 3568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1677622389
transform 1 0 3576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1677622389
transform 1 0 3584 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1677622389
transform -1 0 3688 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2581
timestamp 1677622389
transform 1 0 3688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1677622389
transform 1 0 3696 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_116
timestamp 1677622389
transform 1 0 3704 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2583
timestamp 1677622389
transform 1 0 3744 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_118
timestamp 1677622389
transform 1 0 3752 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2596
timestamp 1677622389
transform 1 0 3792 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1677622389
transform 1 0 3800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1677622389
transform 1 0 3808 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1677622389
transform 1 0 3816 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2599
timestamp 1677622389
transform 1 0 3912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1677622389
transform 1 0 3920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1677622389
transform 1 0 3928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1677622389
transform 1 0 3936 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1677622389
transform 1 0 3944 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2609
timestamp 1677622389
transform 1 0 4040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1677622389
transform 1 0 4048 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2325
timestamp 1677622389
transform 1 0 4068 0 1 3475
box -3 -3 3 3
use FILL  FILL_2611
timestamp 1677622389
transform 1 0 4056 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_209
timestamp 1677622389
transform 1 0 4064 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2612
timestamp 1677622389
transform 1 0 4080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1677622389
transform 1 0 4088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1677622389
transform 1 0 4096 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1677622389
transform 1 0 4104 0 -1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1677622389
transform -1 0 4144 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2635
timestamp 1677622389
transform 1 0 4144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1677622389
transform 1 0 4152 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_21
timestamp 1677622389
transform -1 0 4184 0 -1 3570
box -5 -3 28 105
use FILL  FILL_2637
timestamp 1677622389
transform 1 0 4184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1677622389
transform 1 0 4192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1677622389
transform 1 0 4200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1677622389
transform 1 0 4208 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_119
timestamp 1677622389
transform -1 0 4256 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2641
timestamp 1677622389
transform 1 0 4256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1677622389
transform 1 0 4264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1677622389
transform 1 0 4272 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1677622389
transform 1 0 4280 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1677622389
transform 1 0 4288 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1677622389
transform 1 0 4296 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1677622389
transform -1 0 4400 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2647
timestamp 1677622389
transform 1 0 4400 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1677622389
transform 1 0 4408 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_121
timestamp 1677622389
transform -1 0 4456 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2671
timestamp 1677622389
transform 1 0 4456 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_123
timestamp 1677622389
transform 1 0 4464 0 -1 3570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1677622389
transform -1 0 4600 0 -1 3570
box -8 -3 104 105
use OAI22X1  OAI22X1_124
timestamp 1677622389
transform 1 0 4600 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2672
timestamp 1677622389
transform 1 0 4640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1677622389
transform 1 0 4648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1677622389
transform 1 0 4656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1677622389
transform 1 0 4664 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1677622389
transform 1 0 4672 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_213
timestamp 1677622389
transform 1 0 4768 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2676
timestamp 1677622389
transform 1 0 4784 0 -1 3570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_25
timestamp 1677622389
transform 1 0 4843 0 1 3470
box -10 -3 10 3
use M3_M2  M3_M2_2346
timestamp 1677622389
transform 1 0 156 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1677622389
transform 1 0 212 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1677622389
transform 1 0 188 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1677622389
transform 1 0 228 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2686
timestamp 1677622389
transform 1 0 188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1677622389
transform 1 0 220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1677622389
transform 1 0 228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1677622389
transform 1 0 140 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2451
timestamp 1677622389
transform 1 0 220 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1677622389
transform 1 0 268 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1677622389
transform 1 0 284 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2689
timestamp 1677622389
transform 1 0 260 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2404
timestamp 1677622389
transform 1 0 276 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2690
timestamp 1677622389
transform 1 0 284 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1677622389
transform 1 0 268 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1677622389
transform 1 0 276 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1677622389
transform 1 0 292 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2426
timestamp 1677622389
transform 1 0 292 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1677622389
transform 1 0 276 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2691
timestamp 1677622389
transform 1 0 316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1677622389
transform 1 0 324 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2427
timestamp 1677622389
transform 1 0 324 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2692
timestamp 1677622389
transform 1 0 364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1677622389
transform 1 0 420 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1677622389
transform 1 0 340 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1677622389
transform 1 0 380 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1677622389
transform 1 0 420 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1677622389
transform 1 0 404 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2775
timestamp 1677622389
transform 1 0 460 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2383
timestamp 1677622389
transform 1 0 476 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1677622389
transform 1 0 516 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2694
timestamp 1677622389
transform 1 0 476 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1677622389
transform 1 0 516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1677622389
transform 1 0 572 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1677622389
transform 1 0 580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1677622389
transform 1 0 492 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2429
timestamp 1677622389
transform 1 0 524 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1677622389
transform 1 0 628 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2698
timestamp 1677622389
transform 1 0 628 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2357
timestamp 1677622389
transform 1 0 652 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2777
timestamp 1677622389
transform 1 0 644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2430
timestamp 1677622389
transform 1 0 636 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2778
timestamp 1677622389
transform 1 0 668 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2431
timestamp 1677622389
transform 1 0 676 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1677622389
transform 1 0 708 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2699
timestamp 1677622389
transform 1 0 708 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1677622389
transform 1 0 724 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1677622389
transform 1 0 732 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2779
timestamp 1677622389
transform 1 0 716 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2417
timestamp 1677622389
transform 1 0 724 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2780
timestamp 1677622389
transform 1 0 732 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2432
timestamp 1677622389
transform 1 0 716 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1677622389
transform 1 0 756 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1677622389
transform 1 0 748 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1677622389
transform 1 0 796 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1677622389
transform 1 0 812 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1677622389
transform 1 0 812 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2834
timestamp 1677622389
transform 1 0 820 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1677622389
transform 1 0 1012 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2434
timestamp 1677622389
transform 1 0 1012 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2781
timestamp 1677622389
transform 1 0 1044 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2386
timestamp 1677622389
transform 1 0 1156 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2702
timestamp 1677622389
transform 1 0 1156 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1677622389
transform 1 0 1212 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1677622389
transform 1 0 1236 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2326
timestamp 1677622389
transform 1 0 1260 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1677622389
transform 1 0 1252 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2704
timestamp 1677622389
transform 1 0 1260 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1677622389
transform 1 0 1252 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1677622389
transform 1 0 1316 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1677622389
transform 1 0 1324 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2435
timestamp 1677622389
transform 1 0 1324 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2705
timestamp 1677622389
transform 1 0 1420 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1677622389
transform 1 0 1412 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1677622389
transform 1 0 1428 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1677622389
transform 1 0 1460 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2407
timestamp 1677622389
transform 1 0 1492 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1677622389
transform 1 0 1492 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1677622389
transform 1 0 1564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1677622389
transform 1 0 1516 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2436
timestamp 1677622389
transform 1 0 1516 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2708
timestamp 1677622389
transform 1 0 1628 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2338
timestamp 1677622389
transform 1 0 1676 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2709
timestamp 1677622389
transform 1 0 1692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1677622389
transform 1 0 1660 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2437
timestamp 1677622389
transform 1 0 1660 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2710
timestamp 1677622389
transform 1 0 1748 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1677622389
transform 1 0 1772 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2339
timestamp 1677622389
transform 1 0 1804 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1677622389
transform 1 0 1796 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1677622389
transform 1 0 1804 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1677622389
transform 1 0 1836 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1677622389
transform 1 0 1828 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2712
timestamp 1677622389
transform 1 0 1836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1677622389
transform 1 0 1812 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1677622389
transform 1 0 1828 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1677622389
transform 1 0 1844 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2438
timestamp 1677622389
transform 1 0 1828 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2713
timestamp 1677622389
transform 1 0 1868 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1677622389
transform 1 0 1916 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1677622389
transform 1 0 1932 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1677622389
transform 1 0 1964 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2410
timestamp 1677622389
transform 1 0 1972 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2793
timestamp 1677622389
transform 1 0 1948 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1677622389
transform 1 0 1956 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1677622389
transform 1 0 1972 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1677622389
transform 1 0 1980 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2358
timestamp 1677622389
transform 1 0 1996 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1677622389
transform 1 0 2028 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1677622389
transform 1 0 2020 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1677622389
transform 1 0 2012 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2717
timestamp 1677622389
transform 1 0 2012 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1677622389
transform 1 0 2036 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2351
timestamp 1677622389
transform 1 0 2060 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1677622389
transform 1 0 2052 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2797
timestamp 1677622389
transform 1 0 2068 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2439
timestamp 1677622389
transform 1 0 2060 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1677622389
transform 1 0 2108 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2719
timestamp 1677622389
transform 1 0 2092 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1677622389
transform 1 0 2108 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2418
timestamp 1677622389
transform 1 0 2092 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2798
timestamp 1677622389
transform 1 0 2100 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2419
timestamp 1677622389
transform 1 0 2140 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1677622389
transform 1 0 2220 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1677622389
transform 1 0 2244 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2721
timestamp 1677622389
transform 1 0 2332 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1677622389
transform 1 0 2284 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2420
timestamp 1677622389
transform 1 0 2348 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1677622389
transform 1 0 2380 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2722
timestamp 1677622389
transform 1 0 2372 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1677622389
transform 1 0 2380 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2453
timestamp 1677622389
transform 1 0 2332 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1677622389
transform 1 0 2364 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1677622389
transform 1 0 2404 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1677622389
transform 1 0 2404 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2724
timestamp 1677622389
transform 1 0 2404 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1677622389
transform 1 0 2412 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2341
timestamp 1677622389
transform 1 0 2452 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1677622389
transform 1 0 2444 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2801
timestamp 1677622389
transform 1 0 2436 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2455
timestamp 1677622389
transform 1 0 2436 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2725
timestamp 1677622389
transform 1 0 2452 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1677622389
transform 1 0 2476 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2440
timestamp 1677622389
transform 1 0 2476 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1677622389
transform 1 0 2492 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1677622389
transform 1 0 2508 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2726
timestamp 1677622389
transform 1 0 2508 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1677622389
transform 1 0 2516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1677622389
transform 1 0 2532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1677622389
transform 1 0 2524 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2441
timestamp 1677622389
transform 1 0 2532 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1677622389
transform 1 0 2516 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1677622389
transform 1 0 2564 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1677622389
transform 1 0 2556 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2729
timestamp 1677622389
transform 1 0 2564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1677622389
transform 1 0 2564 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2442
timestamp 1677622389
transform 1 0 2564 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1677622389
transform 1 0 2636 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1677622389
transform 1 0 2644 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1677622389
transform 1 0 2604 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2730
timestamp 1677622389
transform 1 0 2604 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2411
timestamp 1677622389
transform 1 0 2620 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2731
timestamp 1677622389
transform 1 0 2660 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1677622389
transform 1 0 2580 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2412
timestamp 1677622389
transform 1 0 2668 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2806
timestamp 1677622389
transform 1 0 2668 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2443
timestamp 1677622389
transform 1 0 2660 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1677622389
transform 1 0 2580 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1677622389
transform 1 0 2708 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1677622389
transform 1 0 2716 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1677622389
transform 1 0 2732 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1677622389
transform 1 0 2772 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2732
timestamp 1677622389
transform 1 0 2732 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1677622389
transform 1 0 2772 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1677622389
transform 1 0 2828 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1677622389
transform 1 0 2836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1677622389
transform 1 0 2748 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2458
timestamp 1677622389
transform 1 0 2748 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2808
timestamp 1677622389
transform 1 0 2844 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1677622389
transform 1 0 2860 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2329
timestamp 1677622389
transform 1 0 2884 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1677622389
transform 1 0 2900 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2681
timestamp 1677622389
transform 1 0 2900 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2421
timestamp 1677622389
transform 1 0 2892 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2835
timestamp 1677622389
transform 1 0 2892 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2330
timestamp 1677622389
transform 1 0 2916 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2809
timestamp 1677622389
transform 1 0 2908 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2371
timestamp 1677622389
transform 1 0 2924 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2737
timestamp 1677622389
transform 1 0 2924 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1677622389
transform 1 0 2980 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1677622389
transform 1 0 3036 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1677622389
transform 1 0 2972 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2444
timestamp 1677622389
transform 1 0 2972 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2811
timestamp 1677622389
transform 1 0 3060 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1677622389
transform 1 0 3148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1677622389
transform 1 0 3180 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1677622389
transform 1 0 3100 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2422
timestamp 1677622389
transform 1 0 3148 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1677622389
transform 1 0 3172 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1677622389
transform 1 0 3100 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1677622389
transform 1 0 3140 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1677622389
transform 1 0 3244 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1677622389
transform 1 0 3260 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2742
timestamp 1677622389
transform 1 0 3244 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1677622389
transform 1 0 3292 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1677622389
transform 1 0 3212 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2461
timestamp 1677622389
transform 1 0 3212 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1677622389
transform 1 0 3284 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2744
timestamp 1677622389
transform 1 0 3348 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1677622389
transform 1 0 3324 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2445
timestamp 1677622389
transform 1 0 3340 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2745
timestamp 1677622389
transform 1 0 3436 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2393
timestamp 1677622389
transform 1 0 3484 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1677622389
transform 1 0 3476 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2746
timestamp 1677622389
transform 1 0 3492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1677622389
transform 1 0 3508 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1677622389
transform 1 0 3516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1677622389
transform 1 0 3484 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2425
timestamp 1677622389
transform 1 0 3516 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2682
timestamp 1677622389
transform 1 0 3540 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1677622389
transform 1 0 3596 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2373
timestamp 1677622389
transform 1 0 3620 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2749
timestamp 1677622389
transform 1 0 3684 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2331
timestamp 1677622389
transform 1 0 3700 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2817
timestamp 1677622389
transform 1 0 3708 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2332
timestamp 1677622389
transform 1 0 3724 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1677622389
transform 1 0 3812 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2750
timestamp 1677622389
transform 1 0 3796 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1677622389
transform 1 0 3812 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1677622389
transform 1 0 3828 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1677622389
transform 1 0 3804 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1677622389
transform 1 0 3820 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2446
timestamp 1677622389
transform 1 0 3804 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1677622389
transform 1 0 3836 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1677622389
transform 1 0 3860 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2820
timestamp 1677622389
transform 1 0 3892 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2334
timestamp 1677622389
transform 1 0 3916 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1677622389
transform 1 0 3908 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2753
timestamp 1677622389
transform 1 0 3932 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2414
timestamp 1677622389
transform 1 0 3988 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2821
timestamp 1677622389
transform 1 0 3908 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1677622389
transform 1 0 3932 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1677622389
transform 1 0 4020 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2754
timestamp 1677622389
transform 1 0 4020 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1677622389
transform 1 0 4052 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1677622389
transform 1 0 4068 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1677622389
transform 1 0 4084 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2345
timestamp 1677622389
transform 1 0 4156 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1677622389
transform 1 0 4148 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1677622389
transform 1 0 4140 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2679
timestamp 1677622389
transform 1 0 4156 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1677622389
transform 1 0 4148 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2376
timestamp 1677622389
transform 1 0 4164 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2756
timestamp 1677622389
transform 1 0 4164 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2396
timestamp 1677622389
transform 1 0 4180 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2685
timestamp 1677622389
transform 1 0 4196 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2377
timestamp 1677622389
transform 1 0 4220 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1677622389
transform 1 0 4236 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2757
timestamp 1677622389
transform 1 0 4220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1677622389
transform 1 0 4236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1677622389
transform 1 0 4212 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2398
timestamp 1677622389
transform 1 0 4252 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2759
timestamp 1677622389
transform 1 0 4284 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1677622389
transform 1 0 4292 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1677622389
transform 1 0 4308 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1677622389
transform 1 0 4316 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2463
timestamp 1677622389
transform 1 0 4356 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1677622389
transform 1 0 4372 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2399
timestamp 1677622389
transform 1 0 4388 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2760
timestamp 1677622389
transform 1 0 4388 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1677622389
transform 1 0 4404 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2354
timestamp 1677622389
transform 1 0 4428 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1677622389
transform 1 0 4436 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2762
timestamp 1677622389
transform 1 0 4428 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1677622389
transform 1 0 4436 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2448
timestamp 1677622389
transform 1 0 4436 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2763
timestamp 1677622389
transform 1 0 4452 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2355
timestamp 1677622389
transform 1 0 4492 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1677622389
transform 1 0 4516 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1677622389
transform 1 0 4508 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2764
timestamp 1677622389
transform 1 0 4492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1677622389
transform 1 0 4516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1677622389
transform 1 0 4484 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1677622389
transform 1 0 4492 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1677622389
transform 1 0 4508 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2356
timestamp 1677622389
transform 1 0 4532 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2831
timestamp 1677622389
transform 1 0 4532 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2402
timestamp 1677622389
transform 1 0 4588 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2766
timestamp 1677622389
transform 1 0 4588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1677622389
transform 1 0 4564 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2449
timestamp 1677622389
transform 1 0 4636 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1677622389
transform 1 0 4564 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1677622389
transform 1 0 4660 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2767
timestamp 1677622389
transform 1 0 4660 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2450
timestamp 1677622389
transform 1 0 4660 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2768
timestamp 1677622389
transform 1 0 4676 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1677622389
transform 1 0 4756 0 1 3405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_26
timestamp 1677622389
transform 1 0 48 0 1 3370
box -10 -3 10 3
use FILL  FILL_2677
timestamp 1677622389
transform 1 0 72 0 1 3370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1677622389
transform 1 0 80 0 1 3370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1677622389
transform 1 0 88 0 1 3370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1677622389
transform 1 0 96 0 1 3370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1677622389
transform 1 0 104 0 1 3370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1677622389
transform 1 0 112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1677622389
transform 1 0 120 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2465
timestamp 1677622389
transform 1 0 228 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_186
timestamp 1677622389
transform 1 0 128 0 1 3370
box -8 -3 104 105
use FILL  FILL_2685
timestamp 1677622389
transform 1 0 224 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_214
timestamp 1677622389
transform -1 0 248 0 1 3370
box -9 -3 26 105
use FILL  FILL_2686
timestamp 1677622389
transform 1 0 248 0 1 3370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1677622389
transform 1 0 256 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2466
timestamp 1677622389
transform 1 0 284 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1677622389
transform 1 0 300 0 1 3375
box -3 -3 3 3
use AOI22X1  AOI22X1_122
timestamp 1677622389
transform -1 0 304 0 1 3370
box -8 -3 46 105
use FILL  FILL_2688
timestamp 1677622389
transform 1 0 304 0 1 3370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1677622389
transform 1 0 312 0 1 3370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1677622389
transform 1 0 320 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1677622389
transform 1 0 328 0 1 3370
box -8 -3 104 105
use FILL  FILL_2691
timestamp 1677622389
transform 1 0 424 0 1 3370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1677622389
transform 1 0 432 0 1 3370
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1677622389
transform 1 0 440 0 1 3370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1677622389
transform 1 0 448 0 1 3370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1677622389
transform 1 0 456 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2468
timestamp 1677622389
transform 1 0 484 0 1 3375
box -3 -3 3 3
use INVX2  INVX2_217
timestamp 1677622389
transform 1 0 464 0 1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1677622389
transform 1 0 480 0 1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2469
timestamp 1677622389
transform 1 0 588 0 1 3375
box -3 -3 3 3
use FILL  FILL_2710
timestamp 1677622389
transform 1 0 576 0 1 3370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1677622389
transform 1 0 584 0 1 3370
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1677622389
transform 1 0 592 0 1 3370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1677622389
transform 1 0 600 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_7
timestamp 1677622389
transform -1 0 640 0 1 3370
box -8 -3 40 105
use FILL  FILL_2714
timestamp 1677622389
transform 1 0 640 0 1 3370
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1677622389
transform 1 0 648 0 1 3370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1677622389
transform 1 0 656 0 1 3370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1677622389
transform 1 0 664 0 1 3370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1677622389
transform 1 0 672 0 1 3370
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1677622389
transform 1 0 680 0 1 3370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1677622389
transform 1 0 688 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_126
timestamp 1677622389
transform 1 0 696 0 1 3370
box -8 -3 46 105
use FILL  FILL_2731
timestamp 1677622389
transform 1 0 736 0 1 3370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1677622389
transform 1 0 744 0 1 3370
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1677622389
transform 1 0 752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1677622389
transform 1 0 760 0 1 3370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1677622389
transform 1 0 768 0 1 3370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1677622389
transform 1 0 776 0 1 3370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1677622389
transform 1 0 784 0 1 3370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1677622389
transform 1 0 792 0 1 3370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1677622389
transform 1 0 800 0 1 3370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1677622389
transform 1 0 808 0 1 3370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1677622389
transform 1 0 816 0 1 3370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1677622389
transform 1 0 824 0 1 3370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1677622389
transform 1 0 832 0 1 3370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1677622389
transform 1 0 840 0 1 3370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1677622389
transform 1 0 848 0 1 3370
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1677622389
transform 1 0 856 0 1 3370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1677622389
transform 1 0 864 0 1 3370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1677622389
transform 1 0 872 0 1 3370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1677622389
transform 1 0 880 0 1 3370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1677622389
transform 1 0 888 0 1 3370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1677622389
transform 1 0 896 0 1 3370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1677622389
transform 1 0 904 0 1 3370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1677622389
transform 1 0 912 0 1 3370
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1677622389
transform 1 0 920 0 1 3370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1677622389
transform 1 0 928 0 1 3370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1677622389
transform 1 0 936 0 1 3370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1677622389
transform 1 0 944 0 1 3370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1677622389
transform 1 0 952 0 1 3370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1677622389
transform 1 0 960 0 1 3370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1677622389
transform 1 0 968 0 1 3370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1677622389
transform 1 0 976 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_32
timestamp 1677622389
transform 1 0 984 0 1 3370
box -8 -3 32 105
use FILL  FILL_2781
timestamp 1677622389
transform 1 0 1008 0 1 3370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1677622389
transform 1 0 1016 0 1 3370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1677622389
transform 1 0 1024 0 1 3370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1677622389
transform 1 0 1032 0 1 3370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1677622389
transform 1 0 1040 0 1 3370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1677622389
transform 1 0 1048 0 1 3370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1677622389
transform 1 0 1056 0 1 3370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1677622389
transform 1 0 1064 0 1 3370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1677622389
transform 1 0 1072 0 1 3370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1677622389
transform 1 0 1080 0 1 3370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1677622389
transform 1 0 1088 0 1 3370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1677622389
transform 1 0 1096 0 1 3370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1677622389
transform 1 0 1104 0 1 3370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1677622389
transform 1 0 1112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1677622389
transform 1 0 1120 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2470
timestamp 1677622389
transform 1 0 1140 0 1 3375
box -3 -3 3 3
use FILL  FILL_2809
timestamp 1677622389
transform 1 0 1128 0 1 3370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1677622389
transform 1 0 1136 0 1 3370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1677622389
transform 1 0 1144 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1677622389
transform -1 0 1248 0 1 3370
box -8 -3 104 105
use FILL  FILL_2814
timestamp 1677622389
transform 1 0 1248 0 1 3370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1677622389
transform 1 0 1256 0 1 3370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1677622389
transform 1 0 1264 0 1 3370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1677622389
transform 1 0 1272 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_63
timestamp 1677622389
transform 1 0 1280 0 1 3370
box -8 -3 34 105
use FILL  FILL_2833
timestamp 1677622389
transform 1 0 1312 0 1 3370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1677622389
transform 1 0 1320 0 1 3370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1677622389
transform 1 0 1328 0 1 3370
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1677622389
transform 1 0 1336 0 1 3370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1677622389
transform 1 0 1344 0 1 3370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1677622389
transform 1 0 1352 0 1 3370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1677622389
transform 1 0 1360 0 1 3370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1677622389
transform 1 0 1368 0 1 3370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1677622389
transform 1 0 1376 0 1 3370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1677622389
transform 1 0 1384 0 1 3370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1677622389
transform 1 0 1392 0 1 3370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1677622389
transform 1 0 1400 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_127
timestamp 1677622389
transform -1 0 1448 0 1 3370
box -8 -3 46 105
use FILL  FILL_2850
timestamp 1677622389
transform 1 0 1448 0 1 3370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1677622389
transform 1 0 1456 0 1 3370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1677622389
transform 1 0 1464 0 1 3370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1677622389
transform 1 0 1472 0 1 3370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1677622389
transform 1 0 1480 0 1 3370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1677622389
transform 1 0 1488 0 1 3370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1677622389
transform 1 0 1496 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_194
timestamp 1677622389
transform 1 0 1504 0 1 3370
box -8 -3 104 105
use FILL  FILL_2862
timestamp 1677622389
transform 1 0 1600 0 1 3370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1677622389
transform 1 0 1608 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_221
timestamp 1677622389
transform 1 0 1616 0 1 3370
box -9 -3 26 105
use FILL  FILL_2878
timestamp 1677622389
transform 1 0 1632 0 1 3370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1677622389
transform 1 0 1640 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2471
timestamp 1677622389
transform 1 0 1668 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1677622389
transform 1 0 1748 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_195
timestamp 1677622389
transform 1 0 1648 0 1 3370
box -8 -3 104 105
use FILL  FILL_2884
timestamp 1677622389
transform 1 0 1744 0 1 3370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1677622389
transform 1 0 1752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1677622389
transform 1 0 1760 0 1 3370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1677622389
transform 1 0 1768 0 1 3370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1677622389
transform 1 0 1776 0 1 3370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1677622389
transform 1 0 1784 0 1 3370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1677622389
transform 1 0 1792 0 1 3370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1677622389
transform 1 0 1800 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_128
timestamp 1677622389
transform 1 0 1808 0 1 3370
box -8 -3 46 105
use FILL  FILL_2903
timestamp 1677622389
transform 1 0 1848 0 1 3370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1677622389
transform 1 0 1856 0 1 3370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1677622389
transform 1 0 1864 0 1 3370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1677622389
transform 1 0 1872 0 1 3370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1677622389
transform 1 0 1880 0 1 3370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1677622389
transform 1 0 1888 0 1 3370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1677622389
transform 1 0 1896 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_223
timestamp 1677622389
transform -1 0 1920 0 1 3370
box -9 -3 26 105
use FILL  FILL_2910
timestamp 1677622389
transform 1 0 1920 0 1 3370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1677622389
transform 1 0 1928 0 1 3370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1677622389
transform 1 0 1936 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_128
timestamp 1677622389
transform 1 0 1944 0 1 3370
box -8 -3 46 105
use FILL  FILL_2917
timestamp 1677622389
transform 1 0 1984 0 1 3370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1677622389
transform 1 0 1992 0 1 3370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1677622389
transform 1 0 2000 0 1 3370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1677622389
transform 1 0 2008 0 1 3370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1677622389
transform 1 0 2016 0 1 3370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1677622389
transform 1 0 2024 0 1 3370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1677622389
transform 1 0 2032 0 1 3370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1677622389
transform 1 0 2040 0 1 3370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1677622389
transform 1 0 2048 0 1 3370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1677622389
transform 1 0 2056 0 1 3370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1677622389
transform 1 0 2064 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_129
timestamp 1677622389
transform 1 0 2072 0 1 3370
box -8 -3 46 105
use FILL  FILL_2928
timestamp 1677622389
transform 1 0 2112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1677622389
transform 1 0 2120 0 1 3370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1677622389
transform 1 0 2128 0 1 3370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1677622389
transform 1 0 2136 0 1 3370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1677622389
transform 1 0 2144 0 1 3370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1677622389
transform 1 0 2152 0 1 3370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1677622389
transform 1 0 2160 0 1 3370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1677622389
transform 1 0 2168 0 1 3370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1677622389
transform 1 0 2176 0 1 3370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1677622389
transform 1 0 2184 0 1 3370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1677622389
transform 1 0 2192 0 1 3370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1677622389
transform 1 0 2200 0 1 3370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1677622389
transform 1 0 2208 0 1 3370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1677622389
transform 1 0 2216 0 1 3370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1677622389
transform 1 0 2224 0 1 3370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1677622389
transform 1 0 2232 0 1 3370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1677622389
transform 1 0 2240 0 1 3370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1677622389
transform 1 0 2248 0 1 3370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1677622389
transform 1 0 2256 0 1 3370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1677622389
transform 1 0 2264 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_200
timestamp 1677622389
transform 1 0 2272 0 1 3370
box -8 -3 104 105
use FILL  FILL_2951
timestamp 1677622389
transform 1 0 2368 0 1 3370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1677622389
transform 1 0 2376 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2473
timestamp 1677622389
transform 1 0 2404 0 1 3375
box -3 -3 3 3
use AND2X2  AND2X2_8
timestamp 1677622389
transform -1 0 2416 0 1 3370
box -8 -3 40 105
use FILL  FILL_2953
timestamp 1677622389
transform 1 0 2416 0 1 3370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1677622389
transform 1 0 2424 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_226
timestamp 1677622389
transform 1 0 2432 0 1 3370
box -9 -3 26 105
use FILL  FILL_2955
timestamp 1677622389
transform 1 0 2448 0 1 3370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1677622389
transform 1 0 2456 0 1 3370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1677622389
transform 1 0 2464 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1677622389
transform 1 0 2472 0 1 3370
box -9 -3 26 105
use FILL  FILL_2958
timestamp 1677622389
transform 1 0 2488 0 1 3370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1677622389
transform 1 0 2496 0 1 3370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1677622389
transform 1 0 2504 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_131
timestamp 1677622389
transform 1 0 2512 0 1 3370
box -8 -3 46 105
use FILL  FILL_2972
timestamp 1677622389
transform 1 0 2552 0 1 3370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1677622389
transform 1 0 2560 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1677622389
transform 1 0 2568 0 1 3370
box -8 -3 104 105
use FILL  FILL_2974
timestamp 1677622389
transform 1 0 2664 0 1 3370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1677622389
transform 1 0 2672 0 1 3370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1677622389
transform 1 0 2680 0 1 3370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1677622389
transform 1 0 2688 0 1 3370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1677622389
transform 1 0 2696 0 1 3370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1677622389
transform 1 0 2704 0 1 3370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1677622389
transform 1 0 2712 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_230
timestamp 1677622389
transform 1 0 2720 0 1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_204
timestamp 1677622389
transform 1 0 2736 0 1 3370
box -8 -3 104 105
use FILL  FILL_2987
timestamp 1677622389
transform 1 0 2832 0 1 3370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1677622389
transform 1 0 2840 0 1 3370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1677622389
transform 1 0 2848 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1677622389
transform 1 0 2856 0 1 3370
box -8 -3 34 105
use FILL  FILL_2994
timestamp 1677622389
transform 1 0 2888 0 1 3370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1677622389
transform 1 0 2896 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_34
timestamp 1677622389
transform 1 0 2904 0 1 3370
box -8 -3 32 105
use FILL  FILL_3002
timestamp 1677622389
transform 1 0 2928 0 1 3370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1677622389
transform 1 0 2936 0 1 3370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1677622389
transform 1 0 2944 0 1 3370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1677622389
transform 1 0 2952 0 1 3370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1677622389
transform 1 0 2960 0 1 3370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1677622389
transform 1 0 2968 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1677622389
transform -1 0 3072 0 1 3370
box -8 -3 104 105
use FILL  FILL_3008
timestamp 1677622389
transform 1 0 3072 0 1 3370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1677622389
transform 1 0 3080 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_207
timestamp 1677622389
transform 1 0 3088 0 1 3370
box -8 -3 104 105
use FILL  FILL_3010
timestamp 1677622389
transform 1 0 3184 0 1 3370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1677622389
transform 1 0 3192 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1677622389
transform 1 0 3200 0 1 3370
box -8 -3 104 105
use FILL  FILL_3027
timestamp 1677622389
transform 1 0 3296 0 1 3370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1677622389
transform 1 0 3304 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1677622389
transform 1 0 3312 0 1 3370
box -8 -3 104 105
use FILL  FILL_3036
timestamp 1677622389
transform 1 0 3408 0 1 3370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1677622389
transform 1 0 3416 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_233
timestamp 1677622389
transform 1 0 3424 0 1 3370
box -9 -3 26 105
use FILL  FILL_3038
timestamp 1677622389
transform 1 0 3440 0 1 3370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1677622389
transform 1 0 3448 0 1 3370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1677622389
transform 1 0 3456 0 1 3370
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1677622389
transform 1 0 3464 0 1 3370
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1677622389
transform 1 0 3472 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2474
timestamp 1677622389
transform 1 0 3492 0 1 3375
box -3 -3 3 3
use AND2X2  AND2X2_9
timestamp 1677622389
transform 1 0 3480 0 1 3370
box -8 -3 40 105
use FILL  FILL_3055
timestamp 1677622389
transform 1 0 3512 0 1 3370
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1677622389
transform 1 0 3520 0 1 3370
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1677622389
transform 1 0 3528 0 1 3370
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1677622389
transform 1 0 3536 0 1 3370
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1677622389
transform 1 0 3544 0 1 3370
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1677622389
transform 1 0 3552 0 1 3370
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1677622389
transform 1 0 3560 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_234
timestamp 1677622389
transform -1 0 3584 0 1 3370
box -9 -3 26 105
use FILL  FILL_3064
timestamp 1677622389
transform 1 0 3584 0 1 3370
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1677622389
transform 1 0 3592 0 1 3370
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1677622389
transform 1 0 3600 0 1 3370
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1677622389
transform 1 0 3608 0 1 3370
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1677622389
transform 1 0 3616 0 1 3370
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1677622389
transform 1 0 3624 0 1 3370
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1677622389
transform 1 0 3632 0 1 3370
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1677622389
transform 1 0 3640 0 1 3370
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1677622389
transform 1 0 3648 0 1 3370
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1677622389
transform 1 0 3656 0 1 3370
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1677622389
transform 1 0 3664 0 1 3370
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1677622389
transform 1 0 3672 0 1 3370
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1677622389
transform 1 0 3680 0 1 3370
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1677622389
transform 1 0 3688 0 1 3370
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1677622389
transform 1 0 3696 0 1 3370
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1677622389
transform 1 0 3704 0 1 3370
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1677622389
transform 1 0 3712 0 1 3370
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1677622389
transform 1 0 3720 0 1 3370
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1677622389
transform 1 0 3728 0 1 3370
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1677622389
transform 1 0 3736 0 1 3370
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1677622389
transform 1 0 3744 0 1 3370
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1677622389
transform 1 0 3752 0 1 3370
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1677622389
transform 1 0 3760 0 1 3370
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1677622389
transform 1 0 3768 0 1 3370
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1677622389
transform 1 0 3776 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_131
timestamp 1677622389
transform 1 0 3784 0 1 3370
box -8 -3 46 105
use FILL  FILL_3099
timestamp 1677622389
transform 1 0 3824 0 1 3370
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1677622389
transform 1 0 3832 0 1 3370
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1677622389
transform 1 0 3840 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_235
timestamp 1677622389
transform -1 0 3864 0 1 3370
box -9 -3 26 105
use FILL  FILL_3109
timestamp 1677622389
transform 1 0 3864 0 1 3370
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1677622389
transform 1 0 3872 0 1 3370
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1677622389
transform 1 0 3880 0 1 3370
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1677622389
transform 1 0 3888 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1677622389
transform 1 0 3896 0 1 3370
box -8 -3 104 105
use FILL  FILL_3113
timestamp 1677622389
transform 1 0 3992 0 1 3370
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1677622389
transform 1 0 4000 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_236
timestamp 1677622389
transform 1 0 4008 0 1 3370
box -9 -3 26 105
use FILL  FILL_3115
timestamp 1677622389
transform 1 0 4024 0 1 3370
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1677622389
transform 1 0 4032 0 1 3370
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1677622389
transform 1 0 4040 0 1 3370
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1677622389
transform 1 0 4048 0 1 3370
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1677622389
transform -1 0 4088 0 1 3370
box -8 -3 40 105
use FILL  FILL_3119
timestamp 1677622389
transform 1 0 4088 0 1 3370
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1677622389
transform 1 0 4096 0 1 3370
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1677622389
transform 1 0 4104 0 1 3370
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1677622389
transform 1 0 4112 0 1 3370
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1677622389
transform 1 0 4120 0 1 3370
box -8 -3 16 105
use NAND3X1  NAND3X1_17
timestamp 1677622389
transform -1 0 4160 0 1 3370
box -8 -3 40 105
use FILL  FILL_3130
timestamp 1677622389
transform 1 0 4160 0 1 3370
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1677622389
transform 1 0 4168 0 1 3370
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1677622389
transform 1 0 4176 0 1 3370
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1677622389
transform 1 0 4184 0 1 3370
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1677622389
transform 1 0 4192 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_134
timestamp 1677622389
transform -1 0 4240 0 1 3370
box -8 -3 46 105
use FILL  FILL_3135
timestamp 1677622389
transform 1 0 4240 0 1 3370
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1677622389
transform 1 0 4248 0 1 3370
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1677622389
transform 1 0 4256 0 1 3370
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1677622389
transform 1 0 4264 0 1 3370
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1677622389
transform 1 0 4272 0 1 3370
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1677622389
transform 1 0 4280 0 1 3370
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1677622389
transform 1 0 4288 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_239
timestamp 1677622389
transform -1 0 4312 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1677622389
transform 1 0 4312 0 1 3370
box -9 -3 26 105
use FILL  FILL_3149
timestamp 1677622389
transform 1 0 4328 0 1 3370
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1677622389
transform 1 0 4336 0 1 3370
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1677622389
transform 1 0 4344 0 1 3370
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1677622389
transform 1 0 4352 0 1 3370
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1677622389
transform 1 0 4360 0 1 3370
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1677622389
transform 1 0 4368 0 1 3370
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1677622389
transform 1 0 4376 0 1 3370
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1677622389
transform 1 0 4384 0 1 3370
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1677622389
transform 1 0 4392 0 1 3370
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1677622389
transform 1 0 4400 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2475
timestamp 1677622389
transform 1 0 4420 0 1 3375
box -3 -3 3 3
use AOI22X1  AOI22X1_135
timestamp 1677622389
transform -1 0 4448 0 1 3370
box -8 -3 46 105
use FILL  FILL_3162
timestamp 1677622389
transform 1 0 4448 0 1 3370
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1677622389
transform 1 0 4456 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_25
timestamp 1677622389
transform 1 0 4464 0 1 3370
box -5 -3 28 105
use M3_M2  M3_M2_2476
timestamp 1677622389
transform 1 0 4532 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_132
timestamp 1677622389
transform 1 0 4488 0 1 3370
box -8 -3 46 105
use FILL  FILL_3164
timestamp 1677622389
transform 1 0 4528 0 1 3370
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1677622389
transform 1 0 4536 0 1 3370
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1677622389
transform 1 0 4544 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2477
timestamp 1677622389
transform 1 0 4572 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1677622389
transform 1 0 4620 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_217
timestamp 1677622389
transform 1 0 4552 0 1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2479
timestamp 1677622389
transform 1 0 4676 0 1 3375
box -3 -3 3 3
use INVX2  INVX2_241
timestamp 1677622389
transform 1 0 4648 0 1 3370
box -9 -3 26 105
use FILL  FILL_3176
timestamp 1677622389
transform 1 0 4664 0 1 3370
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1677622389
transform 1 0 4672 0 1 3370
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1677622389
transform 1 0 4680 0 1 3370
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1677622389
transform 1 0 4688 0 1 3370
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1677622389
transform 1 0 4696 0 1 3370
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1677622389
transform 1 0 4704 0 1 3370
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1677622389
transform 1 0 4712 0 1 3370
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1677622389
transform 1 0 4720 0 1 3370
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1677622389
transform 1 0 4728 0 1 3370
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1677622389
transform 1 0 4736 0 1 3370
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1677622389
transform 1 0 4744 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_242
timestamp 1677622389
transform 1 0 4752 0 1 3370
box -9 -3 26 105
use FILL  FILL_3187
timestamp 1677622389
transform 1 0 4768 0 1 3370
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1677622389
transform 1 0 4776 0 1 3370
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1677622389
transform 1 0 4784 0 1 3370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_27
timestamp 1677622389
transform 1 0 4819 0 1 3370
box -10 -3 10 3
use M3_M2  M3_M2_2509
timestamp 1677622389
transform 1 0 172 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2838
timestamp 1677622389
transform 1 0 92 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1677622389
transform 1 0 140 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1677622389
transform 1 0 172 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1677622389
transform 1 0 180 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2585
timestamp 1677622389
transform 1 0 140 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1677622389
transform 1 0 180 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2839
timestamp 1677622389
transform 1 0 204 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2587
timestamp 1677622389
transform 1 0 204 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2840
timestamp 1677622389
transform 1 0 220 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2493
timestamp 1677622389
transform 1 0 260 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1677622389
transform 1 0 268 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2841
timestamp 1677622389
transform 1 0 252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1677622389
transform 1 0 268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1677622389
transform 1 0 244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1677622389
transform 1 0 252 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2920
timestamp 1677622389
transform 1 0 260 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2480
timestamp 1677622389
transform 1 0 340 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1677622389
transform 1 0 316 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1677622389
transform 1 0 332 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2921
timestamp 1677622389
transform 1 0 300 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1677622389
transform 1 0 316 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1677622389
transform 1 0 332 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2588
timestamp 1677622389
transform 1 0 316 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1677622389
transform 1 0 332 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1677622389
transform 1 0 308 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1677622389
transform 1 0 348 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2843
timestamp 1677622389
transform 1 0 348 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1677622389
transform 1 0 356 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2589
timestamp 1677622389
transform 1 0 356 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1677622389
transform 1 0 396 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2845
timestamp 1677622389
transform 1 0 380 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1677622389
transform 1 0 396 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1677622389
transform 1 0 404 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1677622389
transform 1 0 364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1677622389
transform 1 0 372 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1677622389
transform 1 0 388 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2590
timestamp 1677622389
transform 1 0 388 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1677622389
transform 1 0 372 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1677622389
transform 1 0 428 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1677622389
transform 1 0 476 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1677622389
transform 1 0 476 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2927
timestamp 1677622389
transform 1 0 436 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1677622389
transform 1 0 444 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1677622389
transform 1 0 460 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1677622389
transform 1 0 476 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1677622389
transform 1 0 484 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2591
timestamp 1677622389
transform 1 0 436 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1677622389
transform 1 0 492 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1677622389
transform 1 0 484 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1677622389
transform 1 0 516 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2848
timestamp 1677622389
transform 1 0 516 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1677622389
transform 1 0 524 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2544
timestamp 1677622389
transform 1 0 548 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2932
timestamp 1677622389
transform 1 0 532 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1677622389
transform 1 0 548 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2515
timestamp 1677622389
transform 1 0 572 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2850
timestamp 1677622389
transform 1 0 572 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2593
timestamp 1677622389
transform 1 0 572 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1677622389
transform 1 0 588 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2851
timestamp 1677622389
transform 1 0 588 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1677622389
transform 1 0 612 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1677622389
transform 1 0 668 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2594
timestamp 1677622389
transform 1 0 668 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2852
timestamp 1677622389
transform 1 0 684 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2516
timestamp 1677622389
transform 1 0 756 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2936
timestamp 1677622389
transform 1 0 796 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2621
timestamp 1677622389
transform 1 0 804 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2853
timestamp 1677622389
transform 1 0 820 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1677622389
transform 1 0 908 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1677622389
transform 1 0 860 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1677622389
transform 1 0 900 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2595
timestamp 1677622389
transform 1 0 860 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1677622389
transform 1 0 820 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2939
timestamp 1677622389
transform 1 0 916 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1677622389
transform 1 0 924 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1677622389
transform 1 0 916 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2855
timestamp 1677622389
transform 1 0 948 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1677622389
transform 1 0 1028 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2940
timestamp 1677622389
transform 1 0 1044 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1677622389
transform 1 0 1100 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1677622389
transform 1 0 1092 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1677622389
transform 1 0 1108 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1677622389
transform 1 0 1156 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1677622389
transform 1 0 1188 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1677622389
transform 1 0 1212 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1677622389
transform 1 0 1220 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2624
timestamp 1677622389
transform 1 0 1236 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1677622389
transform 1 0 1292 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2857
timestamp 1677622389
transform 1 0 1284 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2566
timestamp 1677622389
transform 1 0 1284 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2947
timestamp 1677622389
transform 1 0 1292 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2653
timestamp 1677622389
transform 1 0 1292 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_2858
timestamp 1677622389
transform 1 0 1316 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1677622389
transform 1 0 1324 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1677622389
transform 1 0 1364 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1677622389
transform 1 0 1412 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2597
timestamp 1677622389
transform 1 0 1412 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1677622389
transform 1 0 1364 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1677622389
transform 1 0 1404 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1677622389
transform 1 0 1372 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1677622389
transform 1 0 1468 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2949
timestamp 1677622389
transform 1 0 1484 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2627
timestamp 1677622389
transform 1 0 1516 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1677622389
transform 1 0 1532 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1677622389
transform 1 0 1588 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1677622389
transform 1 0 1628 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1677622389
transform 1 0 1676 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2860
timestamp 1677622389
transform 1 0 1668 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1677622389
transform 1 0 1676 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1677622389
transform 1 0 1684 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2545
timestamp 1677622389
transform 1 0 1756 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2951
timestamp 1677622389
transform 1 0 1748 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1677622389
transform 1 0 1756 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2518
timestamp 1677622389
transform 1 0 1772 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1677622389
transform 1 0 1780 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2862
timestamp 1677622389
transform 1 0 1796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1677622389
transform 1 0 1804 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2569
timestamp 1677622389
transform 1 0 1804 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1677622389
transform 1 0 1804 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1677622389
transform 1 0 1892 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1677622389
transform 1 0 1924 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1677622389
transform 1 0 1916 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2864
timestamp 1677622389
transform 1 0 1916 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1677622389
transform 1 0 1828 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1677622389
transform 1 0 1836 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1677622389
transform 1 0 1828 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1677622389
transform 1 0 1828 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1677622389
transform 1 0 1844 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2955
timestamp 1677622389
transform 1 0 1868 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2600
timestamp 1677622389
transform 1 0 1868 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1677622389
transform 1 0 1876 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1677622389
transform 1 0 1932 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1677622389
transform 1 0 1956 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2865
timestamp 1677622389
transform 1 0 1956 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2483
timestamp 1677622389
transform 1 0 2116 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1677622389
transform 1 0 2052 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1677622389
transform 1 0 2164 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1677622389
transform 1 0 2148 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2866
timestamp 1677622389
transform 1 0 2052 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2547
timestamp 1677622389
transform 1 0 2132 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2867
timestamp 1677622389
transform 1 0 2148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1677622389
transform 1 0 2236 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1677622389
transform 1 0 1988 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1677622389
transform 1 0 2036 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1677622389
transform 1 0 2084 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1677622389
transform 1 0 2004 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1677622389
transform 1 0 2100 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1677622389
transform 1 0 2124 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2959
timestamp 1677622389
transform 1 0 2132 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2644
timestamp 1677622389
transform 1 0 2068 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1677622389
transform 1 0 2148 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2960
timestamp 1677622389
transform 1 0 2188 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1677622389
transform 1 0 2228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1677622389
transform 1 0 2236 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2601
timestamp 1677622389
transform 1 0 2188 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1677622389
transform 1 0 2236 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1677622389
transform 1 0 2284 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1677622389
transform 1 0 2284 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1677622389
transform 1 0 2300 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2869
timestamp 1677622389
transform 1 0 2292 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2549
timestamp 1677622389
transform 1 0 2324 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2870
timestamp 1677622389
transform 1 0 2332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1677622389
transform 1 0 2308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1677622389
transform 1 0 2324 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2603
timestamp 1677622389
transform 1 0 2332 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2871
timestamp 1677622389
transform 1 0 2348 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1677622389
transform 1 0 2356 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1677622389
transform 1 0 2364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1677622389
transform 1 0 2388 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2604
timestamp 1677622389
transform 1 0 2388 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1677622389
transform 1 0 2412 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1677622389
transform 1 0 2500 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1677622389
transform 1 0 2492 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1677622389
transform 1 0 2412 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2872
timestamp 1677622389
transform 1 0 2492 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1677622389
transform 1 0 2452 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2630
timestamp 1677622389
transform 1 0 2428 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1677622389
transform 1 0 2476 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_2873
timestamp 1677622389
transform 1 0 2508 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2646
timestamp 1677622389
transform 1 0 2508 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_2874
timestamp 1677622389
transform 1 0 2644 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1677622389
transform 1 0 2556 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1677622389
transform 1 0 2564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1677622389
transform 1 0 2596 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1677622389
transform 1 0 2556 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1677622389
transform 1 0 2596 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1677622389
transform 1 0 2564 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2875
timestamp 1677622389
transform 1 0 2660 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2632
timestamp 1677622389
transform 1 0 2660 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1677622389
transform 1 0 2684 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1677622389
transform 1 0 2708 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2876
timestamp 1677622389
transform 1 0 2700 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1677622389
transform 1 0 2716 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1677622389
transform 1 0 2684 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1677622389
transform 1 0 2700 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2836
timestamp 1677622389
transform 1 0 2804 0 1 3345
box -2 -2 2 2
use M3_M2  M3_M2_2525
timestamp 1677622389
transform 1 0 2812 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1677622389
transform 1 0 2804 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2973
timestamp 1677622389
transform 1 0 2740 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1677622389
transform 1 0 2796 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2607
timestamp 1677622389
transform 1 0 2684 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3020
timestamp 1677622389
transform 1 0 2700 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2608
timestamp 1677622389
transform 1 0 2796 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1677622389
transform 1 0 2836 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2878
timestamp 1677622389
transform 1 0 2836 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1677622389
transform 1 0 2844 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2575
timestamp 1677622389
transform 1 0 2844 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1677622389
transform 1 0 2868 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1677622389
transform 1 0 2892 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2975
timestamp 1677622389
transform 1 0 2908 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1677622389
transform 1 0 2940 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2527
timestamp 1677622389
transform 1 0 2964 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2880
timestamp 1677622389
transform 1 0 2964 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1677622389
transform 1 0 2972 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2577
timestamp 1677622389
transform 1 0 2972 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3022
timestamp 1677622389
transform 1 0 2972 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1677622389
transform 1 0 2996 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1677622389
transform 1 0 3012 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1677622389
transform 1 0 3036 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1677622389
transform 1 0 3052 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2610
timestamp 1677622389
transform 1 0 3052 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2883
timestamp 1677622389
transform 1 0 3140 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1677622389
transform 1 0 3092 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2647
timestamp 1677622389
transform 1 0 3076 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1677622389
transform 1 0 3156 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2980
timestamp 1677622389
transform 1 0 3156 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2655
timestamp 1677622389
transform 1 0 3148 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1677622389
transform 1 0 3164 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_2884
timestamp 1677622389
transform 1 0 3180 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1677622389
transform 1 0 3212 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1677622389
transform 1 0 3236 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1677622389
transform 1 0 3252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1677622389
transform 1 0 3228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1677622389
transform 1 0 3244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2611
timestamp 1677622389
transform 1 0 3228 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2888
timestamp 1677622389
transform 1 0 3268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1677622389
transform 1 0 3260 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2612
timestamp 1677622389
transform 1 0 3260 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1677622389
transform 1 0 3260 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_2889
timestamp 1677622389
transform 1 0 3292 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1677622389
transform 1 0 3348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1677622389
transform 1 0 3332 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2657
timestamp 1677622389
transform 1 0 3324 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1677622389
transform 1 0 3348 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3025
timestamp 1677622389
transform 1 0 3340 0 1 3305
box -2 -2 2 2
use M3_M2  M3_M2_2658
timestamp 1677622389
transform 1 0 3364 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1677622389
transform 1 0 3388 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2985
timestamp 1677622389
transform 1 0 3380 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1677622389
transform 1 0 3396 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2633
timestamp 1677622389
transform 1 0 3396 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1677622389
transform 1 0 3412 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1677622389
transform 1 0 3436 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2890
timestamp 1677622389
transform 1 0 3412 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2553
timestamp 1677622389
transform 1 0 3436 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2986
timestamp 1677622389
transform 1 0 3420 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1677622389
transform 1 0 3420 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2987
timestamp 1677622389
transform 1 0 3460 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2486
timestamp 1677622389
transform 1 0 3492 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2891
timestamp 1677622389
transform 1 0 3476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1677622389
transform 1 0 3484 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2578
timestamp 1677622389
transform 1 0 3484 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2988
timestamp 1677622389
transform 1 0 3492 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1677622389
transform 1 0 3500 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1677622389
transform 1 0 3508 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1677622389
transform 1 0 3524 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2989
timestamp 1677622389
transform 1 0 3524 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2531
timestamp 1677622389
transform 1 0 3588 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2893
timestamp 1677622389
transform 1 0 3540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1677622389
transform 1 0 3588 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1677622389
transform 1 0 3628 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2503
timestamp 1677622389
transform 1 0 3660 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1677622389
transform 1 0 3668 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2894
timestamp 1677622389
transform 1 0 3652 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2555
timestamp 1677622389
transform 1 0 3660 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2895
timestamp 1677622389
transform 1 0 3668 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1677622389
transform 1 0 3692 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1677622389
transform 1 0 3660 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1677622389
transform 1 0 3684 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1677622389
transform 1 0 3692 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2634
timestamp 1677622389
transform 1 0 3668 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1677622389
transform 1 0 3732 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1677622389
transform 1 0 3740 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2897
timestamp 1677622389
transform 1 0 3732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1677622389
transform 1 0 3740 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1677622389
transform 1 0 3748 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1677622389
transform 1 0 3764 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1677622389
transform 1 0 3780 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1677622389
transform 1 0 3780 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2504
timestamp 1677622389
transform 1 0 3820 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1677622389
transform 1 0 3812 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1677622389
transform 1 0 3860 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1677622389
transform 1 0 3876 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1677622389
transform 1 0 3900 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1677622389
transform 1 0 3876 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2900
timestamp 1677622389
transform 1 0 3876 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1677622389
transform 1 0 3924 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1677622389
transform 1 0 3980 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2536
timestamp 1677622389
transform 1 0 4076 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2901
timestamp 1677622389
transform 1 0 4076 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1677622389
transform 1 0 3996 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1677622389
transform 1 0 4044 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2635
timestamp 1677622389
transform 1 0 4044 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1677622389
transform 1 0 4092 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1677622389
transform 1 0 4108 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2902
timestamp 1677622389
transform 1 0 4108 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1677622389
transform 1 0 4156 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2637
timestamp 1677622389
transform 1 0 4156 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_3003
timestamp 1677622389
transform 1 0 4212 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2638
timestamp 1677622389
transform 1 0 4204 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1677622389
transform 1 0 4284 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1677622389
transform 1 0 4348 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1677622389
transform 1 0 4276 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1677622389
transform 1 0 4316 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1677622389
transform 1 0 4332 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2903
timestamp 1677622389
transform 1 0 4356 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1677622389
transform 1 0 4276 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1677622389
transform 1 0 4332 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2659
timestamp 1677622389
transform 1 0 4292 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1677622389
transform 1 0 4348 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_2904
timestamp 1677622389
transform 1 0 4380 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2538
timestamp 1677622389
transform 1 0 4404 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1677622389
transform 1 0 4396 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2905
timestamp 1677622389
transform 1 0 4404 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1677622389
transform 1 0 4420 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2580
timestamp 1677622389
transform 1 0 4388 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3006
timestamp 1677622389
transform 1 0 4396 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2581
timestamp 1677622389
transform 1 0 4404 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3007
timestamp 1677622389
transform 1 0 4412 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2582
timestamp 1677622389
transform 1 0 4420 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1677622389
transform 1 0 4396 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3008
timestamp 1677622389
transform 1 0 4436 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2507
timestamp 1677622389
transform 1 0 4468 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1677622389
transform 1 0 4484 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2907
timestamp 1677622389
transform 1 0 4460 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2560
timestamp 1677622389
transform 1 0 4468 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3009
timestamp 1677622389
transform 1 0 4468 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1677622389
transform 1 0 4484 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2616
timestamp 1677622389
transform 1 0 4468 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1677622389
transform 1 0 4484 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2837
timestamp 1677622389
transform 1 0 4516 0 1 3345
box -2 -2 2 2
use M3_M2  M3_M2_2561
timestamp 1677622389
transform 1 0 4508 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3011
timestamp 1677622389
transform 1 0 4516 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2650
timestamp 1677622389
transform 1 0 4516 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1677622389
transform 1 0 4564 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1677622389
transform 1 0 4540 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2908
timestamp 1677622389
transform 1 0 4540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1677622389
transform 1 0 4556 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2562
timestamp 1677622389
transform 1 0 4564 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2910
timestamp 1677622389
transform 1 0 4572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1677622389
transform 1 0 4548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1677622389
transform 1 0 4564 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2618
timestamp 1677622389
transform 1 0 4540 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1677622389
transform 1 0 4532 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1677622389
transform 1 0 4572 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3014
timestamp 1677622389
transform 1 0 4580 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2652
timestamp 1677622389
transform 1 0 4556 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1677622389
transform 1 0 4580 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2911
timestamp 1677622389
transform 1 0 4620 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1677622389
transform 1 0 4636 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1677622389
transform 1 0 4620 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3015
timestamp 1677622389
transform 1 0 4628 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2661
timestamp 1677622389
transform 1 0 4636 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1677622389
transform 1 0 4652 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2913
timestamp 1677622389
transform 1 0 4660 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2492
timestamp 1677622389
transform 1 0 4676 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2914
timestamp 1677622389
transform 1 0 4676 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2563
timestamp 1677622389
transform 1 0 4700 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1677622389
transform 1 0 4700 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1677622389
transform 1 0 4756 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1677622389
transform 1 0 4764 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2662
timestamp 1677622389
transform 1 0 4684 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1677622389
transform 1 0 4764 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_2915
timestamp 1677622389
transform 1 0 4788 0 1 3335
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_28
timestamp 1677622389
transform 1 0 24 0 1 3270
box -10 -3 10 3
use FILL  FILL_2678
timestamp 1677622389
transform 1 0 72 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1677622389
transform 1 0 80 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_215
timestamp 1677622389
transform -1 0 192 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2692
timestamp 1677622389
transform 1 0 192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1677622389
transform 1 0 200 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1677622389
transform 1 0 208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1677622389
transform 1 0 216 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1677622389
transform 1 0 224 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_125
timestamp 1677622389
transform 1 0 232 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2697
timestamp 1677622389
transform 1 0 272 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1677622389
transform 1 0 280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1677622389
transform 1 0 288 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_123
timestamp 1677622389
transform -1 0 336 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2700
timestamp 1677622389
transform 1 0 336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1677622389
transform 1 0 344 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_216
timestamp 1677622389
transform 1 0 352 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_124
timestamp 1677622389
transform -1 0 408 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2702
timestamp 1677622389
transform 1 0 408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1677622389
transform 1 0 416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1677622389
transform 1 0 424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1677622389
transform 1 0 432 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_125
timestamp 1677622389
transform 1 0 440 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2719
timestamp 1677622389
transform 1 0 480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1677622389
transform 1 0 488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1677622389
transform 1 0 496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1677622389
transform 1 0 504 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_126
timestamp 1677622389
transform 1 0 512 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2723
timestamp 1677622389
transform 1 0 552 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1677622389
transform 1 0 560 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1677622389
transform 1 0 568 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1677622389
transform 1 0 576 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2726
timestamp 1677622389
transform 1 0 672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1677622389
transform 1 0 680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1677622389
transform 1 0 688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1677622389
transform 1 0 696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1677622389
transform 1 0 704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1677622389
transform 1 0 712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1677622389
transform 1 0 720 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1677622389
transform 1 0 728 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1677622389
transform 1 0 736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1677622389
transform 1 0 744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1677622389
transform 1 0 752 0 -1 3370
box -8 -3 16 105
use BUFX2  BUFX2_22
timestamp 1677622389
transform -1 0 784 0 -1 3370
box -5 -3 28 105
use FILL  FILL_2746
timestamp 1677622389
transform 1 0 784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1677622389
transform 1 0 792 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1677622389
transform 1 0 800 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1677622389
transform 1 0 808 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2764
timestamp 1677622389
transform 1 0 904 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_218
timestamp 1677622389
transform 1 0 912 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2768
timestamp 1677622389
transform 1 0 928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1677622389
transform 1 0 936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1677622389
transform 1 0 944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1677622389
transform 1 0 952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1677622389
transform 1 0 960 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1677622389
transform 1 0 968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1677622389
transform 1 0 976 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1677622389
transform 1 0 984 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1677622389
transform 1 0 992 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1677622389
transform 1 0 1000 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1677622389
transform 1 0 1008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1677622389
transform 1 0 1016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1677622389
transform 1 0 1024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1677622389
transform 1 0 1032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1677622389
transform 1 0 1040 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1677622389
transform 1 0 1048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1677622389
transform 1 0 1056 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1677622389
transform 1 0 1064 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_127
timestamp 1677622389
transform 1 0 1072 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2806
timestamp 1677622389
transform 1 0 1112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1677622389
transform 1 0 1120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1677622389
transform 1 0 1128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1677622389
transform 1 0 1136 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1677622389
transform 1 0 1144 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1677622389
transform 1 0 1152 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1677622389
transform 1 0 1160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1677622389
transform 1 0 1168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1677622389
transform 1 0 1176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1677622389
transform 1 0 1184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1677622389
transform 1 0 1192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1677622389
transform 1 0 1200 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_219
timestamp 1677622389
transform 1 0 1208 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2823
timestamp 1677622389
transform 1 0 1224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1677622389
transform 1 0 1232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1677622389
transform 1 0 1240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1677622389
transform 1 0 1248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1677622389
transform 1 0 1256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1677622389
transform 1 0 1264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1677622389
transform 1 0 1272 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1677622389
transform 1 0 1280 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2834
timestamp 1677622389
transform 1 0 1312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1677622389
transform 1 0 1320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1677622389
transform 1 0 1328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1677622389
transform 1 0 1336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1677622389
transform 1 0 1344 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1677622389
transform 1 0 1352 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2851
timestamp 1677622389
transform 1 0 1448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1677622389
transform 1 0 1456 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_220
timestamp 1677622389
transform 1 0 1464 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2857
timestamp 1677622389
transform 1 0 1480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1677622389
transform 1 0 1488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1677622389
transform 1 0 1496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1677622389
transform 1 0 1504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1677622389
transform 1 0 1512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1677622389
transform 1 0 1520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1677622389
transform 1 0 1528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1677622389
transform 1 0 1536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1677622389
transform 1 0 1544 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1677622389
transform 1 0 1552 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1677622389
transform 1 0 1560 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1677622389
transform 1 0 1568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1677622389
transform 1 0 1576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1677622389
transform 1 0 1584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1677622389
transform 1 0 1592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1677622389
transform 1 0 1600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1677622389
transform 1 0 1608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1677622389
transform 1 0 1616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1677622389
transform 1 0 1624 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1677622389
transform 1 0 1632 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1677622389
transform 1 0 1640 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1677622389
transform 1 0 1648 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_222
timestamp 1677622389
transform -1 0 1672 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2886
timestamp 1677622389
transform 1 0 1672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1677622389
transform 1 0 1680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1677622389
transform 1 0 1688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1677622389
transform 1 0 1696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1677622389
transform 1 0 1704 0 -1 3370
box -8 -3 16 105
use BUFX2  BUFX2_23
timestamp 1677622389
transform -1 0 1736 0 -1 3370
box -5 -3 28 105
use FILL  FILL_2891
timestamp 1677622389
transform 1 0 1736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1677622389
transform 1 0 1744 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2664
timestamp 1677622389
transform 1 0 1764 0 1 3275
box -3 -3 3 3
use BUFX2  BUFX2_24
timestamp 1677622389
transform 1 0 1752 0 -1 3370
box -5 -3 28 105
use FILL  FILL_2897
timestamp 1677622389
transform 1 0 1776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1677622389
transform 1 0 1784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1677622389
transform 1 0 1792 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_224
timestamp 1677622389
transform 1 0 1800 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2912
timestamp 1677622389
transform 1 0 1816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1677622389
transform 1 0 1824 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_196
timestamp 1677622389
transform -1 0 1928 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2914
timestamp 1677622389
transform 1 0 1928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1677622389
transform 1 0 1936 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_197
timestamp 1677622389
transform 1 0 1944 0 -1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2665
timestamp 1677622389
transform 1 0 2092 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_198
timestamp 1677622389
transform 1 0 2040 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_199
timestamp 1677622389
transform 1 0 2136 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_225
timestamp 1677622389
transform 1 0 2232 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2946
timestamp 1677622389
transform 1 0 2248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1677622389
transform 1 0 2256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1677622389
transform 1 0 2264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1677622389
transform 1 0 2272 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1677622389
transform 1 0 2280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1677622389
transform 1 0 2288 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1677622389
transform 1 0 2296 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_130
timestamp 1677622389
transform 1 0 2304 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2965
timestamp 1677622389
transform 1 0 2344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1677622389
transform 1 0 2352 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_228
timestamp 1677622389
transform 1 0 2360 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2967
timestamp 1677622389
transform 1 0 2376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1677622389
transform 1 0 2384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1677622389
transform 1 0 2392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1677622389
transform 1 0 2400 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1677622389
transform -1 0 2504 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2971
timestamp 1677622389
transform 1 0 2504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1677622389
transform 1 0 2512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1677622389
transform 1 0 2520 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_229
timestamp 1677622389
transform 1 0 2528 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2977
timestamp 1677622389
transform 1 0 2544 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1677622389
transform 1 0 2552 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_203
timestamp 1677622389
transform -1 0 2656 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2979
timestamp 1677622389
transform 1 0 2656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1677622389
transform 1 0 2664 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1677622389
transform 1 0 2672 0 -1 3370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1677622389
transform 1 0 2704 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2990
timestamp 1677622389
transform 1 0 2800 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1677622389
transform 1 0 2808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1677622389
transform 1 0 2816 0 -1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_33
timestamp 1677622389
transform 1 0 2824 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2993
timestamp 1677622389
transform 1 0 2848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1677622389
transform 1 0 2856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1677622389
transform 1 0 2864 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1677622389
transform 1 0 2872 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1677622389
transform 1 0 2880 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1677622389
transform 1 0 2888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1677622389
transform 1 0 2896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1677622389
transform 1 0 2904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1677622389
transform 1 0 2912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1677622389
transform 1 0 2920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1677622389
transform 1 0 2928 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_67
timestamp 1677622389
transform -1 0 2968 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3015
timestamp 1677622389
transform 1 0 2968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1677622389
transform 1 0 2976 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1677622389
transform 1 0 2984 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_68
timestamp 1677622389
transform -1 0 3024 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3018
timestamp 1677622389
transform 1 0 3024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1677622389
transform 1 0 3032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1677622389
transform 1 0 3040 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1677622389
transform 1 0 3048 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2666
timestamp 1677622389
transform 1 0 3108 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_208
timestamp 1677622389
transform -1 0 3152 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3022
timestamp 1677622389
transform 1 0 3152 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_231
timestamp 1677622389
transform -1 0 3176 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3023
timestamp 1677622389
transform 1 0 3176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1677622389
transform 1 0 3184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1677622389
transform 1 0 3192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1677622389
transform 1 0 3200 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1677622389
transform 1 0 3208 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_129
timestamp 1677622389
transform -1 0 3256 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3030
timestamp 1677622389
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1677622389
transform 1 0 3264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1677622389
transform 1 0 3272 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_232
timestamp 1677622389
transform -1 0 3296 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3033
timestamp 1677622389
transform 1 0 3296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1677622389
transform 1 0 3304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1677622389
transform 1 0 3312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1677622389
transform 1 0 3320 0 -1 3370
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1677622389
transform -1 0 3360 0 -1 3370
box -8 -3 40 105
use FILL  FILL_3041
timestamp 1677622389
transform 1 0 3360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1677622389
transform 1 0 3368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1677622389
transform 1 0 3376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1677622389
transform 1 0 3384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1677622389
transform 1 0 3392 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_132
timestamp 1677622389
transform 1 0 3400 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3046
timestamp 1677622389
transform 1 0 3440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1677622389
transform 1 0 3448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1677622389
transform 1 0 3456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1677622389
transform 1 0 3464 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1677622389
transform 1 0 3472 0 -1 3370
box -8 -3 16 105
use AND2X2  AND2X2_10
timestamp 1677622389
transform 1 0 3480 0 -1 3370
box -8 -3 40 105
use FILL  FILL_3056
timestamp 1677622389
transform 1 0 3512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1677622389
transform 1 0 3520 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2667
timestamp 1677622389
transform 1 0 3572 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_211
timestamp 1677622389
transform 1 0 3528 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3070
timestamp 1677622389
transform 1 0 3624 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1677622389
transform 1 0 3632 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1677622389
transform 1 0 3640 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_130
timestamp 1677622389
transform -1 0 3688 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3081
timestamp 1677622389
transform 1 0 3688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1677622389
transform 1 0 3696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1677622389
transform 1 0 3704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1677622389
transform 1 0 3712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1677622389
transform 1 0 3720 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_133
timestamp 1677622389
transform -1 0 3768 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3096
timestamp 1677622389
transform 1 0 3768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1677622389
transform 1 0 3776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1677622389
transform 1 0 3784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1677622389
transform 1 0 3792 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1677622389
transform 1 0 3800 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1677622389
transform 1 0 3808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1677622389
transform 1 0 3816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1677622389
transform 1 0 3824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1677622389
transform 1 0 3832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1677622389
transform 1 0 3840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1677622389
transform 1 0 3848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1677622389
transform 1 0 3856 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_213
timestamp 1677622389
transform 1 0 3864 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3123
timestamp 1677622389
transform 1 0 3960 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_237
timestamp 1677622389
transform 1 0 3968 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3124
timestamp 1677622389
transform 1 0 3984 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1677622389
transform -1 0 4088 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3125
timestamp 1677622389
transform 1 0 4088 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_215
timestamp 1677622389
transform 1 0 4096 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3136
timestamp 1677622389
transform 1 0 4192 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_238
timestamp 1677622389
transform 1 0 4200 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3137
timestamp 1677622389
transform 1 0 4216 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1677622389
transform 1 0 4224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1677622389
transform 1 0 4232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1677622389
transform 1 0 4240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1677622389
transform 1 0 4248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1677622389
transform 1 0 4256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1677622389
transform 1 0 4264 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1677622389
transform -1 0 4368 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3156
timestamp 1677622389
transform 1 0 4368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1677622389
transform 1 0 4376 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_133
timestamp 1677622389
transform 1 0 4384 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3165
timestamp 1677622389
transform 1 0 4424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1677622389
transform 1 0 4432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1677622389
transform 1 0 4440 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_136
timestamp 1677622389
transform -1 0 4488 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3168
timestamp 1677622389
transform 1 0 4488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1677622389
transform 1 0 4496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1677622389
transform 1 0 4504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1677622389
transform 1 0 4512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1677622389
transform 1 0 4520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1677622389
transform 1 0 4528 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_134
timestamp 1677622389
transform 1 0 4536 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3189
timestamp 1677622389
transform 1 0 4576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1677622389
transform 1 0 4584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1677622389
transform 1 0 4592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1677622389
transform 1 0 4600 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2668
timestamp 1677622389
transform 1 0 4628 0 1 3275
box -3 -3 3 3
use AOI22X1  AOI22X1_137
timestamp 1677622389
transform 1 0 4608 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3193
timestamp 1677622389
transform 1 0 4648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1677622389
transform 1 0 4656 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_218
timestamp 1677622389
transform 1 0 4664 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_243
timestamp 1677622389
transform -1 0 4776 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3195
timestamp 1677622389
transform 1 0 4776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1677622389
transform 1 0 4784 0 -1 3370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_29
timestamp 1677622389
transform 1 0 4843 0 1 3270
box -10 -3 10 3
use M3_M2  M3_M2_2752
timestamp 1677622389
transform 1 0 100 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1677622389
transform 1 0 116 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3049
timestamp 1677622389
transform 1 0 116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1677622389
transform 1 0 116 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2810
timestamp 1677622389
transform 1 0 116 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1677622389
transform 1 0 164 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3050
timestamp 1677622389
transform 1 0 164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1677622389
transform 1 0 140 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2838
timestamp 1677622389
transform 1 0 140 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3051
timestamp 1677622389
transform 1 0 236 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2811
timestamp 1677622389
transform 1 0 228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1677622389
transform 1 0 260 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1677622389
transform 1 0 268 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1677622389
transform 1 0 324 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1677622389
transform 1 0 348 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1677622389
transform 1 0 316 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1677622389
transform 1 0 268 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1677622389
transform 1 0 356 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3052
timestamp 1677622389
transform 1 0 316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1677622389
transform 1 0 348 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1677622389
transform 1 0 356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1677622389
transform 1 0 268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1677622389
transform 1 0 372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1677622389
transform 1 0 396 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2702
timestamp 1677622389
transform 1 0 412 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3057
timestamp 1677622389
transform 1 0 420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1677622389
transform 1 0 404 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1677622389
transform 1 0 412 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1677622389
transform 1 0 428 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2689
timestamp 1677622389
transform 1 0 444 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3058
timestamp 1677622389
transform 1 0 444 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1677622389
transform 1 0 468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2728
timestamp 1677622389
transform 1 0 564 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3059
timestamp 1677622389
transform 1 0 508 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2754
timestamp 1677622389
transform 1 0 532 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3060
timestamp 1677622389
transform 1 0 564 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1677622389
transform 1 0 484 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2812
timestamp 1677622389
transform 1 0 524 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1677622389
transform 1 0 484 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1677622389
transform 1 0 572 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3162
timestamp 1677622389
transform 1 0 572 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2813
timestamp 1677622389
transform 1 0 572 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1677622389
transform 1 0 612 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1677622389
transform 1 0 644 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3061
timestamp 1677622389
transform 1 0 604 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1677622389
transform 1 0 620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1677622389
transform 1 0 636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1677622389
transform 1 0 612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1677622389
transform 1 0 628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1677622389
transform 1 0 644 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2814
timestamp 1677622389
transform 1 0 628 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1677622389
transform 1 0 692 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3166
timestamp 1677622389
transform 1 0 692 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2690
timestamp 1677622389
transform 1 0 732 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3064
timestamp 1677622389
transform 1 0 724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1677622389
transform 1 0 732 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2731
timestamp 1677622389
transform 1 0 772 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3066
timestamp 1677622389
transform 1 0 772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1677622389
transform 1 0 764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1677622389
transform 1 0 780 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1677622389
transform 1 0 788 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2840
timestamp 1677622389
transform 1 0 764 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3067
timestamp 1677622389
transform 1 0 804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1677622389
transform 1 0 812 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2841
timestamp 1677622389
transform 1 0 812 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1677622389
transform 1 0 828 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1677622389
transform 1 0 860 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3258
timestamp 1677622389
transform 1 0 860 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2732
timestamp 1677622389
transform 1 0 900 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3068
timestamp 1677622389
transform 1 0 892 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2756
timestamp 1677622389
transform 1 0 908 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3069
timestamp 1677622389
transform 1 0 916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1677622389
transform 1 0 884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1677622389
transform 1 0 900 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2779
timestamp 1677622389
transform 1 0 916 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3259
timestamp 1677622389
transform 1 0 924 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2757
timestamp 1677622389
transform 1 0 1020 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3173
timestamp 1677622389
transform 1 0 1012 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1677622389
transform 1 0 996 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2816
timestamp 1677622389
transform 1 0 1004 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3261
timestamp 1677622389
transform 1 0 1020 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1677622389
transform 1 0 1036 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2758
timestamp 1677622389
transform 1 0 1044 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3071
timestamp 1677622389
transform 1 0 1060 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2733
timestamp 1677622389
transform 1 0 1068 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3072
timestamp 1677622389
transform 1 0 1068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1677622389
transform 1 0 1076 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2817
timestamp 1677622389
transform 1 0 1068 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1677622389
transform 1 0 1076 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1677622389
transform 1 0 1116 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3073
timestamp 1677622389
transform 1 0 1092 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2759
timestamp 1677622389
transform 1 0 1108 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3175
timestamp 1677622389
transform 1 0 1108 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2818
timestamp 1677622389
transform 1 0 1092 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3176
timestamp 1677622389
transform 1 0 1116 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1677622389
transform 1 0 1132 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2760
timestamp 1677622389
transform 1 0 1132 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1677622389
transform 1 0 1172 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1677622389
transform 1 0 1148 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3074
timestamp 1677622389
transform 1 0 1140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1677622389
transform 1 0 1156 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1677622389
transform 1 0 1132 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2761
timestamp 1677622389
transform 1 0 1180 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3076
timestamp 1677622389
transform 1 0 1188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1677622389
transform 1 0 1148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1677622389
transform 1 0 1172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1677622389
transform 1 0 1180 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2819
timestamp 1677622389
transform 1 0 1156 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1677622389
transform 1 0 1172 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1677622389
transform 1 0 1172 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1677622389
transform 1 0 1188 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1677622389
transform 1 0 1236 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1677622389
transform 1 0 1252 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1677622389
transform 1 0 1276 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3033
timestamp 1677622389
transform 1 0 1324 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2822
timestamp 1677622389
transform 1 0 1340 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3077
timestamp 1677622389
transform 1 0 1372 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2823
timestamp 1677622389
transform 1 0 1364 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3034
timestamp 1677622389
transform 1 0 1396 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1677622389
transform 1 0 1428 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1677622389
transform 1 0 1444 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2762
timestamp 1677622389
transform 1 0 1444 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3181
timestamp 1677622389
transform 1 0 1444 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1677622389
transform 1 0 1460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1677622389
transform 1 0 1476 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2763
timestamp 1677622389
transform 1 0 1484 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3080
timestamp 1677622389
transform 1 0 1492 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2781
timestamp 1677622389
transform 1 0 1460 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3182
timestamp 1677622389
transform 1 0 1468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2782
timestamp 1677622389
transform 1 0 1492 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3081
timestamp 1677622389
transform 1 0 1540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1677622389
transform 1 0 1524 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2783
timestamp 1677622389
transform 1 0 1532 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1677622389
transform 1 0 1524 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3184
timestamp 1677622389
transform 1 0 1556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1677622389
transform 1 0 1588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1677622389
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2784
timestamp 1677622389
transform 1 0 1588 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3186
timestamp 1677622389
transform 1 0 1596 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2825
timestamp 1677622389
transform 1 0 1596 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3083
timestamp 1677622389
transform 1 0 1684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1677622389
transform 1 0 1700 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1677622389
transform 1 0 1676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1677622389
transform 1 0 1692 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2706
timestamp 1677622389
transform 1 0 1724 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3085
timestamp 1677622389
transform 1 0 1724 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2707
timestamp 1677622389
transform 1 0 1756 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3189
timestamp 1677622389
transform 1 0 1748 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2826
timestamp 1677622389
transform 1 0 1748 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1677622389
transform 1 0 1748 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1677622389
transform 1 0 1772 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3190
timestamp 1677622389
transform 1 0 1772 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2845
timestamp 1677622389
transform 1 0 1764 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1677622389
transform 1 0 1788 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3086
timestamp 1677622389
transform 1 0 1804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1677622389
transform 1 0 1844 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1677622389
transform 1 0 1860 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1677622389
transform 1 0 1836 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1677622389
transform 1 0 1852 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1677622389
transform 1 0 1908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1677622389
transform 1 0 1948 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1677622389
transform 1 0 1956 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2785
timestamp 1677622389
transform 1 0 1972 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3089
timestamp 1677622389
transform 1 0 1988 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2682
timestamp 1677622389
transform 1 0 2028 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1677622389
transform 1 0 2028 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3196
timestamp 1677622389
transform 1 0 2028 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1677622389
transform 1 0 2044 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2846
timestamp 1677622389
transform 1 0 2044 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1677622389
transform 1 0 2076 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1677622389
transform 1 0 2068 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1677622389
transform 1 0 2084 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1677622389
transform 1 0 2092 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3090
timestamp 1677622389
transform 1 0 2068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1677622389
transform 1 0 2076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1677622389
transform 1 0 2092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1677622389
transform 1 0 2108 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1677622389
transform 1 0 2100 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2786
timestamp 1677622389
transform 1 0 2108 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1677622389
transform 1 0 2132 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1677622389
transform 1 0 2124 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3094
timestamp 1677622389
transform 1 0 2140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1677622389
transform 1 0 2124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1677622389
transform 1 0 2164 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1677622389
transform 1 0 2188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1677622389
transform 1 0 2196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1677622389
transform 1 0 2212 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1677622389
transform 1 0 2228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1677622389
transform 1 0 2196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1677622389
transform 1 0 2220 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2847
timestamp 1677622389
transform 1 0 2196 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1677622389
transform 1 0 2228 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1677622389
transform 1 0 2276 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3203
timestamp 1677622389
transform 1 0 2276 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1677622389
transform 1 0 2292 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2848
timestamp 1677622389
transform 1 0 2292 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3026
timestamp 1677622389
transform 1 0 2308 0 1 3245
box -2 -2 2 2
use M3_M2  M3_M2_2710
timestamp 1677622389
transform 1 0 2308 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1677622389
transform 1 0 2316 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1677622389
transform 1 0 2348 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3099
timestamp 1677622389
transform 1 0 2308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1677622389
transform 1 0 2316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1677622389
transform 1 0 2324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1677622389
transform 1 0 2340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1677622389
transform 1 0 2356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1677622389
transform 1 0 2332 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2788
timestamp 1677622389
transform 1 0 2356 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3206
timestamp 1677622389
transform 1 0 2364 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2849
timestamp 1677622389
transform 1 0 2324 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1677622389
transform 1 0 2348 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1677622389
transform 1 0 2380 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1677622389
transform 1 0 2388 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3104
timestamp 1677622389
transform 1 0 2404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1677622389
transform 1 0 2420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1677622389
transform 1 0 2428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1677622389
transform 1 0 2412 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2790
timestamp 1677622389
transform 1 0 2420 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3208
timestamp 1677622389
transform 1 0 2428 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2852
timestamp 1677622389
transform 1 0 2420 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1677622389
transform 1 0 2452 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3107
timestamp 1677622389
transform 1 0 2476 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1677622389
transform 1 0 2468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2853
timestamp 1677622389
transform 1 0 2500 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3108
timestamp 1677622389
transform 1 0 2516 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2764
timestamp 1677622389
transform 1 0 2524 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3210
timestamp 1677622389
transform 1 0 2524 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2739
timestamp 1677622389
transform 1 0 2540 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1677622389
transform 1 0 2564 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1677622389
transform 1 0 2628 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3109
timestamp 1677622389
transform 1 0 2572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1677622389
transform 1 0 2620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1677622389
transform 1 0 2628 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1677622389
transform 1 0 2540 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1677622389
transform 1 0 2628 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2854
timestamp 1677622389
transform 1 0 2540 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1677622389
transform 1 0 2604 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1677622389
transform 1 0 2620 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3112
timestamp 1677622389
transform 1 0 2676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1677622389
transform 1 0 2700 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1677622389
transform 1 0 2684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1677622389
transform 1 0 2692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1677622389
transform 1 0 2740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1677622389
transform 1 0 2740 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2857
timestamp 1677622389
transform 1 0 2740 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3115
timestamp 1677622389
transform 1 0 2804 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2791
timestamp 1677622389
transform 1 0 2804 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1677622389
transform 1 0 2836 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1677622389
transform 1 0 2836 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1677622389
transform 1 0 2852 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3216
timestamp 1677622389
transform 1 0 2844 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1677622389
transform 1 0 2860 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2766
timestamp 1677622389
transform 1 0 2860 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3038
timestamp 1677622389
transform 1 0 2892 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1677622389
transform 1 0 2876 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1677622389
transform 1 0 2860 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1677622389
transform 1 0 2868 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2741
timestamp 1677622389
transform 1 0 2916 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1677622389
transform 1 0 2932 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3039
timestamp 1677622389
transform 1 0 2940 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1677622389
transform 1 0 2924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1677622389
transform 1 0 2908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1677622389
transform 1 0 2916 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1677622389
transform 1 0 2908 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1677622389
transform 1 0 2932 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3221
timestamp 1677622389
transform 1 0 2932 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2768
timestamp 1677622389
transform 1 0 2948 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3040
timestamp 1677622389
transform 1 0 2972 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1677622389
transform 1 0 2988 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2793
timestamp 1677622389
transform 1 0 2988 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1677622389
transform 1 0 3020 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3222
timestamp 1677622389
transform 1 0 3036 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1677622389
transform 1 0 3068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1677622389
transform 1 0 3084 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1677622389
transform 1 0 3116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1677622389
transform 1 0 3076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1677622389
transform 1 0 3092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1677622389
transform 1 0 3108 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2858
timestamp 1677622389
transform 1 0 3076 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1677622389
transform 1 0 3116 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3226
timestamp 1677622389
transform 1 0 3124 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2859
timestamp 1677622389
transform 1 0 3124 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1677622389
transform 1 0 3180 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3122
timestamp 1677622389
transform 1 0 3164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1677622389
transform 1 0 3180 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2796
timestamp 1677622389
transform 1 0 3164 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3227
timestamp 1677622389
transform 1 0 3172 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2797
timestamp 1677622389
transform 1 0 3180 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1677622389
transform 1 0 3196 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3124
timestamp 1677622389
transform 1 0 3196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1677622389
transform 1 0 3188 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2860
timestamp 1677622389
transform 1 0 3188 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1677622389
transform 1 0 3204 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1677622389
transform 1 0 3244 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1677622389
transform 1 0 3300 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1677622389
transform 1 0 3236 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3125
timestamp 1677622389
transform 1 0 3252 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2799
timestamp 1677622389
transform 1 0 3252 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1677622389
transform 1 0 3268 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3229
timestamp 1677622389
transform 1 0 3300 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2827
timestamp 1677622389
transform 1 0 3220 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1677622389
transform 1 0 3212 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1677622389
transform 1 0 3228 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1677622389
transform 1 0 3356 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3027
timestamp 1677622389
transform 1 0 3348 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1677622389
transform 1 0 3340 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1677622389
transform 1 0 3356 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2769
timestamp 1677622389
transform 1 0 3340 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3126
timestamp 1677622389
transform 1 0 3356 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2770
timestamp 1677622389
transform 1 0 3364 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1677622389
transform 1 0 3420 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3028
timestamp 1677622389
transform 1 0 3420 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1677622389
transform 1 0 3412 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1677622389
transform 1 0 3436 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1677622389
transform 1 0 3452 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2771
timestamp 1677622389
transform 1 0 3452 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1677622389
transform 1 0 3468 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3029
timestamp 1677622389
transform 1 0 3468 0 1 3235
box -2 -2 2 2
use M3_M2  M3_M2_2685
timestamp 1677622389
transform 1 0 3492 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3030
timestamp 1677622389
transform 1 0 3492 0 1 3235
box -2 -2 2 2
use M3_M2  M3_M2_2716
timestamp 1677622389
transform 1 0 3500 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3046
timestamp 1677622389
transform 1 0 3500 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1677622389
transform 1 0 3492 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2694
timestamp 1677622389
transform 1 0 3540 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3047
timestamp 1677622389
transform 1 0 3540 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1677622389
transform 1 0 3564 0 1 3235
box -2 -2 2 2
use M3_M2  M3_M2_2742
timestamp 1677622389
transform 1 0 3564 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3128
timestamp 1677622389
transform 1 0 3572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1677622389
transform 1 0 3604 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2743
timestamp 1677622389
transform 1 0 3612 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1677622389
transform 1 0 3612 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3230
timestamp 1677622389
transform 1 0 3612 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2773
timestamp 1677622389
transform 1 0 3628 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1677622389
transform 1 0 3628 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1677622389
transform 1 0 3628 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1677622389
transform 1 0 3652 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1677622389
transform 1 0 3676 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3129
timestamp 1677622389
transform 1 0 3652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1677622389
transform 1 0 3668 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2828
timestamp 1677622389
transform 1 0 3644 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1677622389
transform 1 0 3692 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3231
timestamp 1677622389
transform 1 0 3660 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1677622389
transform 1 0 3676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1677622389
transform 1 0 3684 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2717
timestamp 1677622389
transform 1 0 3740 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3131
timestamp 1677622389
transform 1 0 3716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1677622389
transform 1 0 3724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1677622389
transform 1 0 3740 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2802
timestamp 1677622389
transform 1 0 3724 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1677622389
transform 1 0 3724 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3234
timestamp 1677622389
transform 1 0 3764 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1677622389
transform 1 0 3772 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3134
timestamp 1677622389
transform 1 0 3772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1677622389
transform 1 0 3772 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2830
timestamp 1677622389
transform 1 0 3764 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3135
timestamp 1677622389
transform 1 0 3788 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2803
timestamp 1677622389
transform 1 0 3788 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1677622389
transform 1 0 3828 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1677622389
transform 1 0 3828 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1677622389
transform 1 0 3812 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3136
timestamp 1677622389
transform 1 0 3812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1677622389
transform 1 0 3828 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2745
timestamp 1677622389
transform 1 0 3844 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3236
timestamp 1677622389
transform 1 0 3844 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1677622389
transform 1 0 3860 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2804
timestamp 1677622389
transform 1 0 3868 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1677622389
transform 1 0 3884 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3237
timestamp 1677622389
transform 1 0 3876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1677622389
transform 1 0 3892 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2864
timestamp 1677622389
transform 1 0 3892 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3139
timestamp 1677622389
transform 1 0 3924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1677622389
transform 1 0 3940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1677622389
transform 1 0 3916 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2805
timestamp 1677622389
transform 1 0 3924 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3240
timestamp 1677622389
transform 1 0 3932 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2831
timestamp 1677622389
transform 1 0 3940 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1677622389
transform 1 0 3956 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3141
timestamp 1677622389
transform 1 0 3956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1677622389
transform 1 0 3988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1677622389
transform 1 0 3996 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2832
timestamp 1677622389
transform 1 0 3980 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1677622389
transform 1 0 3988 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1677622389
transform 1 0 4044 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1677622389
transform 1 0 4060 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3243
timestamp 1677622389
transform 1 0 4084 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2806
timestamp 1677622389
transform 1 0 4100 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1677622389
transform 1 0 4172 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3142
timestamp 1677622389
transform 1 0 4276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1677622389
transform 1 0 4228 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2833
timestamp 1677622389
transform 1 0 4276 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3245
timestamp 1677622389
transform 1 0 4332 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2697
timestamp 1677622389
transform 1 0 4364 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1677622389
transform 1 0 4380 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1677622389
transform 1 0 4380 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1677622389
transform 1 0 4372 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1677622389
transform 1 0 4396 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3143
timestamp 1677622389
transform 1 0 4372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1677622389
transform 1 0 4380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1677622389
transform 1 0 4396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1677622389
transform 1 0 4364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1677622389
transform 1 0 4388 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2807
timestamp 1677622389
transform 1 0 4396 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1677622389
transform 1 0 4388 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1677622389
transform 1 0 4436 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3146
timestamp 1677622389
transform 1 0 4436 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1677622389
transform 1 0 4428 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2835
timestamp 1677622389
transform 1 0 4428 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1677622389
transform 1 0 4468 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3249
timestamp 1677622389
transform 1 0 4460 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2721
timestamp 1677622389
transform 1 0 4484 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1677622389
transform 1 0 4508 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3147
timestamp 1677622389
transform 1 0 4484 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2777
timestamp 1677622389
transform 1 0 4500 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3148
timestamp 1677622389
transform 1 0 4508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1677622389
transform 1 0 4484 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1677622389
transform 1 0 4500 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2808
timestamp 1677622389
transform 1 0 4508 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3252
timestamp 1677622389
transform 1 0 4516 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2836
timestamp 1677622389
transform 1 0 4516 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1677622389
transform 1 0 4636 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1677622389
transform 1 0 4668 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1677622389
transform 1 0 4676 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1677622389
transform 1 0 4660 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3149
timestamp 1677622389
transform 1 0 4596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1677622389
transform 1 0 4660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1677622389
transform 1 0 4668 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1677622389
transform 1 0 4684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1677622389
transform 1 0 4572 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2809
timestamp 1677622389
transform 1 0 4596 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1677622389
transform 1 0 4708 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1677622389
transform 1 0 4700 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3153
timestamp 1677622389
transform 1 0 4708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1677622389
transform 1 0 4660 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1677622389
transform 1 0 4676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1677622389
transform 1 0 4692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1677622389
transform 1 0 4700 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2868
timestamp 1677622389
transform 1 0 4572 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1677622389
transform 1 0 4692 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1677622389
transform 1 0 4708 0 1 3185
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_30
timestamp 1677622389
transform 1 0 48 0 1 3170
box -10 -3 10 3
use FILL  FILL_3198
timestamp 1677622389
transform 1 0 72 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_244
timestamp 1677622389
transform -1 0 96 0 1 3170
box -9 -3 26 105
use FILL  FILL_3199
timestamp 1677622389
transform 1 0 96 0 1 3170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1677622389
transform 1 0 104 0 1 3170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1677622389
transform 1 0 112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1677622389
transform 1 0 120 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_219
timestamp 1677622389
transform 1 0 128 0 1 3170
box -8 -3 104 105
use FILL  FILL_3203
timestamp 1677622389
transform 1 0 224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1677622389
transform 1 0 232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1677622389
transform 1 0 240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1677622389
transform 1 0 248 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1677622389
transform 1 0 256 0 1 3170
box -8 -3 104 105
use FILL  FILL_3213
timestamp 1677622389
transform 1 0 352 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_245
timestamp 1677622389
transform -1 0 376 0 1 3170
box -9 -3 26 105
use FILL  FILL_3214
timestamp 1677622389
transform 1 0 376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1677622389
transform 1 0 384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1677622389
transform 1 0 392 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_139
timestamp 1677622389
transform -1 0 440 0 1 3170
box -8 -3 46 105
use FILL  FILL_3217
timestamp 1677622389
transform 1 0 440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1677622389
transform 1 0 448 0 1 3170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1677622389
transform 1 0 456 0 1 3170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1677622389
transform 1 0 464 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1677622389
transform 1 0 472 0 1 3170
box -8 -3 104 105
use FILL  FILL_3236
timestamp 1677622389
transform 1 0 568 0 1 3170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1677622389
transform 1 0 576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1677622389
transform 1 0 584 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_247
timestamp 1677622389
transform 1 0 592 0 1 3170
box -9 -3 26 105
use OAI22X1  OAI22X1_135
timestamp 1677622389
transform 1 0 608 0 1 3170
box -8 -3 46 105
use FILL  FILL_3247
timestamp 1677622389
transform 1 0 648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1677622389
transform 1 0 656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1677622389
transform 1 0 664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1677622389
transform 1 0 672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1677622389
transform 1 0 680 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_248
timestamp 1677622389
transform 1 0 688 0 1 3170
box -9 -3 26 105
use FILL  FILL_3252
timestamp 1677622389
transform 1 0 704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1677622389
transform 1 0 712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1677622389
transform 1 0 720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1677622389
transform 1 0 728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1677622389
transform 1 0 736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1677622389
transform 1 0 744 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2870
timestamp 1677622389
transform 1 0 796 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_141
timestamp 1677622389
transform 1 0 752 0 1 3170
box -8 -3 46 105
use FILL  FILL_3258
timestamp 1677622389
transform 1 0 792 0 1 3170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1677622389
transform 1 0 800 0 1 3170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1677622389
transform 1 0 808 0 1 3170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1677622389
transform 1 0 816 0 1 3170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1677622389
transform 1 0 824 0 1 3170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1677622389
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1677622389
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1677622389
transform 1 0 848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1677622389
transform 1 0 856 0 1 3170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1677622389
transform 1 0 864 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2871
timestamp 1677622389
transform 1 0 892 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_143
timestamp 1677622389
transform 1 0 872 0 1 3170
box -8 -3 46 105
use FILL  FILL_3278
timestamp 1677622389
transform 1 0 912 0 1 3170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1677622389
transform 1 0 920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1677622389
transform 1 0 928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1677622389
transform 1 0 936 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2872
timestamp 1677622389
transform 1 0 956 0 1 3175
box -3 -3 3 3
use FILL  FILL_3288
timestamp 1677622389
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1677622389
transform 1 0 952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1677622389
transform 1 0 960 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_37
timestamp 1677622389
transform 1 0 968 0 1 3170
box -8 -3 32 105
use FILL  FILL_3292
timestamp 1677622389
transform 1 0 992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1677622389
transform 1 0 1000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1677622389
transform 1 0 1008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1677622389
transform 1 0 1016 0 1 3170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1677622389
transform 1 0 1024 0 1 3170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1677622389
transform 1 0 1032 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_249
timestamp 1677622389
transform -1 0 1056 0 1 3170
box -9 -3 26 105
use FILL  FILL_3298
timestamp 1677622389
transform 1 0 1056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1677622389
transform 1 0 1064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1677622389
transform 1 0 1072 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_69
timestamp 1677622389
transform 1 0 1080 0 1 3170
box -8 -3 34 105
use FILL  FILL_3301
timestamp 1677622389
transform 1 0 1112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1677622389
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1677622389
transform 1 0 1128 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_145
timestamp 1677622389
transform 1 0 1136 0 1 3170
box -8 -3 46 105
use FILL  FILL_3306
timestamp 1677622389
transform 1 0 1176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1677622389
transform 1 0 1184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1677622389
transform 1 0 1192 0 1 3170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1677622389
transform 1 0 1200 0 1 3170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1677622389
transform 1 0 1208 0 1 3170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1677622389
transform 1 0 1216 0 1 3170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1677622389
transform 1 0 1224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1677622389
transform 1 0 1232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1677622389
transform 1 0 1240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1677622389
transform 1 0 1248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1677622389
transform 1 0 1256 0 1 3170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1677622389
transform 1 0 1264 0 1 3170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1677622389
transform 1 0 1272 0 1 3170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1677622389
transform 1 0 1280 0 1 3170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1677622389
transform 1 0 1288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1677622389
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1677622389
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1677622389
transform 1 0 1312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1677622389
transform 1 0 1320 0 1 3170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1677622389
transform 1 0 1328 0 1 3170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1677622389
transform 1 0 1336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1677622389
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_72
timestamp 1677622389
transform -1 0 1384 0 1 3170
box -8 -3 34 105
use FILL  FILL_3341
timestamp 1677622389
transform 1 0 1384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1677622389
transform 1 0 1392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1677622389
transform 1 0 1400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1677622389
transform 1 0 1408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1677622389
transform 1 0 1416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1677622389
transform 1 0 1424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1677622389
transform 1 0 1432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1677622389
transform 1 0 1440 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_137
timestamp 1677622389
transform 1 0 1448 0 1 3170
box -8 -3 46 105
use FILL  FILL_3355
timestamp 1677622389
transform 1 0 1488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1677622389
transform 1 0 1496 0 1 3170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1677622389
transform 1 0 1504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1677622389
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1677622389
transform 1 0 1520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1677622389
transform 1 0 1528 0 1 3170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1677622389
transform 1 0 1536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1677622389
transform 1 0 1544 0 1 3170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1677622389
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_138
timestamp 1677622389
transform 1 0 1560 0 1 3170
box -8 -3 46 105
use FILL  FILL_3370
timestamp 1677622389
transform 1 0 1600 0 1 3170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1677622389
transform 1 0 1608 0 1 3170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1677622389
transform 1 0 1616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1677622389
transform 1 0 1624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1677622389
transform 1 0 1632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1677622389
transform 1 0 1640 0 1 3170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1677622389
transform 1 0 1648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1677622389
transform 1 0 1656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1677622389
transform 1 0 1664 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_140
timestamp 1677622389
transform -1 0 1712 0 1 3170
box -8 -3 46 105
use FILL  FILL_3389
timestamp 1677622389
transform 1 0 1712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1677622389
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1677622389
transform 1 0 1728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1677622389
transform 1 0 1736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1677622389
transform 1 0 1744 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_26
timestamp 1677622389
transform 1 0 1752 0 1 3170
box -5 -3 28 105
use FILL  FILL_3399
timestamp 1677622389
transform 1 0 1776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1677622389
transform 1 0 1784 0 1 3170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1677622389
transform 1 0 1792 0 1 3170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1677622389
transform 1 0 1800 0 1 3170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1677622389
transform 1 0 1808 0 1 3170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1677622389
transform 1 0 1816 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_147
timestamp 1677622389
transform 1 0 1824 0 1 3170
box -8 -3 46 105
use FILL  FILL_3411
timestamp 1677622389
transform 1 0 1864 0 1 3170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1677622389
transform 1 0 1872 0 1 3170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1677622389
transform 1 0 1880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1677622389
transform 1 0 1888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1677622389
transform 1 0 1896 0 1 3170
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1677622389
transform 1 0 1904 0 1 3170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1677622389
transform 1 0 1912 0 1 3170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1677622389
transform 1 0 1920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1677622389
transform 1 0 1928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1677622389
transform 1 0 1936 0 1 3170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1677622389
transform 1 0 1944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1677622389
transform 1 0 1952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1677622389
transform 1 0 1960 0 1 3170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1677622389
transform 1 0 1968 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_251
timestamp 1677622389
transform 1 0 1976 0 1 3170
box -9 -3 26 105
use FILL  FILL_3434
timestamp 1677622389
transform 1 0 1992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1677622389
transform 1 0 2000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1677622389
transform 1 0 2008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1677622389
transform 1 0 2016 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_252
timestamp 1677622389
transform 1 0 2024 0 1 3170
box -9 -3 26 105
use FILL  FILL_3444
timestamp 1677622389
transform 1 0 2040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1677622389
transform 1 0 2048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1677622389
transform 1 0 2056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1677622389
transform 1 0 2064 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_150
timestamp 1677622389
transform 1 0 2072 0 1 3170
box -8 -3 46 105
use FILL  FILL_3448
timestamp 1677622389
transform 1 0 2112 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_28
timestamp 1677622389
transform -1 0 2144 0 1 3170
box -5 -3 28 105
use M3_M2  M3_M2_2873
timestamp 1677622389
transform 1 0 2156 0 1 3175
box -3 -3 3 3
use BUFX2  BUFX2_29
timestamp 1677622389
transform 1 0 2144 0 1 3170
box -5 -3 28 105
use FILL  FILL_3449
timestamp 1677622389
transform 1 0 2168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1677622389
transform 1 0 2176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1677622389
transform 1 0 2184 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_151
timestamp 1677622389
transform 1 0 2192 0 1 3170
box -8 -3 46 105
use FILL  FILL_3464
timestamp 1677622389
transform 1 0 2232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1677622389
transform 1 0 2240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1677622389
transform 1 0 2248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1677622389
transform 1 0 2256 0 1 3170
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1677622389
transform 1 0 2264 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_254
timestamp 1677622389
transform 1 0 2272 0 1 3170
box -9 -3 26 105
use FILL  FILL_3473
timestamp 1677622389
transform 1 0 2288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1677622389
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1677622389
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1677622389
transform 1 0 2312 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_152
timestamp 1677622389
transform 1 0 2320 0 1 3170
box -8 -3 46 105
use FILL  FILL_3483
timestamp 1677622389
transform 1 0 2360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1677622389
transform 1 0 2368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1677622389
transform 1 0 2376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1677622389
transform 1 0 2384 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_144
timestamp 1677622389
transform -1 0 2432 0 1 3170
box -8 -3 46 105
use FILL  FILL_3495
timestamp 1677622389
transform 1 0 2432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1677622389
transform 1 0 2440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1677622389
transform 1 0 2448 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_153
timestamp 1677622389
transform 1 0 2456 0 1 3170
box -8 -3 46 105
use FILL  FILL_3501
timestamp 1677622389
transform 1 0 2496 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2874
timestamp 1677622389
transform 1 0 2516 0 1 3175
box -3 -3 3 3
use FILL  FILL_3502
timestamp 1677622389
transform 1 0 2504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1677622389
transform 1 0 2512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1677622389
transform 1 0 2520 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2875
timestamp 1677622389
transform 1 0 2548 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_227
timestamp 1677622389
transform 1 0 2528 0 1 3170
box -8 -3 104 105
use FILL  FILL_3505
timestamp 1677622389
transform 1 0 2624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1677622389
transform 1 0 2632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1677622389
transform 1 0 2640 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2876
timestamp 1677622389
transform 1 0 2660 0 1 3175
box -3 -3 3 3
use FILL  FILL_3508
timestamp 1677622389
transform 1 0 2648 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2877
timestamp 1677622389
transform 1 0 2700 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_154
timestamp 1677622389
transform 1 0 2656 0 1 3170
box -8 -3 46 105
use FILL  FILL_3509
timestamp 1677622389
transform 1 0 2696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1677622389
transform 1 0 2704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1677622389
transform 1 0 2712 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_258
timestamp 1677622389
transform 1 0 2720 0 1 3170
box -9 -3 26 105
use FILL  FILL_3529
timestamp 1677622389
transform 1 0 2736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1677622389
transform 1 0 2744 0 1 3170
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1677622389
transform 1 0 2752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1677622389
transform 1 0 2760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1677622389
transform 1 0 2768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1677622389
transform 1 0 2776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1677622389
transform 1 0 2784 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1677622389
transform 1 0 2792 0 1 3170
box -8 -3 34 105
use FILL  FILL_3536
timestamp 1677622389
transform 1 0 2824 0 1 3170
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1677622389
transform 1 0 2832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1677622389
transform 1 0 2840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1677622389
transform 1 0 2848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1677622389
transform 1 0 2856 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_75
timestamp 1677622389
transform 1 0 2864 0 1 3170
box -8 -3 34 105
use FILL  FILL_3546
timestamp 1677622389
transform 1 0 2896 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_38
timestamp 1677622389
transform 1 0 2904 0 1 3170
box -8 -3 32 105
use FILL  FILL_3550
timestamp 1677622389
transform 1 0 2928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1677622389
transform 1 0 2936 0 1 3170
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1677622389
transform 1 0 2944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1677622389
transform 1 0 2952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1677622389
transform 1 0 2960 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_77
timestamp 1677622389
transform -1 0 3000 0 1 3170
box -8 -3 34 105
use FILL  FILL_3559
timestamp 1677622389
transform 1 0 3000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1677622389
transform 1 0 3008 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_259
timestamp 1677622389
transform -1 0 3032 0 1 3170
box -9 -3 26 105
use FILL  FILL_3561
timestamp 1677622389
transform 1 0 3032 0 1 3170
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1677622389
transform 1 0 3040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1677622389
transform 1 0 3048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1677622389
transform 1 0 3056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1677622389
transform 1 0 3064 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_146
timestamp 1677622389
transform -1 0 3112 0 1 3170
box -8 -3 46 105
use FILL  FILL_3575
timestamp 1677622389
transform 1 0 3112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1677622389
transform 1 0 3120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1677622389
transform 1 0 3128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1677622389
transform 1 0 3136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1677622389
transform 1 0 3144 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2878
timestamp 1677622389
transform 1 0 3164 0 1 3175
box -3 -3 3 3
use OAI22X1  OAI22X1_147
timestamp 1677622389
transform -1 0 3192 0 1 3170
box -8 -3 46 105
use FILL  FILL_3583
timestamp 1677622389
transform 1 0 3192 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2879
timestamp 1677622389
transform 1 0 3212 0 1 3175
box -3 -3 3 3
use FILL  FILL_3584
timestamp 1677622389
transform 1 0 3200 0 1 3170
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1677622389
transform 1 0 3208 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1677622389
transform -1 0 3312 0 1 3170
box -8 -3 104 105
use FILL  FILL_3586
timestamp 1677622389
transform 1 0 3312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1677622389
transform 1 0 3320 0 1 3170
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1677622389
transform 1 0 3328 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_18
timestamp 1677622389
transform -1 0 3368 0 1 3170
box -8 -3 40 105
use FILL  FILL_3608
timestamp 1677622389
transform 1 0 3368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1677622389
transform 1 0 3376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1677622389
transform 1 0 3384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1677622389
transform 1 0 3392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1677622389
transform 1 0 3400 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_19
timestamp 1677622389
transform -1 0 3440 0 1 3170
box -8 -3 40 105
use FILL  FILL_3613
timestamp 1677622389
transform 1 0 3440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1677622389
transform 1 0 3448 0 1 3170
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1677622389
transform 1 0 3456 0 1 3170
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1677622389
transform 1 0 3464 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_20
timestamp 1677622389
transform -1 0 3504 0 1 3170
box -8 -3 40 105
use FILL  FILL_3617
timestamp 1677622389
transform 1 0 3504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1677622389
transform 1 0 3512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1677622389
transform 1 0 3520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1677622389
transform 1 0 3528 0 1 3170
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1677622389
transform 1 0 3536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1677622389
transform 1 0 3544 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1677622389
transform -1 0 3584 0 1 3170
box -8 -3 40 105
use FILL  FILL_3623
timestamp 1677622389
transform 1 0 3584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1677622389
transform 1 0 3592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1677622389
transform 1 0 3600 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_262
timestamp 1677622389
transform 1 0 3608 0 1 3170
box -9 -3 26 105
use FILL  FILL_3635
timestamp 1677622389
transform 1 0 3624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1677622389
transform 1 0 3632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1677622389
transform 1 0 3640 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_157
timestamp 1677622389
transform -1 0 3688 0 1 3170
box -8 -3 46 105
use FILL  FILL_3640
timestamp 1677622389
transform 1 0 3688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1677622389
transform 1 0 3696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1677622389
transform 1 0 3704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1677622389
transform 1 0 3712 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_158
timestamp 1677622389
transform 1 0 3720 0 1 3170
box -8 -3 46 105
use FILL  FILL_3649
timestamp 1677622389
transform 1 0 3760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1677622389
transform 1 0 3768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1677622389
transform 1 0 3776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1677622389
transform 1 0 3784 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_159
timestamp 1677622389
transform 1 0 3792 0 1 3170
box -8 -3 46 105
use FILL  FILL_3656
timestamp 1677622389
transform 1 0 3832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1677622389
transform 1 0 3840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1677622389
transform 1 0 3848 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_31
timestamp 1677622389
transform 1 0 3856 0 1 3170
box -5 -3 28 105
use FILL  FILL_3659
timestamp 1677622389
transform 1 0 3880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1677622389
transform 1 0 3888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1677622389
transform 1 0 3896 0 1 3170
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1677622389
transform 1 0 3904 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_151
timestamp 1677622389
transform 1 0 3912 0 1 3170
box -8 -3 46 105
use FILL  FILL_3665
timestamp 1677622389
transform 1 0 3952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1677622389
transform 1 0 3960 0 1 3170
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1677622389
transform 1 0 3968 0 1 3170
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1677622389
transform 1 0 3976 0 1 3170
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1677622389
transform 1 0 3984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1677622389
transform 1 0 3992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1677622389
transform 1 0 4000 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_265
timestamp 1677622389
transform 1 0 4008 0 1 3170
box -9 -3 26 105
use FILL  FILL_3672
timestamp 1677622389
transform 1 0 4024 0 1 3170
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1677622389
transform 1 0 4032 0 1 3170
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1677622389
transform 1 0 4040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1677622389
transform 1 0 4048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1677622389
transform 1 0 4056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1677622389
transform 1 0 4064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1677622389
transform 1 0 4072 0 1 3170
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1677622389
transform 1 0 4080 0 1 3170
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1677622389
transform 1 0 4088 0 1 3170
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1677622389
transform 1 0 4096 0 1 3170
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1677622389
transform 1 0 4104 0 1 3170
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1677622389
transform 1 0 4112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1677622389
transform 1 0 4120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1677622389
transform 1 0 4128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1677622389
transform 1 0 4136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1677622389
transform 1 0 4144 0 1 3170
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1677622389
transform 1 0 4152 0 1 3170
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1677622389
transform 1 0 4160 0 1 3170
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1677622389
transform 1 0 4168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1677622389
transform 1 0 4176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1677622389
transform 1 0 4184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1677622389
transform 1 0 4192 0 1 3170
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1677622389
transform 1 0 4200 0 1 3170
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1677622389
transform 1 0 4208 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_234
timestamp 1677622389
transform 1 0 4216 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_266
timestamp 1677622389
transform 1 0 4312 0 1 3170
box -9 -3 26 105
use FILL  FILL_3710
timestamp 1677622389
transform 1 0 4328 0 1 3170
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1677622389
transform 1 0 4336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1677622389
transform 1 0 4344 0 1 3170
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1677622389
transform 1 0 4352 0 1 3170
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1677622389
transform 1 0 4360 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_155
timestamp 1677622389
transform 1 0 4368 0 1 3170
box -8 -3 46 105
use FILL  FILL_3726
timestamp 1677622389
transform 1 0 4408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1677622389
transform 1 0 4416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1677622389
transform 1 0 4424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1677622389
transform 1 0 4432 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_33
timestamp 1677622389
transform 1 0 4440 0 1 3170
box -5 -3 28 105
use FILL  FILL_3736
timestamp 1677622389
transform 1 0 4464 0 1 3170
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1677622389
transform 1 0 4472 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_156
timestamp 1677622389
transform 1 0 4480 0 1 3170
box -8 -3 46 105
use FILL  FILL_3738
timestamp 1677622389
transform 1 0 4520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1677622389
transform 1 0 4528 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2880
timestamp 1677622389
transform 1 0 4548 0 1 3175
box -3 -3 3 3
use FILL  FILL_3746
timestamp 1677622389
transform 1 0 4536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1677622389
transform 1 0 4544 0 1 3170
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1677622389
transform 1 0 4552 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2881
timestamp 1677622389
transform 1 0 4572 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_235
timestamp 1677622389
transform 1 0 4560 0 1 3170
box -8 -3 104 105
use OAI22X1  OAI22X1_157
timestamp 1677622389
transform 1 0 4656 0 1 3170
box -8 -3 46 105
use FILL  FILL_3757
timestamp 1677622389
transform 1 0 4696 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_271
timestamp 1677622389
transform 1 0 4704 0 1 3170
box -9 -3 26 105
use FILL  FILL_3758
timestamp 1677622389
transform 1 0 4720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1677622389
transform 1 0 4728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1677622389
transform 1 0 4736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1677622389
transform 1 0 4744 0 1 3170
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1677622389
transform 1 0 4752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1677622389
transform 1 0 4760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1677622389
transform 1 0 4768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1677622389
transform 1 0 4776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1677622389
transform 1 0 4784 0 1 3170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_31
timestamp 1677622389
transform 1 0 4819 0 1 3170
box -10 -3 10 3
use M2_M1  M2_M1_3266
timestamp 1677622389
transform 1 0 100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1677622389
transform 1 0 148 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3001
timestamp 1677622389
transform 1 0 148 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1677622389
transform 1 0 172 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3373
timestamp 1677622389
transform 1 0 196 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2954
timestamp 1677622389
transform 1 0 212 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1677622389
transform 1 0 244 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3267
timestamp 1677622389
transform 1 0 220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1677622389
transform 1 0 236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1677622389
transform 1 0 212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1677622389
transform 1 0 228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1677622389
transform 1 0 244 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3031
timestamp 1677622389
transform 1 0 244 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1677622389
transform 1 0 268 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1677622389
transform 1 0 284 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1677622389
transform 1 0 316 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3269
timestamp 1677622389
transform 1 0 316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1677622389
transform 1 0 364 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2900
timestamp 1677622389
transform 1 0 420 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3378
timestamp 1677622389
transform 1 0 420 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1677622389
transform 1 0 476 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3003
timestamp 1677622389
transform 1 0 476 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3379
timestamp 1677622389
transform 1 0 508 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2922
timestamp 1677622389
transform 1 0 548 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1677622389
transform 1 0 564 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3271
timestamp 1677622389
transform 1 0 548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1677622389
transform 1 0 572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1677622389
transform 1 0 548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1677622389
transform 1 0 564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1677622389
transform 1 0 580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3004
timestamp 1677622389
transform 1 0 564 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1677622389
transform 1 0 580 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1677622389
transform 1 0 548 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1677622389
transform 1 0 564 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3383
timestamp 1677622389
transform 1 0 620 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2924
timestamp 1677622389
transform 1 0 644 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3273
timestamp 1677622389
transform 1 0 644 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2981
timestamp 1677622389
transform 1 0 636 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1677622389
transform 1 0 676 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1677622389
transform 1 0 668 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1677622389
transform 1 0 780 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3263
timestamp 1677622389
transform 1 0 828 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_2926
timestamp 1677622389
transform 1 0 836 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3264
timestamp 1677622389
transform 1 0 844 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1677622389
transform 1 0 668 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1677622389
transform 1 0 684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1677622389
transform 1 0 700 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1677622389
transform 1 0 788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1677622389
transform 1 0 796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1677622389
transform 1 0 812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1677622389
transform 1 0 828 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1677622389
transform 1 0 652 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2982
timestamp 1677622389
transform 1 0 668 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3385
timestamp 1677622389
transform 1 0 676 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2983
timestamp 1677622389
transform 1 0 684 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3386
timestamp 1677622389
transform 1 0 724 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2984
timestamp 1677622389
transform 1 0 748 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3387
timestamp 1677622389
transform 1 0 780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1677622389
transform 1 0 804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1677622389
transform 1 0 820 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3066
timestamp 1677622389
transform 1 0 788 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1677622389
transform 1 0 820 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1677622389
transform 1 0 884 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1677622389
transform 1 0 884 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3281
timestamp 1677622389
transform 1 0 876 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2985
timestamp 1677622389
transform 1 0 876 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3390
timestamp 1677622389
transform 1 0 884 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1677622389
transform 1 0 900 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2903
timestamp 1677622389
transform 1 0 916 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3283
timestamp 1677622389
transform 1 0 916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1677622389
transform 1 0 916 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2928
timestamp 1677622389
transform 1 0 980 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1677622389
transform 1 0 1012 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1677622389
transform 1 0 1052 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1677622389
transform 1 0 1068 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1677622389
transform 1 0 1108 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3284
timestamp 1677622389
transform 1 0 980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1677622389
transform 1 0 996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1677622389
transform 1 0 1012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1677622389
transform 1 0 1020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1677622389
transform 1 0 1036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1677622389
transform 1 0 956 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3067
timestamp 1677622389
transform 1 0 948 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1677622389
transform 1 0 972 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3393
timestamp 1677622389
transform 1 0 980 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2987
timestamp 1677622389
transform 1 0 988 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3394
timestamp 1677622389
transform 1 0 1004 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2988
timestamp 1677622389
transform 1 0 1020 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3395
timestamp 1677622389
transform 1 0 1060 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1677622389
transform 1 0 979 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3007
timestamp 1677622389
transform 1 0 988 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1677622389
transform 1 0 964 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1677622389
transform 1 0 1004 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1677622389
transform 1 0 1020 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1677622389
transform 1 0 1148 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1677622389
transform 1 0 1180 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1677622389
transform 1 0 1156 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1677622389
transform 1 0 1188 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3289
timestamp 1677622389
transform 1 0 1180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1677622389
transform 1 0 1188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1677622389
transform 1 0 1148 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1677622389
transform 1 0 1156 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2989
timestamp 1677622389
transform 1 0 1164 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3398
timestamp 1677622389
transform 1 0 1172 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3008
timestamp 1677622389
transform 1 0 1188 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1677622389
transform 1 0 1188 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1677622389
transform 1 0 1156 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1677622389
transform 1 0 1172 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1677622389
transform 1 0 1220 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3399
timestamp 1677622389
transform 1 0 1220 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3051
timestamp 1677622389
transform 1 0 1212 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1677622389
transform 1 0 1252 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3400
timestamp 1677622389
transform 1 0 1252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1677622389
transform 1 0 1252 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3052
timestamp 1677622389
transform 1 0 1252 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1677622389
transform 1 0 1276 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1677622389
transform 1 0 1292 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3291
timestamp 1677622389
transform 1 0 1292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1677622389
transform 1 0 1300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1677622389
transform 1 0 1292 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3009
timestamp 1677622389
transform 1 0 1292 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3483
timestamp 1677622389
transform 1 0 1316 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1677622389
transform 1 0 1340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1677622389
transform 1 0 1324 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3053
timestamp 1677622389
transform 1 0 1316 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1677622389
transform 1 0 1340 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3403
timestamp 1677622389
transform 1 0 1372 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2906
timestamp 1677622389
transform 1 0 1388 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3293
timestamp 1677622389
transform 1 0 1388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1677622389
transform 1 0 1404 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2956
timestamp 1677622389
transform 1 0 1444 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3404
timestamp 1677622389
transform 1 0 1444 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2907
timestamp 1677622389
transform 1 0 1516 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3295
timestamp 1677622389
transform 1 0 1524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1677622389
transform 1 0 1516 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2908
timestamp 1677622389
transform 1 0 1540 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3406
timestamp 1677622389
transform 1 0 1556 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2909
timestamp 1677622389
transform 1 0 1596 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1677622389
transform 1 0 1572 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3296
timestamp 1677622389
transform 1 0 1580 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2958
timestamp 1677622389
transform 1 0 1596 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3407
timestamp 1677622389
transform 1 0 1572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1677622389
transform 1 0 1596 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3011
timestamp 1677622389
transform 1 0 1596 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3297
timestamp 1677622389
transform 1 0 1644 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2888
timestamp 1677622389
transform 1 0 1684 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3298
timestamp 1677622389
transform 1 0 1676 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1677622389
transform 1 0 1692 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2959
timestamp 1677622389
transform 1 0 1700 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3409
timestamp 1677622389
transform 1 0 1684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1677622389
transform 1 0 1700 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1677622389
transform 1 0 1724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1677622389
transform 1 0 1748 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2889
timestamp 1677622389
transform 1 0 1772 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3301
timestamp 1677622389
transform 1 0 1772 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3036
timestamp 1677622389
transform 1 0 1812 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1677622389
transform 1 0 1836 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1677622389
transform 1 0 1868 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3302
timestamp 1677622389
transform 1 0 1836 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2960
timestamp 1677622389
transform 1 0 1860 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3412
timestamp 1677622389
transform 1 0 1828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1677622389
transform 1 0 1844 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1677622389
transform 1 0 1860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1677622389
transform 1 0 1868 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3037
timestamp 1677622389
transform 1 0 1860 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1677622389
transform 1 0 1940 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3303
timestamp 1677622389
transform 1 0 1932 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1677622389
transform 1 0 1940 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2961
timestamp 1677622389
transform 1 0 1972 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3416
timestamp 1677622389
transform 1 0 1940 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1677622389
transform 1 0 1956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1677622389
transform 1 0 1972 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3038
timestamp 1677622389
transform 1 0 1932 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1677622389
transform 1 0 1956 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1677622389
transform 1 0 2004 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1677622389
transform 1 0 2052 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1677622389
transform 1 0 2044 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1677622389
transform 1 0 2036 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3305
timestamp 1677622389
transform 1 0 2028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1677622389
transform 1 0 2060 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2962
timestamp 1677622389
transform 1 0 2068 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3419
timestamp 1677622389
transform 1 0 2052 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1677622389
transform 1 0 2068 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2963
timestamp 1677622389
transform 1 0 2084 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3307
timestamp 1677622389
transform 1 0 2092 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3055
timestamp 1677622389
transform 1 0 2076 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1677622389
transform 1 0 2052 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1677622389
transform 1 0 2076 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1677622389
transform 1 0 2124 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3421
timestamp 1677622389
transform 1 0 2124 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2965
timestamp 1677622389
transform 1 0 2140 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3308
timestamp 1677622389
transform 1 0 2156 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2990
timestamp 1677622389
transform 1 0 2156 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1677622389
transform 1 0 2172 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3309
timestamp 1677622389
transform 1 0 2172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1677622389
transform 1 0 2180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1677622389
transform 1 0 2204 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3056
timestamp 1677622389
transform 1 0 2204 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1677622389
transform 1 0 2220 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1677622389
transform 1 0 2244 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3310
timestamp 1677622389
transform 1 0 2228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1677622389
transform 1 0 2244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1677622389
transform 1 0 2252 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2937
timestamp 1677622389
transform 1 0 2268 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3312
timestamp 1677622389
transform 1 0 2268 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3040
timestamp 1677622389
transform 1 0 2316 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1677622389
transform 1 0 2372 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1677622389
transform 1 0 2428 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3313
timestamp 1677622389
transform 1 0 2388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1677622389
transform 1 0 2404 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1677622389
transform 1 0 2420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1677622389
transform 1 0 2428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1677622389
transform 1 0 2380 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3057
timestamp 1677622389
transform 1 0 2380 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3426
timestamp 1677622389
transform 1 0 2412 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3058
timestamp 1677622389
transform 1 0 2404 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3317
timestamp 1677622389
transform 1 0 2468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1677622389
transform 1 0 2460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1677622389
transform 1 0 2468 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2940
timestamp 1677622389
transform 1 0 2508 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3318
timestamp 1677622389
transform 1 0 2508 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1677622389
transform 1 0 2524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1677622389
transform 1 0 2532 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1677622389
transform 1 0 2516 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2966
timestamp 1677622389
transform 1 0 2540 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3430
timestamp 1677622389
transform 1 0 2548 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2941
timestamp 1677622389
transform 1 0 2580 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3321
timestamp 1677622389
transform 1 0 2580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1677622389
transform 1 0 2572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1677622389
transform 1 0 2580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3041
timestamp 1677622389
transform 1 0 2580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1677622389
transform 1 0 2604 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1677622389
transform 1 0 2620 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3322
timestamp 1677622389
transform 1 0 2628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1677622389
transform 1 0 2644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1677622389
transform 1 0 2652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1677622389
transform 1 0 2636 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3042
timestamp 1677622389
transform 1 0 2644 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3434
timestamp 1677622389
transform 1 0 2660 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2968
timestamp 1677622389
transform 1 0 2708 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3435
timestamp 1677622389
transform 1 0 2708 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2943
timestamp 1677622389
transform 1 0 2724 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3325
timestamp 1677622389
transform 1 0 2724 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2969
timestamp 1677622389
transform 1 0 2748 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3436
timestamp 1677622389
transform 1 0 2748 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1677622389
transform 1 0 2804 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3043
timestamp 1677622389
transform 1 0 2804 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1677622389
transform 1 0 2836 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1677622389
transform 1 0 2860 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3438
timestamp 1677622389
transform 1 0 2860 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2915
timestamp 1677622389
transform 1 0 2884 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3265
timestamp 1677622389
transform 1 0 2884 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_3059
timestamp 1677622389
transform 1 0 2908 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3326
timestamp 1677622389
transform 1 0 2924 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2992
timestamp 1677622389
transform 1 0 2932 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3485
timestamp 1677622389
transform 1 0 2932 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1677622389
transform 1 0 2956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1677622389
transform 1 0 2980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1677622389
transform 1 0 2988 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1677622389
transform 1 0 2972 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3060
timestamp 1677622389
transform 1 0 2972 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1677622389
transform 1 0 3028 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1677622389
transform 1 0 3020 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3329
timestamp 1677622389
transform 1 0 3028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1677622389
transform 1 0 3036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1677622389
transform 1 0 3020 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2993
timestamp 1677622389
transform 1 0 3036 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3487
timestamp 1677622389
transform 1 0 3036 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3061
timestamp 1677622389
transform 1 0 3036 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1677622389
transform 1 0 3092 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3441
timestamp 1677622389
transform 1 0 3092 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1677622389
transform 1 0 3180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1677622389
transform 1 0 3188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1677622389
transform 1 0 3204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1677622389
transform 1 0 3220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1677622389
transform 1 0 3180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1677622389
transform 1 0 3196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1677622389
transform 1 0 3212 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3012
timestamp 1677622389
transform 1 0 3268 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1677622389
transform 1 0 3292 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1677622389
transform 1 0 3284 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3335
timestamp 1677622389
transform 1 0 3292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1677622389
transform 1 0 3284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1677622389
transform 1 0 3300 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1677622389
transform 1 0 3364 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2994
timestamp 1677622389
transform 1 0 3364 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1677622389
transform 1 0 3380 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3337
timestamp 1677622389
transform 1 0 3380 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2973
timestamp 1677622389
transform 1 0 3412 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3446
timestamp 1677622389
transform 1 0 3412 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1677622389
transform 1 0 3420 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1677622389
transform 1 0 3412 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3447
timestamp 1677622389
transform 1 0 3492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1677622389
transform 1 0 3508 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2974
timestamp 1677622389
transform 1 0 3548 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3448
timestamp 1677622389
transform 1 0 3556 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3013
timestamp 1677622389
transform 1 0 3556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1677622389
transform 1 0 3516 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1677622389
transform 1 0 3636 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3339
timestamp 1677622389
transform 1 0 3628 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2975
timestamp 1677622389
transform 1 0 3636 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3449
timestamp 1677622389
transform 1 0 3636 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2894
timestamp 1677622389
transform 1 0 3700 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1677622389
transform 1 0 3692 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3340
timestamp 1677622389
transform 1 0 3676 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2976
timestamp 1677622389
transform 1 0 3684 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3341
timestamp 1677622389
transform 1 0 3692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1677622389
transform 1 0 3700 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1677622389
transform 1 0 3668 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1677622389
transform 1 0 3684 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3014
timestamp 1677622389
transform 1 0 3676 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1677622389
transform 1 0 3668 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1677622389
transform 1 0 3716 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3452
timestamp 1677622389
transform 1 0 3708 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3045
timestamp 1677622389
transform 1 0 3708 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1677622389
transform 1 0 3764 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3343
timestamp 1677622389
transform 1 0 3732 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1677622389
transform 1 0 3748 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1677622389
transform 1 0 3764 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2996
timestamp 1677622389
transform 1 0 3732 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3453
timestamp 1677622389
transform 1 0 3756 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3015
timestamp 1677622389
transform 1 0 3748 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1677622389
transform 1 0 3772 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1677622389
transform 1 0 3844 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1677622389
transform 1 0 3860 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3346
timestamp 1677622389
transform 1 0 3796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1677622389
transform 1 0 3820 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2978
timestamp 1677622389
transform 1 0 3892 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3455
timestamp 1677622389
transform 1 0 3892 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3016
timestamp 1677622389
transform 1 0 3820 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1677622389
transform 1 0 3876 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1677622389
transform 1 0 3892 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1677622389
transform 1 0 3876 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1677622389
transform 1 0 3900 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1677622389
transform 1 0 3916 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3347
timestamp 1677622389
transform 1 0 3948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1677622389
transform 1 0 3972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1677622389
transform 1 0 4028 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3018
timestamp 1677622389
transform 1 0 3988 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3348
timestamp 1677622389
transform 1 0 4044 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2946
timestamp 1677622389
transform 1 0 4060 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1677622389
transform 1 0 4116 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1677622389
transform 1 0 4108 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3349
timestamp 1677622389
transform 1 0 4076 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1677622389
transform 1 0 4092 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1677622389
transform 1 0 4108 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1677622389
transform 1 0 4084 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1677622389
transform 1 0 4100 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3019
timestamp 1677622389
transform 1 0 4100 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1677622389
transform 1 0 4100 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3352
timestamp 1677622389
transform 1 0 4124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1677622389
transform 1 0 4116 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2997
timestamp 1677622389
transform 1 0 4124 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3461
timestamp 1677622389
transform 1 0 4148 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3063
timestamp 1677622389
transform 1 0 4140 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1677622389
transform 1 0 4164 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1677622389
transform 1 0 4188 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3353
timestamp 1677622389
transform 1 0 4180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1677622389
transform 1 0 4188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1677622389
transform 1 0 4204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1677622389
transform 1 0 4220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1677622389
transform 1 0 4172 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3020
timestamp 1677622389
transform 1 0 4172 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3463
timestamp 1677622389
transform 1 0 4212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1677622389
transform 1 0 4228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1677622389
transform 1 0 4276 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3047
timestamp 1677622389
transform 1 0 4276 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1677622389
transform 1 0 4324 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3357
timestamp 1677622389
transform 1 0 4316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1677622389
transform 1 0 4324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1677622389
transform 1 0 4340 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2999
timestamp 1677622389
transform 1 0 4308 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1677622389
transform 1 0 4316 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3466
timestamp 1677622389
transform 1 0 4332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1677622389
transform 1 0 4348 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3022
timestamp 1677622389
transform 1 0 4348 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3468
timestamp 1677622389
transform 1 0 4364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1677622389
transform 1 0 4372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1677622389
transform 1 0 4404 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3023
timestamp 1677622389
transform 1 0 4404 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3469
timestamp 1677622389
transform 1 0 4420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2950
timestamp 1677622389
transform 1 0 4452 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3362
timestamp 1677622389
transform 1 0 4452 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2980
timestamp 1677622389
transform 1 0 4484 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3470
timestamp 1677622389
transform 1 0 4460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1677622389
transform 1 0 4476 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3024
timestamp 1677622389
transform 1 0 4452 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3472
timestamp 1677622389
transform 1 0 4516 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3025
timestamp 1677622389
transform 1 0 4516 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3363
timestamp 1677622389
transform 1 0 4532 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3048
timestamp 1677622389
transform 1 0 4532 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1677622389
transform 1 0 4580 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1677622389
transform 1 0 4588 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3364
timestamp 1677622389
transform 1 0 4548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1677622389
transform 1 0 4564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1677622389
transform 1 0 4580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1677622389
transform 1 0 4556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1677622389
transform 1 0 4572 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3000
timestamp 1677622389
transform 1 0 4580 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3475
timestamp 1677622389
transform 1 0 4588 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3026
timestamp 1677622389
transform 1 0 4556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1677622389
transform 1 0 4572 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1677622389
transform 1 0 4580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1677622389
transform 1 0 4548 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1677622389
transform 1 0 4572 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1677622389
transform 1 0 4604 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1677622389
transform 1 0 4660 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1677622389
transform 1 0 4660 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1677622389
transform 1 0 4676 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1677622389
transform 1 0 4732 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3367
timestamp 1677622389
transform 1 0 4652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1677622389
transform 1 0 4660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1677622389
transform 1 0 4676 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1677622389
transform 1 0 4692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1677622389
transform 1 0 4708 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1677622389
transform 1 0 4660 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1677622389
transform 1 0 4668 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1677622389
transform 1 0 4684 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3029
timestamp 1677622389
transform 1 0 4660 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1677622389
transform 1 0 4684 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1677622389
transform 1 0 4652 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_3479
timestamp 1677622389
transform 1 0 4732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1677622389
transform 1 0 4788 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3079
timestamp 1677622389
transform 1 0 4788 0 1 3085
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_32
timestamp 1677622389
transform 1 0 24 0 1 3070
box -10 -3 10 3
use FILL  FILL_3207
timestamp 1677622389
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1677622389
transform 1 0 80 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_220
timestamp 1677622389
transform 1 0 88 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3209
timestamp 1677622389
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1677622389
transform 1 0 192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1677622389
transform 1 0 200 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_138
timestamp 1677622389
transform 1 0 208 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3212
timestamp 1677622389
transform 1 0 248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1677622389
transform 1 0 256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1677622389
transform 1 0 264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1677622389
transform 1 0 272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1677622389
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1677622389
transform 1 0 288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1677622389
transform 1 0 296 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1677622389
transform 1 0 304 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3224
timestamp 1677622389
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1677622389
transform 1 0 408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1677622389
transform 1 0 416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1677622389
transform 1 0 424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1677622389
transform 1 0 432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1677622389
transform 1 0 440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1677622389
transform 1 0 448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1677622389
transform 1 0 456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1677622389
transform 1 0 464 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_246
timestamp 1677622389
transform 1 0 472 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3239
timestamp 1677622389
transform 1 0 488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1677622389
transform 1 0 496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1677622389
transform 1 0 504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1677622389
transform 1 0 512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1677622389
transform 1 0 520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1677622389
transform 1 0 528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1677622389
transform 1 0 536 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_140
timestamp 1677622389
transform -1 0 584 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3246
timestamp 1677622389
transform 1 0 584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1677622389
transform 1 0 592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1677622389
transform 1 0 600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1677622389
transform 1 0 608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1677622389
transform 1 0 616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1677622389
transform 1 0 624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1677622389
transform 1 0 632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1677622389
transform 1 0 640 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3080
timestamp 1677622389
transform 1 0 676 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_136
timestamp 1677622389
transform 1 0 648 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1677622389
transform 1 0 688 0 -1 3170
box -8 -3 104 105
use AOI22X1  AOI22X1_142
timestamp 1677622389
transform -1 0 824 0 -1 3170
box -8 -3 46 105
use NOR2X1  NOR2X1_35
timestamp 1677622389
transform 1 0 824 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3273
timestamp 1677622389
transform 1 0 848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1677622389
transform 1 0 856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1677622389
transform 1 0 864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1677622389
transform 1 0 872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1677622389
transform 1 0 880 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_36
timestamp 1677622389
transform 1 0 888 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3281
timestamp 1677622389
transform 1 0 912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1677622389
transform 1 0 920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1677622389
transform 1 0 928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1677622389
transform 1 0 936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1677622389
transform 1 0 944 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_70
timestamp 1677622389
transform 1 0 952 0 -1 3170
box -8 -3 34 105
use AOI22X1  AOI22X1_144
timestamp 1677622389
transform 1 0 984 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1677622389
transform 1 0 1024 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3303
timestamp 1677622389
transform 1 0 1120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1677622389
transform 1 0 1128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1677622389
transform 1 0 1136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1677622389
transform 1 0 1144 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_146
timestamp 1677622389
transform -1 0 1192 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3311
timestamp 1677622389
transform 1 0 1192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1677622389
transform 1 0 1200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1677622389
transform 1 0 1208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1677622389
transform 1 0 1216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1677622389
transform 1 0 1224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1677622389
transform 1 0 1232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1677622389
transform 1 0 1240 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_71
timestamp 1677622389
transform -1 0 1280 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3329
timestamp 1677622389
transform 1 0 1280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1677622389
transform 1 0 1288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1677622389
transform 1 0 1296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1677622389
transform 1 0 1304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1677622389
transform 1 0 1312 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_73
timestamp 1677622389
transform -1 0 1352 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3343
timestamp 1677622389
transform 1 0 1352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1677622389
transform 1 0 1360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1677622389
transform 1 0 1368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1677622389
transform 1 0 1376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1677622389
transform 1 0 1384 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1677622389
transform 1 0 1392 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3356
timestamp 1677622389
transform 1 0 1488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1677622389
transform 1 0 1496 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_250
timestamp 1677622389
transform 1 0 1504 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3362
timestamp 1677622389
transform 1 0 1520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1677622389
transform 1 0 1528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1677622389
transform 1 0 1536 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1677622389
transform 1 0 1544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1677622389
transform 1 0 1552 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_139
timestamp 1677622389
transform -1 0 1600 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3372
timestamp 1677622389
transform 1 0 1600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1677622389
transform 1 0 1608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1677622389
transform 1 0 1616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1677622389
transform 1 0 1624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1677622389
transform 1 0 1632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1677622389
transform 1 0 1640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1677622389
transform 1 0 1648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1677622389
transform 1 0 1656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1677622389
transform 1 0 1664 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_141
timestamp 1677622389
transform -1 0 1712 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3390
timestamp 1677622389
transform 1 0 1712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1677622389
transform 1 0 1720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1677622389
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1677622389
transform 1 0 1736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1677622389
transform 1 0 1744 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3081
timestamp 1677622389
transform 1 0 1772 0 1 3075
box -3 -3 3 3
use BUFX2  BUFX2_27
timestamp 1677622389
transform 1 0 1752 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3400
timestamp 1677622389
transform 1 0 1776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1677622389
transform 1 0 1784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1677622389
transform 1 0 1792 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1677622389
transform 1 0 1800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1677622389
transform 1 0 1808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1677622389
transform 1 0 1816 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_148
timestamp 1677622389
transform 1 0 1824 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3412
timestamp 1677622389
transform 1 0 1864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1677622389
transform 1 0 1872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1677622389
transform 1 0 1880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1677622389
transform 1 0 1888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1677622389
transform 1 0 1896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1677622389
transform 1 0 1904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1677622389
transform 1 0 1912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1677622389
transform 1 0 1920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1677622389
transform 1 0 1928 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_149
timestamp 1677622389
transform 1 0 1936 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3435
timestamp 1677622389
transform 1 0 1976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1677622389
transform 1 0 1984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1677622389
transform 1 0 1992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1677622389
transform 1 0 2000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1677622389
transform 1 0 2008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1677622389
transform 1 0 2016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1677622389
transform 1 0 2024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1677622389
transform 1 0 2032 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_142
timestamp 1677622389
transform -1 0 2080 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3452
timestamp 1677622389
transform 1 0 2080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1677622389
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1677622389
transform 1 0 2096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1677622389
transform 1 0 2104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1677622389
transform 1 0 2112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1677622389
transform 1 0 2120 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_30
timestamp 1677622389
transform 1 0 2128 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3458
timestamp 1677622389
transform 1 0 2152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1677622389
transform 1 0 2160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1677622389
transform 1 0 2168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1677622389
transform 1 0 2176 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_253
timestamp 1677622389
transform 1 0 2184 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3469
timestamp 1677622389
transform 1 0 2200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1677622389
transform 1 0 2208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1677622389
transform 1 0 2216 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3082
timestamp 1677622389
transform 1 0 2252 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_143
timestamp 1677622389
transform 1 0 2224 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3472
timestamp 1677622389
transform 1 0 2264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1677622389
transform 1 0 2272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1677622389
transform 1 0 2280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1677622389
transform 1 0 2288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1677622389
transform 1 0 2296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1677622389
transform 1 0 2304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1677622389
transform 1 0 2312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1677622389
transform 1 0 2320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1677622389
transform 1 0 2328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1677622389
transform 1 0 2336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1677622389
transform 1 0 2344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1677622389
transform 1 0 2352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1677622389
transform 1 0 2360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1677622389
transform 1 0 2368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1677622389
transform 1 0 2376 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3083
timestamp 1677622389
transform 1 0 2412 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_145
timestamp 1677622389
transform 1 0 2384 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3496
timestamp 1677622389
transform 1 0 2424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1677622389
transform 1 0 2432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1677622389
transform 1 0 2440 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_255
timestamp 1677622389
transform 1 0 2448 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3510
timestamp 1677622389
transform 1 0 2464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1677622389
transform 1 0 2472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1677622389
transform 1 0 2480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1677622389
transform 1 0 2488 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_155
timestamp 1677622389
transform 1 0 2496 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3514
timestamp 1677622389
transform 1 0 2536 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1677622389
transform 1 0 2544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1677622389
transform 1 0 2552 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_256
timestamp 1677622389
transform 1 0 2560 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3517
timestamp 1677622389
transform 1 0 2576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1677622389
transform 1 0 2584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1677622389
transform 1 0 2592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1677622389
transform 1 0 2600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1677622389
transform 1 0 2608 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_156
timestamp 1677622389
transform 1 0 2616 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3522
timestamp 1677622389
transform 1 0 2656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1677622389
transform 1 0 2664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1677622389
transform 1 0 2672 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_257
timestamp 1677622389
transform 1 0 2680 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3525
timestamp 1677622389
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1677622389
transform 1 0 2704 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1677622389
transform 1 0 2712 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3537
timestamp 1677622389
transform 1 0 2808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1677622389
transform 1 0 2816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1677622389
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1677622389
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1677622389
transform 1 0 2840 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_76
timestamp 1677622389
transform 1 0 2848 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3547
timestamp 1677622389
transform 1 0 2880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1677622389
transform 1 0 2888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1677622389
transform 1 0 2896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1677622389
transform 1 0 2904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1677622389
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1677622389
transform 1 0 2920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1677622389
transform 1 0 2928 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_39
timestamp 1677622389
transform 1 0 2936 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3562
timestamp 1677622389
transform 1 0 2960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1677622389
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1677622389
transform 1 0 2976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1677622389
transform 1 0 2984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1677622389
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_78
timestamp 1677622389
transform -1 0 3032 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3567
timestamp 1677622389
transform 1 0 3032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1677622389
transform 1 0 3040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1677622389
transform 1 0 3048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1677622389
transform 1 0 3056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1677622389
transform 1 0 3064 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_79
timestamp 1677622389
transform -1 0 3104 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3577
timestamp 1677622389
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1677622389
transform 1 0 3112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1677622389
transform 1 0 3120 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_260
timestamp 1677622389
transform -1 0 3144 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3588
timestamp 1677622389
transform 1 0 3144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1677622389
transform 1 0 3152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1677622389
transform 1 0 3160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1677622389
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1677622389
transform 1 0 3176 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_148
timestamp 1677622389
transform -1 0 3224 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3593
timestamp 1677622389
transform 1 0 3224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1677622389
transform 1 0 3232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1677622389
transform 1 0 3240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1677622389
transform 1 0 3248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1677622389
transform 1 0 3256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1677622389
transform 1 0 3264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1677622389
transform 1 0 3272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1677622389
transform 1 0 3280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1677622389
transform 1 0 3288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1677622389
transform 1 0 3296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1677622389
transform 1 0 3304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1677622389
transform 1 0 3312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1677622389
transform 1 0 3320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1677622389
transform 1 0 3328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1677622389
transform 1 0 3336 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_261
timestamp 1677622389
transform -1 0 3360 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3627
timestamp 1677622389
transform 1 0 3360 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1677622389
transform 1 0 3368 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3628
timestamp 1677622389
transform 1 0 3464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1677622389
transform 1 0 3472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1677622389
transform 1 0 3480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1677622389
transform 1 0 3488 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1677622389
transform 1 0 3496 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3632
timestamp 1677622389
transform 1 0 3592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1677622389
transform 1 0 3600 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_263
timestamp 1677622389
transform 1 0 3608 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3636
timestamp 1677622389
transform 1 0 3624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1677622389
transform 1 0 3632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1677622389
transform 1 0 3640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1677622389
transform 1 0 3648 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_149
timestamp 1677622389
transform 1 0 3656 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3644
timestamp 1677622389
transform 1 0 3696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1677622389
transform 1 0 3704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1677622389
transform 1 0 3712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1677622389
transform 1 0 3720 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_150
timestamp 1677622389
transform 1 0 3728 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3652
timestamp 1677622389
transform 1 0 3768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1677622389
transform 1 0 3776 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1677622389
transform 1 0 3784 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_264
timestamp 1677622389
transform 1 0 3880 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3662
timestamp 1677622389
transform 1 0 3896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1677622389
transform 1 0 3904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1677622389
transform 1 0 3912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1677622389
transform 1 0 3920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1677622389
transform 1 0 3928 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1677622389
transform 1 0 3936 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3677
timestamp 1677622389
transform 1 0 4032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1677622389
transform 1 0 4040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1677622389
transform 1 0 4048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1677622389
transform 1 0 4056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1677622389
transform 1 0 4064 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_152
timestamp 1677622389
transform -1 0 4112 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3692
timestamp 1677622389
transform 1 0 4112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1677622389
transform 1 0 4120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1677622389
transform 1 0 4128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1677622389
transform 1 0 4136 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_32
timestamp 1677622389
transform 1 0 4144 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3703
timestamp 1677622389
transform 1 0 4168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1677622389
transform 1 0 4176 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_153
timestamp 1677622389
transform 1 0 4184 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3715
timestamp 1677622389
transform 1 0 4224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1677622389
transform 1 0 4232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1677622389
transform 1 0 4240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1677622389
transform 1 0 4248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1677622389
transform 1 0 4256 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_267
timestamp 1677622389
transform -1 0 4280 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3720
timestamp 1677622389
transform 1 0 4280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1677622389
transform 1 0 4288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1677622389
transform 1 0 4296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1677622389
transform 1 0 4304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1677622389
transform 1 0 4312 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_154
timestamp 1677622389
transform 1 0 4320 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3725
timestamp 1677622389
transform 1 0 4360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1677622389
transform 1 0 4368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1677622389
transform 1 0 4376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1677622389
transform 1 0 4384 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_268
timestamp 1677622389
transform -1 0 4408 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3730
timestamp 1677622389
transform 1 0 4408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1677622389
transform 1 0 4416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1677622389
transform 1 0 4424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1677622389
transform 1 0 4432 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_160
timestamp 1677622389
transform -1 0 4480 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3741
timestamp 1677622389
transform 1 0 4480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1677622389
transform 1 0 4488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1677622389
transform 1 0 4496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1677622389
transform 1 0 4504 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_269
timestamp 1677622389
transform -1 0 4528 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3745
timestamp 1677622389
transform 1 0 4528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1677622389
transform 1 0 4536 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_158
timestamp 1677622389
transform -1 0 4584 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3750
timestamp 1677622389
transform 1 0 4584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1677622389
transform 1 0 4592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1677622389
transform 1 0 4600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1677622389
transform 1 0 4608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1677622389
transform 1 0 4616 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_270
timestamp 1677622389
transform -1 0 4640 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3755
timestamp 1677622389
transform 1 0 4640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1677622389
transform 1 0 4648 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_159
timestamp 1677622389
transform 1 0 4656 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1677622389
transform 1 0 4696 0 -1 3170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_33
timestamp 1677622389
transform 1 0 4843 0 1 3070
box -10 -3 10 3
use M3_M2  M3_M2_3122
timestamp 1677622389
transform 1 0 180 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3494
timestamp 1677622389
transform 1 0 108 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1677622389
transform 1 0 164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1677622389
transform 1 0 172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1677622389
transform 1 0 84 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3185
timestamp 1677622389
transform 1 0 124 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3497
timestamp 1677622389
transform 1 0 180 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3168
timestamp 1677622389
transform 1 0 196 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3498
timestamp 1677622389
transform 1 0 204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1677622389
transform 1 0 220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1677622389
transform 1 0 188 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1677622389
transform 1 0 196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1677622389
transform 1 0 212 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3186
timestamp 1677622389
transform 1 0 220 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1677622389
transform 1 0 236 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1677622389
transform 1 0 252 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3590
timestamp 1677622389
transform 1 0 252 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3134
timestamp 1677622389
transform 1 0 292 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3500
timestamp 1677622389
transform 1 0 268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1677622389
transform 1 0 284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1677622389
transform 1 0 292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1677622389
transform 1 0 276 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3187
timestamp 1677622389
transform 1 0 284 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1677622389
transform 1 0 276 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3503
timestamp 1677622389
transform 1 0 364 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3123
timestamp 1677622389
transform 1 0 404 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1677622389
transform 1 0 412 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3504
timestamp 1677622389
transform 1 0 404 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1677622389
transform 1 0 412 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1677622389
transform 1 0 420 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3136
timestamp 1677622389
transform 1 0 460 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3505
timestamp 1677622389
transform 1 0 444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1677622389
transform 1 0 460 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1677622389
transform 1 0 468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1677622389
transform 1 0 484 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3137
timestamp 1677622389
transform 1 0 516 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3507
timestamp 1677622389
transform 1 0 516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1677622389
transform 1 0 540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1677622389
transform 1 0 524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1677622389
transform 1 0 532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1677622389
transform 1 0 548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1677622389
transform 1 0 564 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3138
timestamp 1677622389
transform 1 0 580 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3599
timestamp 1677622389
transform 1 0 596 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3139
timestamp 1677622389
transform 1 0 636 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3510
timestamp 1677622389
transform 1 0 636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1677622389
transform 1 0 652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1677622389
transform 1 0 644 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3140
timestamp 1677622389
transform 1 0 676 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3601
timestamp 1677622389
transform 1 0 668 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3108
timestamp 1677622389
transform 1 0 732 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3512
timestamp 1677622389
transform 1 0 748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1677622389
transform 1 0 796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1677622389
transform 1 0 716 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3109
timestamp 1677622389
transform 1 0 828 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1677622389
transform 1 0 900 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3514
timestamp 1677622389
transform 1 0 900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1677622389
transform 1 0 916 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3200
timestamp 1677622389
transform 1 0 900 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1677622389
transform 1 0 932 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3603
timestamp 1677622389
transform 1 0 924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1677622389
transform 1 0 932 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3201
timestamp 1677622389
transform 1 0 924 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1677622389
transform 1 0 948 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1677622389
transform 1 0 972 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1677622389
transform 1 0 964 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3491
timestamp 1677622389
transform 1 0 972 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3095
timestamp 1677622389
transform 1 0 1004 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1677622389
transform 1 0 996 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3516
timestamp 1677622389
transform 1 0 996 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1677622389
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1677622389
transform 1 0 1028 0 1 3055
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1677622389
transform 1 0 1028 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3230
timestamp 1677622389
transform 1 0 1028 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3490
timestamp 1677622389
transform 1 0 1044 0 1 3055
box -2 -2 2 2
use M3_M2  M3_M2_3111
timestamp 1677622389
transform 1 0 1052 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1677622389
transform 1 0 1076 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3605
timestamp 1677622389
transform 1 0 1076 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1677622389
transform 1 0 1100 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1677622389
transform 1 0 1116 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3231
timestamp 1677622389
transform 1 0 1124 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1677622389
transform 1 0 1156 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1677622389
transform 1 0 1180 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3518
timestamp 1677622389
transform 1 0 1156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1677622389
transform 1 0 1164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1677622389
transform 1 0 1148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1677622389
transform 1 0 1148 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1677622389
transform 1 0 1180 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3203
timestamp 1677622389
transform 1 0 1164 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1677622389
transform 1 0 1164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1677622389
transform 1 0 1196 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3492
timestamp 1677622389
transform 1 0 1244 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3085
timestamp 1677622389
transform 1 0 1300 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3520
timestamp 1677622389
transform 1 0 1292 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3233
timestamp 1677622389
transform 1 0 1300 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1677622389
transform 1 0 1316 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3609
timestamp 1677622389
transform 1 0 1316 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3086
timestamp 1677622389
transform 1 0 1396 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1677622389
transform 1 0 1332 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1677622389
transform 1 0 1404 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1677622389
transform 1 0 1380 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3521
timestamp 1677622389
transform 1 0 1380 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1677622389
transform 1 0 1332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1677622389
transform 1 0 1444 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3234
timestamp 1677622389
transform 1 0 1444 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1677622389
transform 1 0 1524 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3523
timestamp 1677622389
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1677622389
transform 1 0 1540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1677622389
transform 1 0 1508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1677622389
transform 1 0 1524 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3235
timestamp 1677622389
transform 1 0 1516 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3525
timestamp 1677622389
transform 1 0 1556 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3205
timestamp 1677622389
transform 1 0 1564 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3613
timestamp 1677622389
transform 1 0 1596 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3099
timestamp 1677622389
transform 1 0 1620 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1677622389
transform 1 0 1668 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1677622389
transform 1 0 1692 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1677622389
transform 1 0 1684 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3526
timestamp 1677622389
transform 1 0 1668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1677622389
transform 1 0 1620 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3206
timestamp 1677622389
transform 1 0 1620 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1677622389
transform 1 0 1668 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1677622389
transform 1 0 1724 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1677622389
transform 1 0 1748 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3527
timestamp 1677622389
transform 1 0 1748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1677622389
transform 1 0 1756 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3147
timestamp 1677622389
transform 1 0 1780 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1677622389
transform 1 0 1780 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3615
timestamp 1677622389
transform 1 0 1780 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3188
timestamp 1677622389
transform 1 0 1788 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1677622389
transform 1 0 1788 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1677622389
transform 1 0 1828 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3529
timestamp 1677622389
transform 1 0 1844 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3149
timestamp 1677622389
transform 1 0 1900 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3530
timestamp 1677622389
transform 1 0 1900 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3189
timestamp 1677622389
transform 1 0 1908 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1677622389
transform 1 0 1948 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1677622389
transform 1 0 1988 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3531
timestamp 1677622389
transform 1 0 1948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1677622389
transform 1 0 2004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1677622389
transform 1 0 1924 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3238
timestamp 1677622389
transform 1 0 1972 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3533
timestamp 1677622389
transform 1 0 2060 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1677622389
transform 1 0 2076 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3171
timestamp 1677622389
transform 1 0 2084 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3617
timestamp 1677622389
transform 1 0 2052 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3190
timestamp 1677622389
transform 1 0 2060 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3618
timestamp 1677622389
transform 1 0 2068 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3208
timestamp 1677622389
transform 1 0 2068 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1677622389
transform 1 0 2076 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1677622389
transform 1 0 2092 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3619
timestamp 1677622389
transform 1 0 2100 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1677622389
transform 1 0 2092 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1677622389
transform 1 0 2100 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1677622389
transform 1 0 2116 0 1 2985
box -2 -2 2 2
use M3_M2  M3_M2_3102
timestamp 1677622389
transform 1 0 2164 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1677622389
transform 1 0 2156 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1677622389
transform 1 0 2188 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3535
timestamp 1677622389
transform 1 0 2156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1677622389
transform 1 0 2172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1677622389
transform 1 0 2156 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1677622389
transform 1 0 2148 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3240
timestamp 1677622389
transform 1 0 2140 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1677622389
transform 1 0 2172 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3621
timestamp 1677622389
transform 1 0 2188 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3241
timestamp 1677622389
transform 1 0 2196 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3537
timestamp 1677622389
transform 1 0 2220 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3193
timestamp 1677622389
transform 1 0 2220 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3622
timestamp 1677622389
transform 1 0 2228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1677622389
transform 1 0 2228 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3087
timestamp 1677622389
transform 1 0 2268 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3538
timestamp 1677622389
transform 1 0 2268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1677622389
transform 1 0 2284 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3088
timestamp 1677622389
transform 1 0 2316 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1677622389
transform 1 0 2324 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3539
timestamp 1677622389
transform 1 0 2324 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1677622389
transform 1 0 2316 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3242
timestamp 1677622389
transform 1 0 2308 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1677622389
transform 1 0 2356 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3540
timestamp 1677622389
transform 1 0 2380 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1677622389
transform 1 0 2388 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3194
timestamp 1677622389
transform 1 0 2380 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1677622389
transform 1 0 2396 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1677622389
transform 1 0 2412 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1677622389
transform 1 0 2468 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1677622389
transform 1 0 2420 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3542
timestamp 1677622389
transform 1 0 2460 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3196
timestamp 1677622389
transform 1 0 2420 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3624
timestamp 1677622389
transform 1 0 2484 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3243
timestamp 1677622389
transform 1 0 2484 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3543
timestamp 1677622389
transform 1 0 2540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1677622389
transform 1 0 2508 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3244
timestamp 1677622389
transform 1 0 2524 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3544
timestamp 1677622389
transform 1 0 2604 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3117
timestamp 1677622389
transform 1 0 2644 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1677622389
transform 1 0 2620 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3545
timestamp 1677622389
transform 1 0 2620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1677622389
transform 1 0 2636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1677622389
transform 1 0 2660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1677622389
transform 1 0 2628 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1677622389
transform 1 0 2644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1677622389
transform 1 0 2652 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3245
timestamp 1677622389
transform 1 0 2652 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1677622389
transform 1 0 2668 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1677622389
transform 1 0 2700 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3548
timestamp 1677622389
transform 1 0 2700 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3118
timestamp 1677622389
transform 1 0 2796 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1677622389
transform 1 0 2740 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3549
timestamp 1677622389
transform 1 0 2740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1677622389
transform 1 0 2796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1677622389
transform 1 0 2716 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3247
timestamp 1677622389
transform 1 0 2732 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1677622389
transform 1 0 2828 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3672
timestamp 1677622389
transform 1 0 2828 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1677622389
transform 1 0 2844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1677622389
transform 1 0 2844 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3248
timestamp 1677622389
transform 1 0 2844 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1677622389
transform 1 0 2860 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3552
timestamp 1677622389
transform 1 0 2868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1677622389
transform 1 0 2860 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3209
timestamp 1677622389
transform 1 0 2876 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3632
timestamp 1677622389
transform 1 0 2956 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3091
timestamp 1677622389
transform 1 0 2980 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3493
timestamp 1677622389
transform 1 0 2988 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1677622389
transform 1 0 3036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1677622389
transform 1 0 3140 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3173
timestamp 1677622389
transform 1 0 3220 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3634
timestamp 1677622389
transform 1 0 3228 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3104
timestamp 1677622389
transform 1 0 3252 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3635
timestamp 1677622389
transform 1 0 3268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1677622389
transform 1 0 3284 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3174
timestamp 1677622389
transform 1 0 3292 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3555
timestamp 1677622389
transform 1 0 3300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1677622389
transform 1 0 3292 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1677622389
transform 1 0 3308 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3210
timestamp 1677622389
transform 1 0 3292 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1677622389
transform 1 0 3380 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1677622389
transform 1 0 3340 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1677622389
transform 1 0 3372 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1677622389
transform 1 0 3340 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3556
timestamp 1677622389
transform 1 0 3364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1677622389
transform 1 0 3420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1677622389
transform 1 0 3340 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3211
timestamp 1677622389
transform 1 0 3364 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1677622389
transform 1 0 3436 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1677622389
transform 1 0 3508 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1677622389
transform 1 0 3476 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1677622389
transform 1 0 3492 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3558
timestamp 1677622389
transform 1 0 3476 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1677622389
transform 1 0 3492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1677622389
transform 1 0 3508 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1677622389
transform 1 0 3524 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1677622389
transform 1 0 3460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1677622389
transform 1 0 3468 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3197
timestamp 1677622389
transform 1 0 3476 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3641
timestamp 1677622389
transform 1 0 3492 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1677622389
transform 1 0 3500 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1677622389
transform 1 0 3516 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3198
timestamp 1677622389
transform 1 0 3524 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3562
timestamp 1677622389
transform 1 0 3540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1677622389
transform 1 0 3532 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3212
timestamp 1677622389
transform 1 0 3492 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1677622389
transform 1 0 3540 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1677622389
transform 1 0 3556 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3645
timestamp 1677622389
transform 1 0 3556 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3176
timestamp 1677622389
transform 1 0 3644 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3563
timestamp 1677622389
transform 1 0 3652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1677622389
transform 1 0 3668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1677622389
transform 1 0 3644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1677622389
transform 1 0 3660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1677622389
transform 1 0 3676 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3214
timestamp 1677622389
transform 1 0 3660 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1677622389
transform 1 0 3692 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1677622389
transform 1 0 3756 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1677622389
transform 1 0 3780 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1677622389
transform 1 0 3788 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3565
timestamp 1677622389
transform 1 0 3708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1677622389
transform 1 0 3740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1677622389
transform 1 0 3788 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3215
timestamp 1677622389
transform 1 0 3740 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1677622389
transform 1 0 3788 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1677622389
transform 1 0 3836 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1677622389
transform 1 0 3852 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1677622389
transform 1 0 3908 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1677622389
transform 1 0 3948 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3567
timestamp 1677622389
transform 1 0 3932 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3178
timestamp 1677622389
transform 1 0 3980 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3650
timestamp 1677622389
transform 1 0 3908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3199
timestamp 1677622389
transform 1 0 3940 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3568
timestamp 1677622389
transform 1 0 4012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1677622389
transform 1 0 4020 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3249
timestamp 1677622389
transform 1 0 4004 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3651
timestamp 1677622389
transform 1 0 4028 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3218
timestamp 1677622389
transform 1 0 4020 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1677622389
transform 1 0 4052 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1677622389
transform 1 0 4076 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1677622389
transform 1 0 4108 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3570
timestamp 1677622389
transform 1 0 4100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1677622389
transform 1 0 4116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1677622389
transform 1 0 4132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1677622389
transform 1 0 4108 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1677622389
transform 1 0 4124 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3219
timestamp 1677622389
transform 1 0 4124 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3573
timestamp 1677622389
transform 1 0 4172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1677622389
transform 1 0 4164 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3220
timestamp 1677622389
transform 1 0 4164 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1677622389
transform 1 0 4196 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1677622389
transform 1 0 4204 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1677622389
transform 1 0 4220 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3574
timestamp 1677622389
transform 1 0 4204 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3180
timestamp 1677622389
transform 1 0 4212 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3655
timestamp 1677622389
transform 1 0 4196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1677622389
transform 1 0 4212 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3221
timestamp 1677622389
transform 1 0 4196 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1677622389
transform 1 0 4228 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1677622389
transform 1 0 4228 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1677622389
transform 1 0 4252 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1677622389
transform 1 0 4340 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1677622389
transform 1 0 4268 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3575
timestamp 1677622389
transform 1 0 4292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1677622389
transform 1 0 4348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1677622389
transform 1 0 4268 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3222
timestamp 1677622389
transform 1 0 4292 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1677622389
transform 1 0 4332 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1677622389
transform 1 0 4284 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1677622389
transform 1 0 4332 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1677622389
transform 1 0 4396 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1677622389
transform 1 0 4372 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3577
timestamp 1677622389
transform 1 0 4396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1677622389
transform 1 0 4452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1677622389
transform 1 0 4372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3224
timestamp 1677622389
transform 1 0 4388 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1677622389
transform 1 0 4468 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1677622389
transform 1 0 4460 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1677622389
transform 1 0 4484 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1677622389
transform 1 0 4500 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3579
timestamp 1677622389
transform 1 0 4548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1677622389
transform 1 0 4580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1677622389
transform 1 0 4500 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3226
timestamp 1677622389
transform 1 0 4500 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1677622389
transform 1 0 4620 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3660
timestamp 1677622389
transform 1 0 4612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1677622389
transform 1 0 4628 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3166
timestamp 1677622389
transform 1 0 4676 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3582
timestamp 1677622389
transform 1 0 4652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1677622389
transform 1 0 4668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1677622389
transform 1 0 4644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1677622389
transform 1 0 4660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1677622389
transform 1 0 4692 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3227
timestamp 1677622389
transform 1 0 4684 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1677622389
transform 1 0 4868 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1677622389
transform 1 0 4732 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3584
timestamp 1677622389
transform 1 0 4732 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1677622389
transform 1 0 4788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1677622389
transform 1 0 4708 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3228
timestamp 1677622389
transform 1 0 4708 0 1 2995
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_34
timestamp 1677622389
transform 1 0 48 0 1 2970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_237
timestamp 1677622389
transform 1 0 72 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_272
timestamp 1677622389
transform -1 0 184 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_161
timestamp 1677622389
transform -1 0 224 0 1 2970
box -8 -3 46 105
use FILL  FILL_3767
timestamp 1677622389
transform 1 0 224 0 1 2970
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1677622389
transform 1 0 232 0 1 2970
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1677622389
transform 1 0 240 0 1 2970
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1677622389
transform 1 0 248 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_160
timestamp 1677622389
transform -1 0 296 0 1 2970
box -8 -3 46 105
use FILL  FILL_3785
timestamp 1677622389
transform 1 0 296 0 1 2970
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1677622389
transform 1 0 304 0 1 2970
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1677622389
transform 1 0 312 0 1 2970
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1677622389
transform 1 0 320 0 1 2970
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1677622389
transform 1 0 328 0 1 2970
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1677622389
transform 1 0 336 0 1 2970
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1677622389
transform 1 0 344 0 1 2970
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1677622389
transform 1 0 352 0 1 2970
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1677622389
transform 1 0 360 0 1 2970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1677622389
transform 1 0 368 0 1 2970
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1677622389
transform 1 0 376 0 1 2970
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1677622389
transform 1 0 384 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_274
timestamp 1677622389
transform -1 0 408 0 1 2970
box -9 -3 26 105
use FILL  FILL_3800
timestamp 1677622389
transform 1 0 408 0 1 2970
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1677622389
transform 1 0 416 0 1 2970
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1677622389
transform 1 0 424 0 1 2970
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1677622389
transform 1 0 432 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_163
timestamp 1677622389
transform -1 0 480 0 1 2970
box -8 -3 46 105
use FILL  FILL_3806
timestamp 1677622389
transform 1 0 480 0 1 2970
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1677622389
transform 1 0 488 0 1 2970
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1677622389
transform 1 0 496 0 1 2970
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1677622389
transform 1 0 504 0 1 2970
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1677622389
transform 1 0 512 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_165
timestamp 1677622389
transform 1 0 520 0 1 2970
box -8 -3 46 105
use FILL  FILL_3817
timestamp 1677622389
transform 1 0 560 0 1 2970
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1677622389
transform 1 0 568 0 1 2970
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1677622389
transform 1 0 576 0 1 2970
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1677622389
transform 1 0 584 0 1 2970
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1677622389
transform 1 0 592 0 1 2970
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1677622389
transform 1 0 600 0 1 2970
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1677622389
transform 1 0 608 0 1 2970
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1677622389
transform 1 0 616 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3254
timestamp 1677622389
transform 1 0 644 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_162
timestamp 1677622389
transform -1 0 664 0 1 2970
box -8 -3 46 105
use FILL  FILL_3832
timestamp 1677622389
transform 1 0 664 0 1 2970
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1677622389
transform 1 0 672 0 1 2970
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1677622389
transform 1 0 680 0 1 2970
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1677622389
transform 1 0 688 0 1 2970
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1677622389
transform 1 0 696 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3255
timestamp 1677622389
transform 1 0 756 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_239
timestamp 1677622389
transform 1 0 704 0 1 2970
box -8 -3 104 105
use FILL  FILL_3837
timestamp 1677622389
transform 1 0 800 0 1 2970
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1677622389
transform 1 0 808 0 1 2970
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1677622389
transform 1 0 816 0 1 2970
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1677622389
transform 1 0 824 0 1 2970
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1677622389
transform 1 0 832 0 1 2970
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1677622389
transform 1 0 840 0 1 2970
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1677622389
transform 1 0 848 0 1 2970
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1677622389
transform 1 0 856 0 1 2970
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1677622389
transform 1 0 864 0 1 2970
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1677622389
transform 1 0 872 0 1 2970
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1677622389
transform 1 0 880 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3256
timestamp 1677622389
transform 1 0 900 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1677622389
transform 1 0 916 0 1 2975
box -3 -3 3 3
use OAI21X1  OAI21X1_80
timestamp 1677622389
transform 1 0 888 0 1 2970
box -8 -3 34 105
use FILL  FILL_3866
timestamp 1677622389
transform 1 0 920 0 1 2970
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1677622389
transform 1 0 928 0 1 2970
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1677622389
transform 1 0 936 0 1 2970
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1677622389
transform 1 0 944 0 1 2970
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1677622389
transform 1 0 952 0 1 2970
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1677622389
transform 1 0 960 0 1 2970
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1677622389
transform 1 0 968 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_166
timestamp 1677622389
transform 1 0 976 0 1 2970
box -8 -3 46 105
use FILL  FILL_3880
timestamp 1677622389
transform 1 0 1016 0 1 2970
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1677622389
transform 1 0 1024 0 1 2970
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1677622389
transform 1 0 1032 0 1 2970
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1677622389
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1677622389
transform 1 0 1048 0 1 2970
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1677622389
transform 1 0 1056 0 1 2970
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1677622389
transform 1 0 1064 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_41
timestamp 1677622389
transform 1 0 1072 0 1 2970
box -8 -3 32 105
use FILL  FILL_3899
timestamp 1677622389
transform 1 0 1096 0 1 2970
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1677622389
transform 1 0 1104 0 1 2970
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1677622389
transform 1 0 1112 0 1 2970
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1677622389
transform 1 0 1120 0 1 2970
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1677622389
transform 1 0 1128 0 1 2970
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1677622389
transform 1 0 1136 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3258
timestamp 1677622389
transform 1 0 1156 0 1 2975
box -3 -3 3 3
use FILL  FILL_3912
timestamp 1677622389
transform 1 0 1144 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_82
timestamp 1677622389
transform 1 0 1152 0 1 2970
box -8 -3 34 105
use FILL  FILL_3913
timestamp 1677622389
transform 1 0 1184 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3259
timestamp 1677622389
transform 1 0 1204 0 1 2975
box -3 -3 3 3
use FILL  FILL_3919
timestamp 1677622389
transform 1 0 1192 0 1 2970
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1677622389
transform 1 0 1200 0 1 2970
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1677622389
transform 1 0 1208 0 1 2970
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1677622389
transform 1 0 1216 0 1 2970
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1677622389
transform 1 0 1224 0 1 2970
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1677622389
transform 1 0 1232 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_84
timestamp 1677622389
transform -1 0 1272 0 1 2970
box -8 -3 34 105
use FILL  FILL_3926
timestamp 1677622389
transform 1 0 1272 0 1 2970
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1677622389
transform 1 0 1280 0 1 2970
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1677622389
transform 1 0 1288 0 1 2970
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1677622389
transform 1 0 1296 0 1 2970
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1677622389
transform 1 0 1304 0 1 2970
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1677622389
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1677622389
transform 1 0 1320 0 1 2970
box -8 -3 104 105
use FILL  FILL_3939
timestamp 1677622389
transform 1 0 1416 0 1 2970
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1677622389
transform 1 0 1424 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_279
timestamp 1677622389
transform 1 0 1432 0 1 2970
box -9 -3 26 105
use FILL  FILL_3951
timestamp 1677622389
transform 1 0 1448 0 1 2970
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1677622389
transform 1 0 1456 0 1 2970
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1677622389
transform 1 0 1464 0 1 2970
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1677622389
transform 1 0 1472 0 1 2970
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1677622389
transform 1 0 1480 0 1 2970
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1677622389
transform 1 0 1488 0 1 2970
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1677622389
transform 1 0 1496 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_163
timestamp 1677622389
transform -1 0 1544 0 1 2970
box -8 -3 46 105
use FILL  FILL_3964
timestamp 1677622389
transform 1 0 1544 0 1 2970
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1677622389
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1677622389
transform 1 0 1560 0 1 2970
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1677622389
transform 1 0 1568 0 1 2970
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1677622389
transform 1 0 1576 0 1 2970
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1677622389
transform 1 0 1584 0 1 2970
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1677622389
transform 1 0 1592 0 1 2970
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1677622389
transform 1 0 1600 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_242
timestamp 1677622389
transform 1 0 1608 0 1 2970
box -8 -3 104 105
use FILL  FILL_3977
timestamp 1677622389
transform 1 0 1704 0 1 2970
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1677622389
transform 1 0 1712 0 1 2970
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1677622389
transform 1 0 1720 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_281
timestamp 1677622389
transform 1 0 1728 0 1 2970
box -9 -3 26 105
use FILL  FILL_3987
timestamp 1677622389
transform 1 0 1744 0 1 2970
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1677622389
transform 1 0 1752 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_34
timestamp 1677622389
transform 1 0 1760 0 1 2970
box -5 -3 28 105
use FILL  FILL_3992
timestamp 1677622389
transform 1 0 1784 0 1 2970
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1677622389
transform 1 0 1792 0 1 2970
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1677622389
transform 1 0 1800 0 1 2970
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1677622389
transform 1 0 1808 0 1 2970
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1677622389
transform 1 0 1816 0 1 2970
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1677622389
transform 1 0 1824 0 1 2970
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1677622389
transform 1 0 1832 0 1 2970
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1677622389
transform 1 0 1840 0 1 2970
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1677622389
transform 1 0 1848 0 1 2970
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1677622389
transform 1 0 1856 0 1 2970
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1677622389
transform 1 0 1864 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_282
timestamp 1677622389
transform 1 0 1872 0 1 2970
box -9 -3 26 105
use FILL  FILL_4010
timestamp 1677622389
transform 1 0 1888 0 1 2970
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1677622389
transform 1 0 1896 0 1 2970
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1677622389
transform 1 0 1904 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3260
timestamp 1677622389
transform 1 0 1988 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_244
timestamp 1677622389
transform 1 0 1912 0 1 2970
box -8 -3 104 105
use FILL  FILL_4018
timestamp 1677622389
transform 1 0 2008 0 1 2970
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1677622389
transform 1 0 2016 0 1 2970
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1677622389
transform 1 0 2024 0 1 2970
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1677622389
transform 1 0 2032 0 1 2970
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1677622389
transform 1 0 2040 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_166
timestamp 1677622389
transform 1 0 2048 0 1 2970
box -8 -3 46 105
use FILL  FILL_4035
timestamp 1677622389
transform 1 0 2088 0 1 2970
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1677622389
transform 1 0 2096 0 1 2970
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1677622389
transform 1 0 2104 0 1 2970
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1677622389
transform 1 0 2112 0 1 2970
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1677622389
transform 1 0 2120 0 1 2970
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1677622389
transform 1 0 2128 0 1 2970
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1677622389
transform 1 0 2136 0 1 2970
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1677622389
transform 1 0 2144 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_168
timestamp 1677622389
transform 1 0 2152 0 1 2970
box -8 -3 46 105
use FILL  FILL_4053
timestamp 1677622389
transform 1 0 2192 0 1 2970
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1677622389
transform 1 0 2200 0 1 2970
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1677622389
transform 1 0 2208 0 1 2970
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1677622389
transform 1 0 2216 0 1 2970
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1677622389
transform 1 0 2224 0 1 2970
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1677622389
transform 1 0 2232 0 1 2970
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1677622389
transform 1 0 2240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1677622389
transform 1 0 2248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1677622389
transform 1 0 2256 0 1 2970
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1677622389
transform 1 0 2264 0 1 2970
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1677622389
transform 1 0 2272 0 1 2970
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1677622389
transform 1 0 2280 0 1 2970
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1677622389
transform 1 0 2288 0 1 2970
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1677622389
transform 1 0 2296 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3261
timestamp 1677622389
transform 1 0 2316 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1677622389
transform 1 0 2332 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_170
timestamp 1677622389
transform 1 0 2304 0 1 2970
box -8 -3 46 105
use FILL  FILL_4071
timestamp 1677622389
transform 1 0 2344 0 1 2970
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1677622389
transform 1 0 2352 0 1 2970
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1677622389
transform 1 0 2360 0 1 2970
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1677622389
transform 1 0 2368 0 1 2970
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1677622389
transform 1 0 2376 0 1 2970
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1677622389
transform 1 0 2384 0 1 2970
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1677622389
transform 1 0 2392 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1677622389
transform -1 0 2496 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_247
timestamp 1677622389
transform 1 0 2496 0 1 2970
box -8 -3 104 105
use FILL  FILL_4083
timestamp 1677622389
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1677622389
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1677622389
transform 1 0 2608 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_172
timestamp 1677622389
transform 1 0 2616 0 1 2970
box -8 -3 46 105
use FILL  FILL_4086
timestamp 1677622389
transform 1 0 2656 0 1 2970
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1677622389
transform 1 0 2664 0 1 2970
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1677622389
transform 1 0 2672 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_284
timestamp 1677622389
transform 1 0 2680 0 1 2970
box -9 -3 26 105
use FILL  FILL_4089
timestamp 1677622389
transform 1 0 2696 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3263
timestamp 1677622389
transform 1 0 2732 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_249
timestamp 1677622389
transform 1 0 2704 0 1 2970
box -8 -3 104 105
use FILL  FILL_4103
timestamp 1677622389
transform 1 0 2800 0 1 2970
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1677622389
transform 1 0 2808 0 1 2970
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1677622389
transform 1 0 2816 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_43
timestamp 1677622389
transform 1 0 2824 0 1 2970
box -8 -3 32 105
use FILL  FILL_4109
timestamp 1677622389
transform 1 0 2848 0 1 2970
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1677622389
transform 1 0 2856 0 1 2970
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1677622389
transform 1 0 2864 0 1 2970
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1677622389
transform 1 0 2872 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_88
timestamp 1677622389
transform 1 0 2880 0 1 2970
box -8 -3 34 105
use FILL  FILL_4116
timestamp 1677622389
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1677622389
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1677622389
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1677622389
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1677622389
transform 1 0 2944 0 1 2970
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1677622389
transform 1 0 2952 0 1 2970
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1677622389
transform 1 0 2960 0 1 2970
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1677622389
transform 1 0 2968 0 1 2970
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1677622389
transform 1 0 2976 0 1 2970
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1677622389
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1677622389
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1677622389
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1677622389
transform 1 0 3008 0 1 2970
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1677622389
transform 1 0 3016 0 1 2970
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1677622389
transform 1 0 3024 0 1 2970
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1677622389
transform 1 0 3032 0 1 2970
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1677622389
transform 1 0 3040 0 1 2970
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1677622389
transform 1 0 3048 0 1 2970
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1677622389
transform 1 0 3056 0 1 2970
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1677622389
transform 1 0 3064 0 1 2970
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1677622389
transform 1 0 3072 0 1 2970
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1677622389
transform 1 0 3080 0 1 2970
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1677622389
transform 1 0 3088 0 1 2970
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1677622389
transform 1 0 3096 0 1 2970
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1677622389
transform 1 0 3104 0 1 2970
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1677622389
transform 1 0 3112 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_287
timestamp 1677622389
transform -1 0 3136 0 1 2970
box -9 -3 26 105
use FILL  FILL_4159
timestamp 1677622389
transform 1 0 3136 0 1 2970
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1677622389
transform 1 0 3144 0 1 2970
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1677622389
transform 1 0 3152 0 1 2970
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1677622389
transform 1 0 3160 0 1 2970
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1677622389
transform 1 0 3168 0 1 2970
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1677622389
transform 1 0 3176 0 1 2970
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1677622389
transform 1 0 3184 0 1 2970
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1677622389
transform 1 0 3192 0 1 2970
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1677622389
transform 1 0 3200 0 1 2970
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1677622389
transform 1 0 3208 0 1 2970
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1677622389
transform 1 0 3216 0 1 2970
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1677622389
transform 1 0 3224 0 1 2970
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1677622389
transform 1 0 3232 0 1 2970
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1677622389
transform 1 0 3240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1677622389
transform 1 0 3248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1677622389
transform 1 0 3256 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3264
timestamp 1677622389
transform 1 0 3276 0 1 2975
box -3 -3 3 3
use FILL  FILL_4181
timestamp 1677622389
transform 1 0 3264 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_168
timestamp 1677622389
transform -1 0 3312 0 1 2970
box -8 -3 46 105
use FILL  FILL_4182
timestamp 1677622389
transform 1 0 3312 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3265
timestamp 1677622389
transform 1 0 3332 0 1 2975
box -3 -3 3 3
use FILL  FILL_4186
timestamp 1677622389
transform 1 0 3320 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1677622389
transform 1 0 3328 0 1 2970
box -8 -3 104 105
use FILL  FILL_4188
timestamp 1677622389
transform 1 0 3424 0 1 2970
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1677622389
transform 1 0 3432 0 1 2970
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1677622389
transform 1 0 3440 0 1 2970
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1677622389
transform 1 0 3448 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3266
timestamp 1677622389
transform 1 0 3500 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_175
timestamp 1677622389
transform -1 0 3496 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_170
timestamp 1677622389
transform 1 0 3496 0 1 2970
box -8 -3 46 105
use FILL  FILL_4207
timestamp 1677622389
transform 1 0 3536 0 1 2970
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1677622389
transform 1 0 3544 0 1 2970
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1677622389
transform 1 0 3552 0 1 2970
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1677622389
transform 1 0 3560 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3267
timestamp 1677622389
transform 1 0 3580 0 1 2975
box -3 -3 3 3
use FILL  FILL_4221
timestamp 1677622389
transform 1 0 3568 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_288
timestamp 1677622389
transform 1 0 3576 0 1 2970
box -9 -3 26 105
use FILL  FILL_4223
timestamp 1677622389
transform 1 0 3592 0 1 2970
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1677622389
transform 1 0 3600 0 1 2970
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1677622389
transform 1 0 3608 0 1 2970
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1677622389
transform 1 0 3616 0 1 2970
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1677622389
transform 1 0 3624 0 1 2970
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1677622389
transform 1 0 3632 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3268
timestamp 1677622389
transform 1 0 3676 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_172
timestamp 1677622389
transform -1 0 3680 0 1 2970
box -8 -3 46 105
use FILL  FILL_4234
timestamp 1677622389
transform 1 0 3680 0 1 2970
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1677622389
transform 1 0 3688 0 1 2970
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1677622389
transform 1 0 3696 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3269
timestamp 1677622389
transform 1 0 3716 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_253
timestamp 1677622389
transform -1 0 3800 0 1 2970
box -8 -3 104 105
use FILL  FILL_4237
timestamp 1677622389
transform 1 0 3800 0 1 2970
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1677622389
transform 1 0 3808 0 1 2970
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1677622389
transform 1 0 3816 0 1 2970
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1677622389
transform 1 0 3824 0 1 2970
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1677622389
transform 1 0 3832 0 1 2970
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1677622389
transform 1 0 3840 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3270
timestamp 1677622389
transform 1 0 3860 0 1 2975
box -3 -3 3 3
use FILL  FILL_4261
timestamp 1677622389
transform 1 0 3848 0 1 2970
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1677622389
transform 1 0 3856 0 1 2970
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1677622389
transform 1 0 3864 0 1 2970
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1677622389
transform 1 0 3872 0 1 2970
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1677622389
transform 1 0 3880 0 1 2970
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1677622389
transform 1 0 3888 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1677622389
transform 1 0 3896 0 1 2970
box -8 -3 104 105
use FILL  FILL_4271
timestamp 1677622389
transform 1 0 3992 0 1 2970
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1677622389
transform 1 0 4000 0 1 2970
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1677622389
transform 1 0 4008 0 1 2970
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1677622389
transform 1 0 4016 0 1 2970
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1677622389
transform 1 0 4024 0 1 2970
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1677622389
transform 1 0 4032 0 1 2970
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1677622389
transform 1 0 4040 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_292
timestamp 1677622389
transform 1 0 4048 0 1 2970
box -9 -3 26 105
use FILL  FILL_4290
timestamp 1677622389
transform 1 0 4064 0 1 2970
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1677622389
transform 1 0 4072 0 1 2970
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1677622389
transform 1 0 4080 0 1 2970
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1677622389
transform 1 0 4088 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_177
timestamp 1677622389
transform -1 0 4136 0 1 2970
box -8 -3 46 105
use FILL  FILL_4298
timestamp 1677622389
transform 1 0 4136 0 1 2970
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1677622389
transform 1 0 4144 0 1 2970
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1677622389
transform 1 0 4152 0 1 2970
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1677622389
transform 1 0 4160 0 1 2970
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1677622389
transform 1 0 4168 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_175
timestamp 1677622389
transform 1 0 4176 0 1 2970
box -8 -3 46 105
use FILL  FILL_4308
timestamp 1677622389
transform 1 0 4216 0 1 2970
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1677622389
transform 1 0 4224 0 1 2970
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1677622389
transform 1 0 4232 0 1 2970
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1677622389
transform 1 0 4240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1677622389
transform 1 0 4248 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1677622389
transform 1 0 4256 0 1 2970
box -8 -3 104 105
use FILL  FILL_4317
timestamp 1677622389
transform 1 0 4352 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3271
timestamp 1677622389
transform 1 0 4460 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_256
timestamp 1677622389
transform 1 0 4360 0 1 2970
box -8 -3 104 105
use FILL  FILL_4318
timestamp 1677622389
transform 1 0 4456 0 1 2970
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1677622389
transform 1 0 4464 0 1 2970
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1677622389
transform 1 0 4472 0 1 2970
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1677622389
transform 1 0 4480 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1677622389
transform 1 0 4488 0 1 2970
box -8 -3 104 105
use FILL  FILL_4337
timestamp 1677622389
transform 1 0 4584 0 1 2970
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1677622389
transform 1 0 4592 0 1 2970
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1677622389
transform 1 0 4600 0 1 2970
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1677622389
transform 1 0 4608 0 1 2970
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1677622389
transform 1 0 4616 0 1 2970
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1677622389
transform 1 0 4624 0 1 2970
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1677622389
transform 1 0 4632 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_179
timestamp 1677622389
transform 1 0 4640 0 1 2970
box -8 -3 46 105
use FILL  FILL_4356
timestamp 1677622389
transform 1 0 4680 0 1 2970
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1677622389
transform 1 0 4688 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1677622389
transform 1 0 4696 0 1 2970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_35
timestamp 1677622389
transform 1 0 4819 0 1 2970
box -10 -3 10 3
use M2_M1  M2_M1_3682
timestamp 1677622389
transform 1 0 100 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1677622389
transform 1 0 108 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3353
timestamp 1677622389
transform 1 0 100 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1677622389
transform 1 0 164 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3683
timestamp 1677622389
transform 1 0 164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1677622389
transform 1 0 180 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3272
timestamp 1677622389
transform 1 0 212 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1677622389
transform 1 0 220 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3684
timestamp 1677622389
transform 1 0 212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1677622389
transform 1 0 220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1677622389
transform 1 0 204 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3354
timestamp 1677622389
transform 1 0 204 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1677622389
transform 1 0 212 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3775
timestamp 1677622389
transform 1 0 236 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3373
timestamp 1677622389
transform 1 0 244 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1677622389
transform 1 0 236 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1677622389
transform 1 0 268 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3686
timestamp 1677622389
transform 1 0 268 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1677622389
transform 1 0 284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1677622389
transform 1 0 260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1677622389
transform 1 0 276 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3408
timestamp 1677622389
transform 1 0 300 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3688
timestamp 1677622389
transform 1 0 316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1677622389
transform 1 0 364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1677622389
transform 1 0 396 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1677622389
transform 1 0 404 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3355
timestamp 1677622389
transform 1 0 364 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1677622389
transform 1 0 404 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1677622389
transform 1 0 396 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3781
timestamp 1677622389
transform 1 0 444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3273
timestamp 1677622389
transform 1 0 484 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3689
timestamp 1677622389
transform 1 0 460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1677622389
transform 1 0 468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1677622389
transform 1 0 484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1677622389
transform 1 0 476 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3375
timestamp 1677622389
transform 1 0 468 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3692
timestamp 1677622389
transform 1 0 524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1677622389
transform 1 0 516 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3336
timestamp 1677622389
transform 1 0 524 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1677622389
transform 1 0 548 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3693
timestamp 1677622389
transform 1 0 540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1677622389
transform 1 0 572 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3337
timestamp 1677622389
transform 1 0 564 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3784
timestamp 1677622389
transform 1 0 604 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3357
timestamp 1677622389
transform 1 0 604 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1677622389
transform 1 0 596 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1677622389
transform 1 0 668 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3695
timestamp 1677622389
transform 1 0 620 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3322
timestamp 1677622389
transform 1 0 652 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1677622389
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1677622389
transform 1 0 700 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3358
timestamp 1677622389
transform 1 0 644 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1677622389
transform 1 0 700 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1677622389
transform 1 0 732 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3696
timestamp 1677622389
transform 1 0 732 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1677622389
transform 1 0 748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1677622389
transform 1 0 756 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3277
timestamp 1677622389
transform 1 0 804 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1677622389
transform 1 0 820 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3678
timestamp 1677622389
transform 1 0 876 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3360
timestamp 1677622389
transform 1 0 876 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1677622389
transform 1 0 876 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3697
timestamp 1677622389
transform 1 0 900 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3409
timestamp 1677622389
transform 1 0 900 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3788
timestamp 1677622389
transform 1 0 916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1677622389
transform 1 0 924 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3361
timestamp 1677622389
transform 1 0 916 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1677622389
transform 1 0 948 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3679
timestamp 1677622389
transform 1 0 948 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1677622389
transform 1 0 948 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3362
timestamp 1677622389
transform 1 0 948 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3869
timestamp 1677622389
transform 1 0 956 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3398
timestamp 1677622389
transform 1 0 956 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1677622389
transform 1 0 988 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1677622389
transform 1 0 1036 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3699
timestamp 1677622389
transform 1 0 1124 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3379
timestamp 1677622389
transform 1 0 1156 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3700
timestamp 1677622389
transform 1 0 1180 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3296
timestamp 1677622389
transform 1 0 1220 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3790
timestamp 1677622389
transform 1 0 1196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1677622389
transform 1 0 1204 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3363
timestamp 1677622389
transform 1 0 1196 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3701
timestamp 1677622389
transform 1 0 1228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1677622389
transform 1 0 1220 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3380
timestamp 1677622389
transform 1 0 1204 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1677622389
transform 1 0 1228 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3871
timestamp 1677622389
transform 1 0 1252 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3365
timestamp 1677622389
transform 1 0 1260 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1677622389
transform 1 0 1252 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3702
timestamp 1677622389
transform 1 0 1276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1677622389
transform 1 0 1300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1677622389
transform 1 0 1292 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3399
timestamp 1677622389
transform 1 0 1276 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1677622389
transform 1 0 1292 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1677622389
transform 1 0 1316 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1677622389
transform 1 0 1324 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3704
timestamp 1677622389
transform 1 0 1324 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3366
timestamp 1677622389
transform 1 0 1348 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3872
timestamp 1677622389
transform 1 0 1356 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3305
timestamp 1677622389
transform 1 0 1364 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3793
timestamp 1677622389
transform 1 0 1380 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3413
timestamp 1677622389
transform 1 0 1388 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3675
timestamp 1677622389
transform 1 0 1404 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1677622389
transform 1 0 1428 0 1 2955
box -2 -2 2 2
use M3_M2  M3_M2_3306
timestamp 1677622389
transform 1 0 1420 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3705
timestamp 1677622389
transform 1 0 1468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1677622389
transform 1 0 1460 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3367
timestamp 1677622389
transform 1 0 1468 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1677622389
transform 1 0 1460 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3706
timestamp 1677622389
transform 1 0 1508 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3280
timestamp 1677622389
transform 1 0 1540 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3707
timestamp 1677622389
transform 1 0 1540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1677622389
transform 1 0 1532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1677622389
transform 1 0 1556 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3382
timestamp 1677622389
transform 1 0 1532 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1677622389
transform 1 0 1580 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3708
timestamp 1677622389
transform 1 0 1580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1677622389
transform 1 0 1580 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3368
timestamp 1677622389
transform 1 0 1580 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1677622389
transform 1 0 1620 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3709
timestamp 1677622389
transform 1 0 1668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1677622389
transform 1 0 1620 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3369
timestamp 1677622389
transform 1 0 1644 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3799
timestamp 1677622389
transform 1 0 1724 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3323
timestamp 1677622389
transform 1 0 1764 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3710
timestamp 1677622389
transform 1 0 1772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1677622389
transform 1 0 1756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1677622389
transform 1 0 1804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1677622389
transform 1 0 1844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1677622389
transform 1 0 1860 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1677622389
transform 1 0 1852 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3383
timestamp 1677622389
transform 1 0 1844 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3803
timestamp 1677622389
transform 1 0 1876 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3400
timestamp 1677622389
transform 1 0 1876 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3804
timestamp 1677622389
transform 1 0 1908 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3384
timestamp 1677622389
transform 1 0 1908 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3713
timestamp 1677622389
transform 1 0 1940 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3401
timestamp 1677622389
transform 1 0 1932 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1677622389
transform 1 0 1964 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3714
timestamp 1677622389
transform 1 0 1964 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1677622389
transform 1 0 1972 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3385
timestamp 1677622389
transform 1 0 1948 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1677622389
transform 1 0 1988 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1677622389
transform 1 0 1988 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3715
timestamp 1677622389
transform 1 0 2004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1677622389
transform 1 0 2052 0 1 2895
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1677622389
transform 1 0 2084 0 1 2895
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1677622389
transform 1 0 2124 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3283
timestamp 1677622389
transform 1 0 2148 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1677622389
transform 1 0 2164 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1677622389
transform 1 0 2180 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1677622389
transform 1 0 2140 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1677622389
transform 1 0 2164 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3716
timestamp 1677622389
transform 1 0 2140 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1677622389
transform 1 0 2148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1677622389
transform 1 0 2156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1677622389
transform 1 0 2172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1677622389
transform 1 0 2164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1677622389
transform 1 0 2180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1677622389
transform 1 0 2188 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3386
timestamp 1677622389
transform 1 0 2156 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1677622389
transform 1 0 2180 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1677622389
transform 1 0 2204 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1677622389
transform 1 0 2204 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3720
timestamp 1677622389
transform 1 0 2220 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3286
timestamp 1677622389
transform 1 0 2268 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1677622389
transform 1 0 2300 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3721
timestamp 1677622389
transform 1 0 2308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1677622389
transform 1 0 2268 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3404
timestamp 1677622389
transform 1 0 2236 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1677622389
transform 1 0 2236 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1677622389
transform 1 0 2300 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1677622389
transform 1 0 2324 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3722
timestamp 1677622389
transform 1 0 2332 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3387
timestamp 1677622389
transform 1 0 2332 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1677622389
transform 1 0 2372 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3723
timestamp 1677622389
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1677622389
transform 1 0 2348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1677622389
transform 1 0 2364 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3338
timestamp 1677622389
transform 1 0 2372 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3813
timestamp 1677622389
transform 1 0 2380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1677622389
transform 1 0 2404 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3339
timestamp 1677622389
transform 1 0 2404 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1677622389
transform 1 0 2452 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1677622389
transform 1 0 2436 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1677622389
transform 1 0 2476 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3725
timestamp 1677622389
transform 1 0 2524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1677622389
transform 1 0 2436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1677622389
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1677622389
transform 1 0 2476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1677622389
transform 1 0 2540 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3327
timestamp 1677622389
transform 1 0 2572 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1677622389
transform 1 0 2604 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3726
timestamp 1677622389
transform 1 0 2580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1677622389
transform 1 0 2588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1677622389
transform 1 0 2604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1677622389
transform 1 0 2564 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3328
timestamp 1677622389
transform 1 0 2612 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1677622389
transform 1 0 2588 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3819
timestamp 1677622389
transform 1 0 2596 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1677622389
transform 1 0 2612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1677622389
transform 1 0 2620 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3388
timestamp 1677622389
transform 1 0 2612 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3729
timestamp 1677622389
transform 1 0 2628 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3341
timestamp 1677622389
transform 1 0 2628 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1677622389
transform 1 0 2644 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3822
timestamp 1677622389
transform 1 0 2676 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1677622389
transform 1 0 2692 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3390
timestamp 1677622389
transform 1 0 2660 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1677622389
transform 1 0 2692 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1677622389
transform 1 0 2716 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3730
timestamp 1677622389
transform 1 0 2716 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3290
timestamp 1677622389
transform 1 0 2820 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1677622389
transform 1 0 2812 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3731
timestamp 1677622389
transform 1 0 2732 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1677622389
transform 1 0 2820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1677622389
transform 1 0 2756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1677622389
transform 1 0 2812 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3392
timestamp 1677622389
transform 1 0 2732 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3826
timestamp 1677622389
transform 1 0 2836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1677622389
transform 1 0 2844 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3313
timestamp 1677622389
transform 1 0 2868 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3680
timestamp 1677622389
transform 1 0 2876 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3291
timestamp 1677622389
transform 1 0 2900 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1677622389
transform 1 0 2892 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1677622389
transform 1 0 2892 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3873
timestamp 1677622389
transform 1 0 2892 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1677622389
transform 1 0 2908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1677622389
transform 1 0 2932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1677622389
transform 1 0 2924 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3343
timestamp 1677622389
transform 1 0 2932 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1677622389
transform 1 0 2948 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3681
timestamp 1677622389
transform 1 0 2964 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1677622389
transform 1 0 2972 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1677622389
transform 1 0 3012 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3292
timestamp 1677622389
transform 1 0 3060 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1677622389
transform 1 0 3044 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1677622389
transform 1 0 3060 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3735
timestamp 1677622389
transform 1 0 3036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1677622389
transform 1 0 3044 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3344
timestamp 1677622389
transform 1 0 3036 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1677622389
transform 1 0 3052 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3737
timestamp 1677622389
transform 1 0 3060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1677622389
transform 1 0 3052 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3345
timestamp 1677622389
transform 1 0 3060 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3831
timestamp 1677622389
transform 1 0 3068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1677622389
transform 1 0 3084 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3418
timestamp 1677622389
transform 1 0 3108 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1677622389
transform 1 0 3172 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3739
timestamp 1677622389
transform 1 0 3220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1677622389
transform 1 0 3140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1677622389
transform 1 0 3172 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3405
timestamp 1677622389
transform 1 0 3180 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1677622389
transform 1 0 3260 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3740
timestamp 1677622389
transform 1 0 3268 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1677622389
transform 1 0 3284 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3330
timestamp 1677622389
transform 1 0 3300 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3834
timestamp 1677622389
transform 1 0 3276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1677622389
transform 1 0 3300 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3346
timestamp 1677622389
transform 1 0 3308 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1677622389
transform 1 0 3324 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3742
timestamp 1677622389
transform 1 0 3324 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3293
timestamp 1677622389
transform 1 0 3372 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3743
timestamp 1677622389
transform 1 0 3364 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3301
timestamp 1677622389
transform 1 0 3460 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3744
timestamp 1677622389
transform 1 0 3500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1677622389
transform 1 0 3532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1677622389
transform 1 0 3516 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1677622389
transform 1 0 3540 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3394
timestamp 1677622389
transform 1 0 3540 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3746
timestamp 1677622389
transform 1 0 3556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1677622389
transform 1 0 3604 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3395
timestamp 1677622389
transform 1 0 3604 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3747
timestamp 1677622389
transform 1 0 3660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1677622389
transform 1 0 3652 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3419
timestamp 1677622389
transform 1 0 3652 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3748
timestamp 1677622389
transform 1 0 3708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1677622389
transform 1 0 3724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1677622389
transform 1 0 3748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1677622389
transform 1 0 3764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1677622389
transform 1 0 3772 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1677622389
transform 1 0 3828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1677622389
transform 1 0 3836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1677622389
transform 1 0 3860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1677622389
transform 1 0 3852 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1677622389
transform 1 0 3900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1677622389
transform 1 0 3892 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3406
timestamp 1677622389
transform 1 0 3900 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3847
timestamp 1677622389
transform 1 0 3916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1677622389
transform 1 0 3924 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3396
timestamp 1677622389
transform 1 0 3924 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3750
timestamp 1677622389
transform 1 0 3940 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1677622389
transform 1 0 3956 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3331
timestamp 1677622389
transform 1 0 3964 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3848
timestamp 1677622389
transform 1 0 3964 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1677622389
transform 1 0 3980 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3420
timestamp 1677622389
transform 1 0 3980 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3753
timestamp 1677622389
transform 1 0 4012 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3332
timestamp 1677622389
transform 1 0 4020 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3849
timestamp 1677622389
transform 1 0 4020 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3333
timestamp 1677622389
transform 1 0 4068 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3754
timestamp 1677622389
transform 1 0 4076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1677622389
transform 1 0 4108 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3334
timestamp 1677622389
transform 1 0 4116 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3756
timestamp 1677622389
transform 1 0 4132 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1677622389
transform 1 0 4100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1677622389
transform 1 0 4124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1677622389
transform 1 0 4164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1677622389
transform 1 0 4180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1677622389
transform 1 0 4196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1677622389
transform 1 0 4204 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3347
timestamp 1677622389
transform 1 0 4164 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3852
timestamp 1677622389
transform 1 0 4172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1677622389
transform 1 0 4188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1677622389
transform 1 0 4220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1677622389
transform 1 0 4252 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3348
timestamp 1677622389
transform 1 0 4252 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3855
timestamp 1677622389
transform 1 0 4260 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3397
timestamp 1677622389
transform 1 0 4260 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3856
timestamp 1677622389
transform 1 0 4284 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3318
timestamp 1677622389
transform 1 0 4324 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1677622389
transform 1 0 4324 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1677622389
transform 1 0 4340 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1677622389
transform 1 0 4356 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3762
timestamp 1677622389
transform 1 0 4348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1677622389
transform 1 0 4356 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1677622389
transform 1 0 4356 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3335
timestamp 1677622389
transform 1 0 4372 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3764
timestamp 1677622389
transform 1 0 4380 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3302
timestamp 1677622389
transform 1 0 4404 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3765
timestamp 1677622389
transform 1 0 4404 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1677622389
transform 1 0 4372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1677622389
transform 1 0 4388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1677622389
transform 1 0 4396 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3350
timestamp 1677622389
transform 1 0 4404 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1677622389
transform 1 0 4396 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1677622389
transform 1 0 4436 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1677622389
transform 1 0 4452 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3766
timestamp 1677622389
transform 1 0 4452 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1677622389
transform 1 0 4444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1677622389
transform 1 0 4460 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3352
timestamp 1677622389
transform 1 0 4468 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3863
timestamp 1677622389
transform 1 0 4484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1677622389
transform 1 0 4564 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3422
timestamp 1677622389
transform 1 0 4556 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3768
timestamp 1677622389
transform 1 0 4572 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1677622389
transform 1 0 4572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1677622389
transform 1 0 4596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1677622389
transform 1 0 4612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1677622389
transform 1 0 4588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1677622389
transform 1 0 4604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1677622389
transform 1 0 4620 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3371
timestamp 1677622389
transform 1 0 4612 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1677622389
transform 1 0 4588 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1677622389
transform 1 0 4668 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3868
timestamp 1677622389
transform 1 0 4668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1677622389
transform 1 0 4764 0 1 2935
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_36
timestamp 1677622389
transform 1 0 24 0 1 2870
box -10 -3 10 3
use FILL  FILL_3768
timestamp 1677622389
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1677622389
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1677622389
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_273
timestamp 1677622389
transform 1 0 96 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3771
timestamp 1677622389
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1677622389
transform 1 0 120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1677622389
transform 1 0 128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1677622389
transform 1 0 136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1677622389
transform 1 0 144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1677622389
transform 1 0 152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1677622389
transform 1 0 160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1677622389
transform 1 0 168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1677622389
transform 1 0 176 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_162
timestamp 1677622389
transform -1 0 224 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3780
timestamp 1677622389
transform 1 0 224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1677622389
transform 1 0 232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1677622389
transform 1 0 240 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_161
timestamp 1677622389
transform -1 0 288 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3787
timestamp 1677622389
transform 1 0 288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1677622389
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1677622389
transform 1 0 304 0 -1 2970
box -8 -3 104 105
use INVX2  INVX2_275
timestamp 1677622389
transform -1 0 416 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3802
timestamp 1677622389
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1677622389
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1677622389
transform 1 0 432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1677622389
transform 1 0 440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1677622389
transform 1 0 448 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_164
timestamp 1677622389
transform -1 0 496 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3812
timestamp 1677622389
transform 1 0 496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1677622389
transform 1 0 504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1677622389
transform 1 0 512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1677622389
transform 1 0 520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1677622389
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1677622389
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_276
timestamp 1677622389
transform 1 0 544 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3821
timestamp 1677622389
transform 1 0 560 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_277
timestamp 1677622389
transform 1 0 568 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3825
timestamp 1677622389
transform 1 0 584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1677622389
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1677622389
transform 1 0 600 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1677622389
transform 1 0 608 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3838
timestamp 1677622389
transform 1 0 704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1677622389
transform 1 0 712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1677622389
transform 1 0 720 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_278
timestamp 1677622389
transform 1 0 728 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3841
timestamp 1677622389
transform 1 0 744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1677622389
transform 1 0 752 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1677622389
transform 1 0 760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1677622389
transform 1 0 768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1677622389
transform 1 0 776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1677622389
transform 1 0 784 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3424
timestamp 1677622389
transform 1 0 804 0 1 2875
box -3 -3 3 3
use FILL  FILL_3847
timestamp 1677622389
transform 1 0 792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1677622389
transform 1 0 800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1677622389
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1677622389
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_40
timestamp 1677622389
transform 1 0 824 0 -1 2970
box -8 -3 32 105
use FILL  FILL_3857
timestamp 1677622389
transform 1 0 848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1677622389
transform 1 0 856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1677622389
transform 1 0 864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1677622389
transform 1 0 872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1677622389
transform 1 0 880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1677622389
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1677622389
transform 1 0 896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1677622389
transform 1 0 904 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_81
timestamp 1677622389
transform 1 0 912 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3873
timestamp 1677622389
transform 1 0 944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1677622389
transform 1 0 952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1677622389
transform 1 0 960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1677622389
transform 1 0 968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1677622389
transform 1 0 976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1677622389
transform 1 0 984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1677622389
transform 1 0 992 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3425
timestamp 1677622389
transform 1 0 1012 0 1 2875
box -3 -3 3 3
use FILL  FILL_3884
timestamp 1677622389
transform 1 0 1000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1677622389
transform 1 0 1008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1677622389
transform 1 0 1016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1677622389
transform 1 0 1024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1677622389
transform 1 0 1032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1677622389
transform 1 0 1040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1677622389
transform 1 0 1048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1677622389
transform 1 0 1056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1677622389
transform 1 0 1064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1677622389
transform 1 0 1072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1677622389
transform 1 0 1080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1677622389
transform 1 0 1088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1677622389
transform 1 0 1096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1677622389
transform 1 0 1104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1677622389
transform 1 0 1112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1677622389
transform 1 0 1120 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3426
timestamp 1677622389
transform 1 0 1140 0 1 2875
box -3 -3 3 3
use NOR2X1  NOR2X1_42
timestamp 1677622389
transform 1 0 1128 0 -1 2970
box -8 -3 32 105
use FILL  FILL_3914
timestamp 1677622389
transform 1 0 1152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1677622389
transform 1 0 1160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1677622389
transform 1 0 1168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1677622389
transform 1 0 1176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1677622389
transform 1 0 1184 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_83
timestamp 1677622389
transform 1 0 1192 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3924
timestamp 1677622389
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1677622389
transform 1 0 1232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1677622389
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1677622389
transform 1 0 1248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1677622389
transform 1 0 1256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1677622389
transform 1 0 1264 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_85
timestamp 1677622389
transform -1 0 1304 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3936
timestamp 1677622389
transform 1 0 1304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1677622389
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1677622389
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1677622389
transform 1 0 1328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1677622389
transform 1 0 1336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1677622389
transform 1 0 1344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1677622389
transform 1 0 1352 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1677622389
transform -1 0 1392 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3945
timestamp 1677622389
transform 1 0 1392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1677622389
transform 1 0 1400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1677622389
transform 1 0 1408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1677622389
transform 1 0 1416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1677622389
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1677622389
transform 1 0 1432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1677622389
transform 1 0 1440 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_280
timestamp 1677622389
transform -1 0 1464 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3956
timestamp 1677622389
transform 1 0 1464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1677622389
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1677622389
transform 1 0 1480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1677622389
transform 1 0 1488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1677622389
transform 1 0 1496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1677622389
transform 1 0 1504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1677622389
transform 1 0 1512 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_164
timestamp 1677622389
transform -1 0 1560 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3970
timestamp 1677622389
transform 1 0 1560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1677622389
transform 1 0 1568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1677622389
transform 1 0 1576 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1677622389
transform -1 0 1680 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3979
timestamp 1677622389
transform 1 0 1680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1677622389
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1677622389
transform 1 0 1696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1677622389
transform 1 0 1704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1677622389
transform 1 0 1712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1677622389
transform 1 0 1720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1677622389
transform 1 0 1728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1677622389
transform 1 0 1736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1677622389
transform 1 0 1744 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_35
timestamp 1677622389
transform 1 0 1752 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3993
timestamp 1677622389
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1677622389
transform 1 0 1784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1677622389
transform 1 0 1792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1677622389
transform 1 0 1800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1677622389
transform 1 0 1808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1677622389
transform 1 0 1816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1677622389
transform 1 0 1824 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_167
timestamp 1677622389
transform 1 0 1832 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4011
timestamp 1677622389
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1677622389
transform 1 0 1880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1677622389
transform 1 0 1888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1677622389
transform 1 0 1896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1677622389
transform 1 0 1904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1677622389
transform 1 0 1912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1677622389
transform 1 0 1920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1677622389
transform 1 0 1928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1677622389
transform 1 0 1936 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3427
timestamp 1677622389
transform 1 0 1956 0 1 2875
box -3 -3 3 3
use OAI22X1  OAI22X1_165
timestamp 1677622389
transform 1 0 1944 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4023
timestamp 1677622389
transform 1 0 1984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1677622389
transform 1 0 1992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1677622389
transform 1 0 2000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1677622389
transform 1 0 2008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1677622389
transform 1 0 2016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1677622389
transform 1 0 2024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1677622389
transform 1 0 2032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1677622389
transform 1 0 2040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1677622389
transform 1 0 2048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1677622389
transform 1 0 2056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1677622389
transform 1 0 2064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1677622389
transform 1 0 2072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1677622389
transform 1 0 2080 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3428
timestamp 1677622389
transform 1 0 2100 0 1 2875
box -3 -3 3 3
use INVX2  INVX2_283
timestamp 1677622389
transform -1 0 2104 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4043
timestamp 1677622389
transform 1 0 2104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1677622389
transform 1 0 2112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1677622389
transform 1 0 2120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1677622389
transform 1 0 2128 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3429
timestamp 1677622389
transform 1 0 2148 0 1 2875
box -3 -3 3 3
use FILL  FILL_4051
timestamp 1677622389
transform 1 0 2136 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_169
timestamp 1677622389
transform 1 0 2144 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4054
timestamp 1677622389
transform 1 0 2184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1677622389
transform 1 0 2192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1677622389
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1677622389
transform 1 0 2208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1677622389
transform 1 0 2216 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1677622389
transform -1 0 2320 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4078
timestamp 1677622389
transform 1 0 2320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1677622389
transform 1 0 2328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1677622389
transform 1 0 2336 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_171
timestamp 1677622389
transform 1 0 2344 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4081
timestamp 1677622389
transform 1 0 2384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1677622389
transform 1 0 2392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1677622389
transform 1 0 2400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1677622389
transform 1 0 2408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1677622389
transform 1 0 2416 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_285
timestamp 1677622389
transform 1 0 2424 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_248
timestamp 1677622389
transform -1 0 2536 0 -1 2970
box -8 -3 104 105
use INVX2  INVX2_286
timestamp 1677622389
transform -1 0 2552 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4094
timestamp 1677622389
transform 1 0 2552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1677622389
transform 1 0 2560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1677622389
transform 1 0 2568 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_173
timestamp 1677622389
transform 1 0 2576 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4097
timestamp 1677622389
transform 1 0 2616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1677622389
transform 1 0 2624 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1677622389
transform 1 0 2632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1677622389
transform 1 0 2640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1677622389
transform 1 0 2648 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_174
timestamp 1677622389
transform 1 0 2656 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4102
timestamp 1677622389
transform 1 0 2696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1677622389
transform 1 0 2704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1677622389
transform 1 0 2712 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1677622389
transform 1 0 2720 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4108
timestamp 1677622389
transform 1 0 2816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1677622389
transform 1 0 2824 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_87
timestamp 1677622389
transform 1 0 2832 0 -1 2970
box -8 -3 34 105
use FILL  FILL_4113
timestamp 1677622389
transform 1 0 2864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1677622389
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1677622389
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1677622389
transform 1 0 2888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1677622389
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_44
timestamp 1677622389
transform 1 0 2904 0 -1 2970
box -8 -3 32 105
use FILL  FILL_4122
timestamp 1677622389
transform 1 0 2928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1677622389
transform 1 0 2936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1677622389
transform 1 0 2944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1677622389
transform 1 0 2952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1677622389
transform 1 0 2960 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_89
timestamp 1677622389
transform -1 0 3000 0 -1 2970
box -8 -3 34 105
use FILL  FILL_4136
timestamp 1677622389
transform 1 0 3000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1677622389
transform 1 0 3008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1677622389
transform 1 0 3016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1677622389
transform 1 0 3024 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3430
timestamp 1677622389
transform 1 0 3044 0 1 2875
box -3 -3 3 3
use FILL  FILL_4144
timestamp 1677622389
transform 1 0 3032 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_167
timestamp 1677622389
transform 1 0 3040 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4151
timestamp 1677622389
transform 1 0 3080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1677622389
transform 1 0 3088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1677622389
transform 1 0 3096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1677622389
transform 1 0 3104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1677622389
transform 1 0 3112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1677622389
transform 1 0 3120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1677622389
transform 1 0 3128 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1677622389
transform -1 0 3232 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4175
timestamp 1677622389
transform 1 0 3232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1677622389
transform 1 0 3240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1677622389
transform 1 0 3248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1677622389
transform 1 0 3256 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_169
timestamp 1677622389
transform -1 0 3304 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4184
timestamp 1677622389
transform 1 0 3304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1677622389
transform 1 0 3312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1677622389
transform 1 0 3320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1677622389
transform 1 0 3328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1677622389
transform 1 0 3336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1677622389
transform 1 0 3344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1677622389
transform 1 0 3352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1677622389
transform 1 0 3360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1677622389
transform 1 0 3368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1677622389
transform 1 0 3376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1677622389
transform 1 0 3384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1677622389
transform 1 0 3392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1677622389
transform 1 0 3400 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3431
timestamp 1677622389
transform 1 0 3420 0 1 2875
box -3 -3 3 3
use FILL  FILL_4199
timestamp 1677622389
transform 1 0 3408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1677622389
transform 1 0 3416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1677622389
transform 1 0 3424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1677622389
transform 1 0 3432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1677622389
transform 1 0 3440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1677622389
transform 1 0 3448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1677622389
transform 1 0 3456 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3432
timestamp 1677622389
transform 1 0 3476 0 1 2875
box -3 -3 3 3
use FILL  FILL_4212
timestamp 1677622389
transform 1 0 3464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1677622389
transform 1 0 3472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1677622389
transform 1 0 3480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1677622389
transform 1 0 3488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1677622389
transform 1 0 3496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1677622389
transform 1 0 3504 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_171
timestamp 1677622389
transform 1 0 3512 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4218
timestamp 1677622389
transform 1 0 3552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1677622389
transform 1 0 3560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1677622389
transform 1 0 3568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1677622389
transform 1 0 3576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1677622389
transform 1 0 3584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1677622389
transform 1 0 3592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1677622389
transform 1 0 3600 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_289
timestamp 1677622389
transform -1 0 3624 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4232
timestamp 1677622389
transform 1 0 3624 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1677622389
transform 1 0 3632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1677622389
transform 1 0 3640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1677622389
transform 1 0 3648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1677622389
transform 1 0 3656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1677622389
transform 1 0 3664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1677622389
transform 1 0 3672 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_290
timestamp 1677622389
transform -1 0 3696 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4244
timestamp 1677622389
transform 1 0 3696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1677622389
transform 1 0 3704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1677622389
transform 1 0 3712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1677622389
transform 1 0 3720 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3433
timestamp 1677622389
transform 1 0 3748 0 1 2875
box -3 -3 3 3
use AOI22X1  AOI22X1_176
timestamp 1677622389
transform 1 0 3728 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4248
timestamp 1677622389
transform 1 0 3768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1677622389
transform 1 0 3776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1677622389
transform 1 0 3784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1677622389
transform 1 0 3792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1677622389
transform 1 0 3800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1677622389
transform 1 0 3808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1677622389
transform 1 0 3816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1677622389
transform 1 0 3824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1677622389
transform 1 0 3832 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_22
timestamp 1677622389
transform -1 0 3872 0 -1 2970
box -8 -3 40 105
use FILL  FILL_4266
timestamp 1677622389
transform 1 0 3872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1677622389
transform 1 0 3880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1677622389
transform 1 0 3888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1677622389
transform 1 0 3896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1677622389
transform 1 0 3904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1677622389
transform 1 0 3912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1677622389
transform 1 0 3920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1677622389
transform 1 0 3928 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_173
timestamp 1677622389
transform 1 0 3936 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4277
timestamp 1677622389
transform 1 0 3976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1677622389
transform 1 0 3984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1677622389
transform 1 0 3992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1677622389
transform 1 0 4000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1677622389
transform 1 0 4008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1677622389
transform 1 0 4016 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_291
timestamp 1677622389
transform 1 0 4024 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4289
timestamp 1677622389
transform 1 0 4040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1677622389
transform 1 0 4048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1677622389
transform 1 0 4056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1677622389
transform 1 0 4064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1677622389
transform 1 0 4072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1677622389
transform 1 0 4080 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_174
timestamp 1677622389
transform -1 0 4128 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4300
timestamp 1677622389
transform 1 0 4128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1677622389
transform 1 0 4136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1677622389
transform 1 0 4144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1677622389
transform 1 0 4152 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3434
timestamp 1677622389
transform 1 0 4196 0 1 2875
box -3 -3 3 3
use OAI22X1  OAI22X1_176
timestamp 1677622389
transform 1 0 4160 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4309
timestamp 1677622389
transform 1 0 4200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1677622389
transform 1 0 4208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1677622389
transform 1 0 4216 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3435
timestamp 1677622389
transform 1 0 4236 0 1 2875
box -3 -3 3 3
use FILL  FILL_4313
timestamp 1677622389
transform 1 0 4224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1677622389
transform 1 0 4232 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_178
timestamp 1677622389
transform -1 0 4280 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4323
timestamp 1677622389
transform 1 0 4280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1677622389
transform 1 0 4288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1677622389
transform 1 0 4296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1677622389
transform 1 0 4304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1677622389
transform 1 0 4312 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_293
timestamp 1677622389
transform -1 0 4336 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4328
timestamp 1677622389
transform 1 0 4336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1677622389
transform 1 0 4344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1677622389
transform 1 0 4352 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_177
timestamp 1677622389
transform -1 0 4400 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4331
timestamp 1677622389
transform 1 0 4400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1677622389
transform 1 0 4408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1677622389
transform 1 0 4416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1677622389
transform 1 0 4424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1677622389
transform 1 0 4432 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_179
timestamp 1677622389
transform -1 0 4480 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4336
timestamp 1677622389
transform 1 0 4480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1677622389
transform 1 0 4488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1677622389
transform 1 0 4496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1677622389
transform 1 0 4504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1677622389
transform 1 0 4512 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_294
timestamp 1677622389
transform -1 0 4536 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4346
timestamp 1677622389
transform 1 0 4536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1677622389
transform 1 0 4544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1677622389
transform 1 0 4552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1677622389
transform 1 0 4560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1677622389
transform 1 0 4568 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_178
timestamp 1677622389
transform -1 0 4616 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4351
timestamp 1677622389
transform 1 0 4616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1677622389
transform 1 0 4624 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1677622389
transform 1 0 4632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1677622389
transform 1 0 4640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1677622389
transform 1 0 4648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1677622389
transform 1 0 4656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1677622389
transform 1 0 4664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1677622389
transform 1 0 4672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1677622389
transform 1 0 4680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1677622389
transform 1 0 4688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1677622389
transform 1 0 4696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1677622389
transform 1 0 4704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1677622389
transform 1 0 4712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1677622389
transform 1 0 4720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1677622389
transform 1 0 4728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1677622389
transform 1 0 4736 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_295
timestamp 1677622389
transform -1 0 4760 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4371
timestamp 1677622389
transform 1 0 4760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1677622389
transform 1 0 4768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1677622389
transform 1 0 4776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1677622389
transform 1 0 4784 0 -1 2970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_37
timestamp 1677622389
transform 1 0 4843 0 1 2870
box -10 -3 10 3
use M3_M2  M3_M2_3488
timestamp 1677622389
transform 1 0 156 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3893
timestamp 1677622389
transform 1 0 156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1677622389
transform 1 0 156 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3554
timestamp 1677622389
transform 1 0 156 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1677622389
transform 1 0 196 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3894
timestamp 1677622389
transform 1 0 196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1677622389
transform 1 0 172 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3462
timestamp 1677622389
transform 1 0 300 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3895
timestamp 1677622389
transform 1 0 268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1677622389
transform 1 0 284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1677622389
transform 1 0 300 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3530
timestamp 1677622389
transform 1 0 268 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3987
timestamp 1677622389
transform 1 0 276 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3555
timestamp 1677622389
transform 1 0 284 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3988
timestamp 1677622389
transform 1 0 332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1677622389
transform 1 0 388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1677622389
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1677622389
transform 1 0 356 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3556
timestamp 1677622389
transform 1 0 356 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1677622389
transform 1 0 396 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1677622389
transform 1 0 444 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1677622389
transform 1 0 492 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1677622389
transform 1 0 492 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3900
timestamp 1677622389
transform 1 0 516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1677622389
transform 1 0 548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1677622389
transform 1 0 468 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3558
timestamp 1677622389
transform 1 0 468 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3902
timestamp 1677622389
transform 1 0 564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1677622389
transform 1 0 588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1677622389
transform 1 0 572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1677622389
transform 1 0 580 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3532
timestamp 1677622389
transform 1 0 596 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1677622389
transform 1 0 580 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1677622389
transform 1 0 620 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3904
timestamp 1677622389
transform 1 0 628 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3533
timestamp 1677622389
transform 1 0 620 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1677622389
transform 1 0 628 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3993
timestamp 1677622389
transform 1 0 692 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3580
timestamp 1677622389
transform 1 0 692 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1677622389
transform 1 0 708 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3905
timestamp 1677622389
transform 1 0 732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1677622389
transform 1 0 708 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3560
timestamp 1677622389
transform 1 0 724 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1677622389
transform 1 0 780 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1677622389
transform 1 0 748 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3882
timestamp 1677622389
transform 1 0 796 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3562
timestamp 1677622389
transform 1 0 796 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1677622389
transform 1 0 828 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1677622389
transform 1 0 844 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3906
timestamp 1677622389
transform 1 0 828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1677622389
transform 1 0 844 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3534
timestamp 1677622389
transform 1 0 812 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3995
timestamp 1677622389
transform 1 0 820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1677622389
transform 1 0 836 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3563
timestamp 1677622389
transform 1 0 820 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1677622389
transform 1 0 836 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3997
timestamp 1677622389
transform 1 0 884 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3564
timestamp 1677622389
transform 1 0 884 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3908
timestamp 1677622389
transform 1 0 940 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3535
timestamp 1677622389
transform 1 0 932 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1677622389
transform 1 0 940 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3909
timestamp 1677622389
transform 1 0 964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1677622389
transform 1 0 964 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3566
timestamp 1677622389
transform 1 0 980 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3883
timestamp 1677622389
transform 1 0 1012 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3518
timestamp 1677622389
transform 1 0 1012 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1677622389
transform 1 0 1036 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1677622389
transform 1 0 1060 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3910
timestamp 1677622389
transform 1 0 1036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1677622389
transform 1 0 1052 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1677622389
transform 1 0 1060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1677622389
transform 1 0 1028 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3567
timestamp 1677622389
transform 1 0 1044 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4000
timestamp 1677622389
transform 1 0 1092 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1677622389
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3583
timestamp 1677622389
transform 1 0 1108 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3913
timestamp 1677622389
transform 1 0 1140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1677622389
transform 1 0 1156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1677622389
transform 1 0 1172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1677622389
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3437
timestamp 1677622389
transform 1 0 1196 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1677622389
transform 1 0 1196 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1677622389
transform 1 0 1212 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1677622389
transform 1 0 1236 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1677622389
transform 1 0 1228 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3916
timestamp 1677622389
transform 1 0 1276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1677622389
transform 1 0 1228 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3536
timestamp 1677622389
transform 1 0 1292 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1677622389
transform 1 0 1276 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3917
timestamp 1677622389
transform 1 0 1324 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1677622389
transform 1 0 1340 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4004
timestamp 1677622389
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1677622389
transform 1 0 1356 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3465
timestamp 1677622389
transform 1 0 1380 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1677622389
transform 1 0 1396 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3918
timestamp 1677622389
transform 1 0 1388 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3493
timestamp 1677622389
transform 1 0 1460 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1677622389
transform 1 0 1468 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3919
timestamp 1677622389
transform 1 0 1476 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1677622389
transform 1 0 1492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1677622389
transform 1 0 1460 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1677622389
transform 1 0 1468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1677622389
transform 1 0 1484 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3537
timestamp 1677622389
transform 1 0 1492 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4008
timestamp 1677622389
transform 1 0 1500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1677622389
transform 1 0 1508 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3569
timestamp 1677622389
transform 1 0 1484 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1677622389
transform 1 0 1468 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1677622389
transform 1 0 1508 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1677622389
transform 1 0 1532 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1677622389
transform 1 0 1556 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4010
timestamp 1677622389
transform 1 0 1580 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3494
timestamp 1677622389
transform 1 0 1596 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3921
timestamp 1677622389
transform 1 0 1596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1677622389
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1677622389
transform 1 0 1604 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3539
timestamp 1677622389
transform 1 0 1612 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1677622389
transform 1 0 1644 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1677622389
transform 1 0 1644 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1677622389
transform 1 0 1668 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1677622389
transform 1 0 1684 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1677622389
transform 1 0 1676 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3923
timestamp 1677622389
transform 1 0 1684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1677622389
transform 1 0 1676 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3496
timestamp 1677622389
transform 1 0 1748 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3924
timestamp 1677622389
transform 1 0 1748 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1677622389
transform 1 0 1772 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3586
timestamp 1677622389
transform 1 0 1772 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1677622389
transform 1 0 1804 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3925
timestamp 1677622389
transform 1 0 1804 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3440
timestamp 1677622389
transform 1 0 1836 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1677622389
transform 1 0 1828 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4014
timestamp 1677622389
transform 1 0 1844 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3469
timestamp 1677622389
transform 1 0 1860 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3926
timestamp 1677622389
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1677622389
transform 1 0 1940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1677622389
transform 1 0 1860 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3587
timestamp 1677622389
transform 1 0 1860 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1677622389
transform 1 0 1956 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1677622389
transform 1 0 1964 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1677622389
transform 1 0 1980 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3928
timestamp 1677622389
transform 1 0 1956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1677622389
transform 1 0 1972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1677622389
transform 1 0 1988 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1677622389
transform 1 0 1948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1677622389
transform 1 0 2012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1677622389
transform 1 0 1980 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1677622389
transform 1 0 1988 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3541
timestamp 1677622389
transform 1 0 1996 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1677622389
transform 1 0 1988 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1677622389
transform 1 0 2068 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1677622389
transform 1 0 2084 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3932
timestamp 1677622389
transform 1 0 2124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1677622389
transform 1 0 2180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1677622389
transform 1 0 2100 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3589
timestamp 1677622389
transform 1 0 2100 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1677622389
transform 1 0 2172 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1677622389
transform 1 0 2212 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3934
timestamp 1677622389
transform 1 0 2268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1677622389
transform 1 0 2316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1677622389
transform 1 0 2236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1677622389
transform 1 0 2332 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3543
timestamp 1677622389
transform 1 0 2332 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4021
timestamp 1677622389
transform 1 0 2340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1677622389
transform 1 0 2356 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3591
timestamp 1677622389
transform 1 0 2348 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3937
timestamp 1677622389
transform 1 0 2380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1677622389
transform 1 0 2388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1677622389
transform 1 0 2404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1677622389
transform 1 0 2412 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3441
timestamp 1677622389
transform 1 0 2436 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1677622389
transform 1 0 2452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1677622389
transform 1 0 2492 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3939
timestamp 1677622389
transform 1 0 2452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1677622389
transform 1 0 2460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1677622389
transform 1 0 2492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1677622389
transform 1 0 2540 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3450
timestamp 1677622389
transform 1 0 2564 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3942
timestamp 1677622389
transform 1 0 2556 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3544
timestamp 1677622389
transform 1 0 2556 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4026
timestamp 1677622389
transform 1 0 2588 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3442
timestamp 1677622389
transform 1 0 2620 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3943
timestamp 1677622389
transform 1 0 2612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1677622389
transform 1 0 2628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1677622389
transform 1 0 2636 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3592
timestamp 1677622389
transform 1 0 2628 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3944
timestamp 1677622389
transform 1 0 2644 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3502
timestamp 1677622389
transform 1 0 2676 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1677622389
transform 1 0 2700 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4029
timestamp 1677622389
transform 1 0 2700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1677622389
transform 1 0 2716 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3545
timestamp 1677622389
transform 1 0 2716 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1677622389
transform 1 0 2740 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3946
timestamp 1677622389
transform 1 0 2756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1677622389
transform 1 0 2748 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3593
timestamp 1677622389
transform 1 0 2748 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3947
timestamp 1677622389
transform 1 0 2780 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3594
timestamp 1677622389
transform 1 0 2812 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3948
timestamp 1677622389
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1677622389
transform 1 0 2844 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1677622389
transform 1 0 2860 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3547
timestamp 1677622389
transform 1 0 2860 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4032
timestamp 1677622389
transform 1 0 2868 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3472
timestamp 1677622389
transform 1 0 2924 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3886
timestamp 1677622389
transform 1 0 2924 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3548
timestamp 1677622389
transform 1 0 2916 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4065
timestamp 1677622389
transform 1 0 2908 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1677622389
transform 1 0 2932 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3443
timestamp 1677622389
transform 1 0 2964 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1677622389
transform 1 0 2956 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3949
timestamp 1677622389
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1677622389
transform 1 0 2972 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1677622389
transform 1 0 2948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1677622389
transform 1 0 2956 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3549
timestamp 1677622389
transform 1 0 2964 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3888
timestamp 1677622389
transform 1 0 2996 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1677622389
transform 1 0 3012 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3474
timestamp 1677622389
transform 1 0 3044 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3951
timestamp 1677622389
transform 1 0 3036 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3504
timestamp 1677622389
transform 1 0 3076 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3952
timestamp 1677622389
transform 1 0 3052 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3523
timestamp 1677622389
transform 1 0 3060 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3953
timestamp 1677622389
transform 1 0 3076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1677622389
transform 1 0 3044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1677622389
transform 1 0 3052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1677622389
transform 1 0 3068 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3550
timestamp 1677622389
transform 1 0 3076 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4039
timestamp 1677622389
transform 1 0 3084 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3571
timestamp 1677622389
transform 1 0 3068 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1677622389
transform 1 0 3068 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4040
timestamp 1677622389
transform 1 0 3108 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3451
timestamp 1677622389
transform 1 0 3148 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1677622389
transform 1 0 3172 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3954
timestamp 1677622389
transform 1 0 3156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1677622389
transform 1 0 3132 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3572
timestamp 1677622389
transform 1 0 3156 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1677622389
transform 1 0 3276 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1677622389
transform 1 0 3260 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3889
timestamp 1677622389
transform 1 0 3268 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1677622389
transform 1 0 3260 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3457
timestamp 1677622389
transform 1 0 3300 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3880
timestamp 1677622389
transform 1 0 3300 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1677622389
transform 1 0 3292 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3524
timestamp 1677622389
transform 1 0 3300 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3890
timestamp 1677622389
transform 1 0 3332 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3476
timestamp 1677622389
transform 1 0 3356 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1677622389
transform 1 0 3348 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3957
timestamp 1677622389
transform 1 0 3356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1677622389
transform 1 0 3356 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3596
timestamp 1677622389
transform 1 0 3364 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3891
timestamp 1677622389
transform 1 0 3388 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1677622389
transform 1 0 3436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1677622389
transform 1 0 3452 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_3507
timestamp 1677622389
transform 1 0 3452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1677622389
transform 1 0 3468 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1677622389
transform 1 0 3484 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3892
timestamp 1677622389
transform 1 0 3476 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3508
timestamp 1677622389
transform 1 0 3484 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3959
timestamp 1677622389
transform 1 0 3492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1677622389
transform 1 0 3516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1677622389
transform 1 0 3484 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1677622389
transform 1 0 3500 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3597
timestamp 1677622389
transform 1 0 3508 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1677622389
transform 1 0 3532 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4045
timestamp 1677622389
transform 1 0 3524 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3598
timestamp 1677622389
transform 1 0 3540 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1677622389
transform 1 0 3556 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1677622389
transform 1 0 3604 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3961
timestamp 1677622389
transform 1 0 3604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1677622389
transform 1 0 3660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1677622389
transform 1 0 3668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1677622389
transform 1 0 3580 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3573
timestamp 1677622389
transform 1 0 3580 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4047
timestamp 1677622389
transform 1 0 3700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1677622389
transform 1 0 3716 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3574
timestamp 1677622389
transform 1 0 3732 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1677622389
transform 1 0 3764 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1677622389
transform 1 0 3772 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3964
timestamp 1677622389
transform 1 0 3780 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3481
timestamp 1677622389
transform 1 0 3820 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3965
timestamp 1677622389
transform 1 0 3820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1677622389
transform 1 0 3836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1677622389
transform 1 0 3828 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3482
timestamp 1677622389
transform 1 0 3852 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3967
timestamp 1677622389
transform 1 0 3852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1677622389
transform 1 0 3852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1677622389
transform 1 0 3916 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3458
timestamp 1677622389
transform 1 0 3932 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1677622389
transform 1 0 3924 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3969
timestamp 1677622389
transform 1 0 3956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1677622389
transform 1 0 3932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1677622389
transform 1 0 3948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1677622389
transform 1 0 3964 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1677622389
transform 1 0 3972 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1677622389
transform 1 0 3988 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3511
timestamp 1677622389
transform 1 0 4044 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3971
timestamp 1677622389
transform 1 0 4028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1677622389
transform 1 0 4044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1677622389
transform 1 0 4020 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3453
timestamp 1677622389
transform 1 0 4076 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4056
timestamp 1677622389
transform 1 0 4076 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3575
timestamp 1677622389
transform 1 0 4076 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1677622389
transform 1 0 4100 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1677622389
transform 1 0 4132 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1677622389
transform 1 0 4124 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1677622389
transform 1 0 4092 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3973
timestamp 1677622389
transform 1 0 4116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1677622389
transform 1 0 4092 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3552
timestamp 1677622389
transform 1 0 4132 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1677622389
transform 1 0 4180 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1677622389
transform 1 0 4204 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1677622389
transform 1 0 4204 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3512
timestamp 1677622389
transform 1 0 4220 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1677622389
transform 1 0 4292 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1677622389
transform 1 0 4276 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1677622389
transform 1 0 4244 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1677622389
transform 1 0 4268 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1677622389
transform 1 0 4268 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3975
timestamp 1677622389
transform 1 0 4276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1677622389
transform 1 0 4244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1677622389
transform 1 0 4340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1677622389
transform 1 0 4348 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3576
timestamp 1677622389
transform 1 0 4332 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1677622389
transform 1 0 4444 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1677622389
transform 1 0 4404 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1677622389
transform 1 0 4452 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1677622389
transform 1 0 4380 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1677622389
transform 1 0 4404 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3978
timestamp 1677622389
transform 1 0 4404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1677622389
transform 1 0 4468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1677622389
transform 1 0 4452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1677622389
transform 1 0 4508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1677622389
transform 1 0 4540 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3446
timestamp 1677622389
transform 1 0 4556 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3980
timestamp 1677622389
transform 1 0 4572 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3515
timestamp 1677622389
transform 1 0 4660 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3981
timestamp 1677622389
transform 1 0 4612 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3528
timestamp 1677622389
transform 1 0 4636 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1677622389
transform 1 0 4660 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1677622389
transform 1 0 4612 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4062
timestamp 1677622389
transform 1 0 4660 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3516
timestamp 1677622389
transform 1 0 4708 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3982
timestamp 1677622389
transform 1 0 4708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1677622389
transform 1 0 4764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1677622389
transform 1 0 4772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1677622389
transform 1 0 4684 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3577
timestamp 1677622389
transform 1 0 4684 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1677622389
transform 1 0 4708 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4064
timestamp 1677622389
transform 1 0 4788 0 1 2805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_38
timestamp 1677622389
transform 1 0 48 0 1 2770
box -10 -3 10 3
use FILL  FILL_4375
timestamp 1677622389
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1677622389
transform 1 0 80 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_296
timestamp 1677622389
transform -1 0 104 0 1 2770
box -9 -3 26 105
use FILL  FILL_4378
timestamp 1677622389
transform 1 0 104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1677622389
transform 1 0 112 0 1 2770
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1677622389
transform 1 0 120 0 1 2770
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1677622389
transform 1 0 128 0 1 2770
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1677622389
transform 1 0 136 0 1 2770
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1677622389
transform 1 0 144 0 1 2770
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1677622389
transform 1 0 152 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_259
timestamp 1677622389
transform 1 0 160 0 1 2770
box -8 -3 104 105
use FILL  FILL_4385
timestamp 1677622389
transform 1 0 256 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_180
timestamp 1677622389
transform -1 0 304 0 1 2770
box -8 -3 46 105
use FILL  FILL_4386
timestamp 1677622389
transform 1 0 304 0 1 2770
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1677622389
transform 1 0 312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1677622389
transform 1 0 320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1677622389
transform 1 0 328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1677622389
transform 1 0 336 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1677622389
transform 1 0 344 0 1 2770
box -8 -3 104 105
use FILL  FILL_4391
timestamp 1677622389
transform 1 0 440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1677622389
transform 1 0 448 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_263
timestamp 1677622389
transform 1 0 456 0 1 2770
box -8 -3 104 105
use FILL  FILL_4400
timestamp 1677622389
transform 1 0 552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1677622389
transform 1 0 560 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_183
timestamp 1677622389
transform 1 0 568 0 1 2770
box -8 -3 46 105
use FILL  FILL_4411
timestamp 1677622389
transform 1 0 608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1677622389
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1677622389
transform 1 0 624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1677622389
transform 1 0 632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1677622389
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1677622389
transform 1 0 648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1677622389
transform 1 0 656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1677622389
transform 1 0 664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1677622389
transform 1 0 672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1677622389
transform 1 0 680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1677622389
transform 1 0 688 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1677622389
transform 1 0 696 0 1 2770
box -8 -3 104 105
use FILL  FILL_4425
timestamp 1677622389
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1677622389
transform 1 0 800 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_184
timestamp 1677622389
transform -1 0 848 0 1 2770
box -8 -3 46 105
use FILL  FILL_4427
timestamp 1677622389
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1677622389
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1677622389
transform 1 0 864 0 1 2770
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1677622389
transform 1 0 872 0 1 2770
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1677622389
transform 1 0 880 0 1 2770
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1677622389
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1677622389
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1677622389
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1677622389
transform 1 0 912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1677622389
transform 1 0 920 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_90
timestamp 1677622389
transform 1 0 928 0 1 2770
box -8 -3 34 105
use FILL  FILL_4457
timestamp 1677622389
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1677622389
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1677622389
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1677622389
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1677622389
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1677622389
transform 1 0 1000 0 1 2770
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1677622389
transform 1 0 1008 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_186
timestamp 1677622389
transform 1 0 1016 0 1 2770
box -8 -3 46 105
use FILL  FILL_4475
timestamp 1677622389
transform 1 0 1056 0 1 2770
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1677622389
transform 1 0 1064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1677622389
transform 1 0 1072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1677622389
transform 1 0 1080 0 1 2770
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1677622389
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1677622389
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1677622389
transform 1 0 1104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1677622389
transform 1 0 1112 0 1 2770
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1677622389
transform 1 0 1120 0 1 2770
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1677622389
transform 1 0 1128 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_188
timestamp 1677622389
transform 1 0 1136 0 1 2770
box -8 -3 46 105
use FILL  FILL_4495
timestamp 1677622389
transform 1 0 1176 0 1 2770
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1677622389
transform 1 0 1184 0 1 2770
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1677622389
transform 1 0 1192 0 1 2770
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1677622389
transform 1 0 1200 0 1 2770
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1677622389
transform 1 0 1208 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1677622389
transform 1 0 1216 0 1 2770
box -8 -3 104 105
use FILL  FILL_4500
timestamp 1677622389
transform 1 0 1312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1677622389
transform 1 0 1320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1677622389
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1677622389
transform 1 0 1336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1677622389
transform 1 0 1344 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_91
timestamp 1677622389
transform -1 0 1384 0 1 2770
box -8 -3 34 105
use FILL  FILL_4515
timestamp 1677622389
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1677622389
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1677622389
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1677622389
transform 1 0 1408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1677622389
transform 1 0 1416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1677622389
transform 1 0 1424 0 1 2770
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1677622389
transform 1 0 1432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1677622389
transform 1 0 1440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1677622389
transform 1 0 1448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1677622389
transform 1 0 1456 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_181
timestamp 1677622389
transform -1 0 1504 0 1 2770
box -8 -3 46 105
use FILL  FILL_4536
timestamp 1677622389
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1677622389
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1677622389
transform 1 0 1520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1677622389
transform 1 0 1528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1677622389
transform 1 0 1536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1677622389
transform 1 0 1544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1677622389
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1677622389
transform 1 0 1560 0 1 2770
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1677622389
transform 1 0 1568 0 1 2770
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1677622389
transform 1 0 1576 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_183
timestamp 1677622389
transform -1 0 1624 0 1 2770
box -8 -3 46 105
use FILL  FILL_4552
timestamp 1677622389
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1677622389
transform 1 0 1632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1677622389
transform 1 0 1640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1677622389
transform 1 0 1648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1677622389
transform 1 0 1656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1677622389
transform 1 0 1664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1677622389
transform 1 0 1672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1677622389
transform 1 0 1680 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1677622389
transform -1 0 1784 0 1 2770
box -8 -3 104 105
use FILL  FILL_4562
timestamp 1677622389
transform 1 0 1784 0 1 2770
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1677622389
transform 1 0 1792 0 1 2770
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1677622389
transform 1 0 1800 0 1 2770
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1677622389
transform 1 0 1808 0 1 2770
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1677622389
transform 1 0 1816 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_304
timestamp 1677622389
transform -1 0 1840 0 1 2770
box -9 -3 26 105
use FILL  FILL_4572
timestamp 1677622389
transform 1 0 1840 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_270
timestamp 1677622389
transform 1 0 1848 0 1 2770
box -8 -3 104 105
use FILL  FILL_4573
timestamp 1677622389
transform 1 0 1944 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_190
timestamp 1677622389
transform 1 0 1952 0 1 2770
box -8 -3 46 105
use FILL  FILL_4584
timestamp 1677622389
transform 1 0 1992 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_306
timestamp 1677622389
transform 1 0 2000 0 1 2770
box -9 -3 26 105
use FILL  FILL_4585
timestamp 1677622389
transform 1 0 2016 0 1 2770
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1677622389
transform 1 0 2024 0 1 2770
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1677622389
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1677622389
transform 1 0 2040 0 1 2770
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1677622389
transform 1 0 2048 0 1 2770
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1677622389
transform 1 0 2056 0 1 2770
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1677622389
transform 1 0 2064 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3599
timestamp 1677622389
transform 1 0 2084 0 1 2775
box -3 -3 3 3
use FILL  FILL_4592
timestamp 1677622389
transform 1 0 2072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1677622389
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_272
timestamp 1677622389
transform 1 0 2088 0 1 2770
box -8 -3 104 105
use FILL  FILL_4599
timestamp 1677622389
transform 1 0 2184 0 1 2770
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1677622389
transform 1 0 2192 0 1 2770
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1677622389
transform 1 0 2200 0 1 2770
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1677622389
transform 1 0 2208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1677622389
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_273
timestamp 1677622389
transform 1 0 2224 0 1 2770
box -8 -3 104 105
use FILL  FILL_4616
timestamp 1677622389
transform 1 0 2320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1677622389
transform 1 0 2328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1677622389
transform 1 0 2336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1677622389
transform 1 0 2344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1677622389
transform 1 0 2352 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_192
timestamp 1677622389
transform 1 0 2360 0 1 2770
box -8 -3 46 105
use FILL  FILL_4634
timestamp 1677622389
transform 1 0 2400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1677622389
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1677622389
transform 1 0 2416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1677622389
transform 1 0 2424 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_309
timestamp 1677622389
transform 1 0 2432 0 1 2770
box -9 -3 26 105
use FILL  FILL_4642
timestamp 1677622389
transform 1 0 2448 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1677622389
transform -1 0 2552 0 1 2770
box -8 -3 104 105
use FILL  FILL_4643
timestamp 1677622389
transform 1 0 2552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1677622389
transform 1 0 2560 0 1 2770
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1677622389
transform 1 0 2568 0 1 2770
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1677622389
transform 1 0 2576 0 1 2770
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1677622389
transform 1 0 2584 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_193
timestamp 1677622389
transform 1 0 2592 0 1 2770
box -8 -3 46 105
use FILL  FILL_4654
timestamp 1677622389
transform 1 0 2632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1677622389
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1677622389
transform 1 0 2648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1677622389
transform 1 0 2656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1677622389
transform 1 0 2664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1677622389
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_311
timestamp 1677622389
transform 1 0 2680 0 1 2770
box -9 -3 26 105
use FILL  FILL_4666
timestamp 1677622389
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1677622389
transform 1 0 2704 0 1 2770
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1677622389
transform 1 0 2712 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_312
timestamp 1677622389
transform 1 0 2720 0 1 2770
box -9 -3 26 105
use FILL  FILL_4669
timestamp 1677622389
transform 1 0 2736 0 1 2770
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1677622389
transform 1 0 2744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1677622389
transform 1 0 2752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1677622389
transform 1 0 2760 0 1 2770
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1677622389
transform 1 0 2768 0 1 2770
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1677622389
transform 1 0 2776 0 1 2770
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1677622389
transform 1 0 2784 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_93
timestamp 1677622389
transform 1 0 2792 0 1 2770
box -8 -3 34 105
use FILL  FILL_4676
timestamp 1677622389
transform 1 0 2824 0 1 2770
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1677622389
transform 1 0 2832 0 1 2770
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1677622389
transform 1 0 2840 0 1 2770
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1677622389
transform 1 0 2848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1677622389
transform 1 0 2856 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_94
timestamp 1677622389
transform 1 0 2864 0 1 2770
box -8 -3 34 105
use M3_M2  M3_M2_3600
timestamp 1677622389
transform 1 0 2908 0 1 2775
box -3 -3 3 3
use FILL  FILL_4689
timestamp 1677622389
transform 1 0 2896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1677622389
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1677622389
transform 1 0 2912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1677622389
transform 1 0 2920 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_47
timestamp 1677622389
transform 1 0 2928 0 1 2770
box -8 -3 32 105
use FILL  FILL_4697
timestamp 1677622389
transform 1 0 2952 0 1 2770
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1677622389
transform 1 0 2960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1677622389
transform 1 0 2968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1677622389
transform 1 0 2976 0 1 2770
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1677622389
transform 1 0 2984 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_97
timestamp 1677622389
transform -1 0 3024 0 1 2770
box -8 -3 34 105
use FILL  FILL_4706
timestamp 1677622389
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1677622389
transform 1 0 3032 0 1 2770
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1677622389
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_185
timestamp 1677622389
transform 1 0 3048 0 1 2770
box -8 -3 46 105
use FILL  FILL_4712
timestamp 1677622389
transform 1 0 3088 0 1 2770
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1677622389
transform 1 0 3096 0 1 2770
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1677622389
transform 1 0 3104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1677622389
transform 1 0 3112 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3601
timestamp 1677622389
transform 1 0 3196 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1677622389
transform 1 0 3220 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_277
timestamp 1677622389
transform 1 0 3120 0 1 2770
box -8 -3 104 105
use FILL  FILL_4720
timestamp 1677622389
transform 1 0 3216 0 1 2770
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1677622389
transform 1 0 3224 0 1 2770
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1677622389
transform 1 0 3232 0 1 2770
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1677622389
transform 1 0 3240 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3603
timestamp 1677622389
transform 1 0 3276 0 1 2775
box -3 -3 3 3
use INVX2  INVX2_314
timestamp 1677622389
transform 1 0 3248 0 1 2770
box -9 -3 26 105
use FILL  FILL_4733
timestamp 1677622389
transform 1 0 3264 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_23
timestamp 1677622389
transform -1 0 3304 0 1 2770
box -8 -3 40 105
use FILL  FILL_4734
timestamp 1677622389
transform 1 0 3304 0 1 2770
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1677622389
transform 1 0 3312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1677622389
transform 1 0 3320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1677622389
transform 1 0 3328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1677622389
transform 1 0 3336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1677622389
transform 1 0 3344 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_315
timestamp 1677622389
transform 1 0 3352 0 1 2770
box -9 -3 26 105
use FILL  FILL_4740
timestamp 1677622389
transform 1 0 3368 0 1 2770
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1677622389
transform 1 0 3376 0 1 2770
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1677622389
transform 1 0 3384 0 1 2770
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1677622389
transform 1 0 3392 0 1 2770
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1677622389
transform 1 0 3400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1677622389
transform 1 0 3408 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_24
timestamp 1677622389
transform -1 0 3448 0 1 2770
box -8 -3 40 105
use FILL  FILL_4752
timestamp 1677622389
transform 1 0 3448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1677622389
transform 1 0 3456 0 1 2770
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1677622389
transform 1 0 3464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1677622389
transform 1 0 3472 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3604
timestamp 1677622389
transform 1 0 3508 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_188
timestamp 1677622389
transform -1 0 3520 0 1 2770
box -8 -3 46 105
use FILL  FILL_4762
timestamp 1677622389
transform 1 0 3520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1677622389
transform 1 0 3528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1677622389
transform 1 0 3536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1677622389
transform 1 0 3544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1677622389
transform 1 0 3552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1677622389
transform 1 0 3560 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3605
timestamp 1677622389
transform 1 0 3668 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_279
timestamp 1677622389
transform 1 0 3568 0 1 2770
box -8 -3 104 105
use FILL  FILL_4775
timestamp 1677622389
transform 1 0 3664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1677622389
transform 1 0 3672 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_316
timestamp 1677622389
transform -1 0 3696 0 1 2770
box -9 -3 26 105
use FILL  FILL_4777
timestamp 1677622389
transform 1 0 3696 0 1 2770
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1677622389
transform 1 0 3704 0 1 2770
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1677622389
transform 1 0 3712 0 1 2770
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1677622389
transform 1 0 3720 0 1 2770
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1677622389
transform 1 0 3728 0 1 2770
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1677622389
transform 1 0 3736 0 1 2770
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1677622389
transform 1 0 3744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1677622389
transform 1 0 3752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1677622389
transform 1 0 3760 0 1 2770
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1677622389
transform 1 0 3768 0 1 2770
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1677622389
transform 1 0 3776 0 1 2770
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1677622389
transform 1 0 3784 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3606
timestamp 1677622389
transform 1 0 3804 0 1 2775
box -3 -3 3 3
use FILL  FILL_4801
timestamp 1677622389
transform 1 0 3792 0 1 2770
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1677622389
transform 1 0 3800 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_189
timestamp 1677622389
transform 1 0 3808 0 1 2770
box -8 -3 46 105
use FILL  FILL_4803
timestamp 1677622389
transform 1 0 3848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1677622389
transform 1 0 3856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1677622389
transform 1 0 3864 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_317
timestamp 1677622389
transform 1 0 3872 0 1 2770
box -9 -3 26 105
use FILL  FILL_4806
timestamp 1677622389
transform 1 0 3888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1677622389
transform 1 0 3896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1677622389
transform 1 0 3904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1677622389
transform 1 0 3912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1677622389
transform 1 0 3920 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_190
timestamp 1677622389
transform 1 0 3928 0 1 2770
box -8 -3 46 105
use FILL  FILL_4814
timestamp 1677622389
transform 1 0 3968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1677622389
transform 1 0 3976 0 1 2770
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1677622389
transform 1 0 3984 0 1 2770
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1677622389
transform 1 0 3992 0 1 2770
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1677622389
transform 1 0 4000 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_196
timestamp 1677622389
transform 1 0 4008 0 1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3607
timestamp 1677622389
transform 1 0 4060 0 1 2775
box -3 -3 3 3
use FILL  FILL_4825
timestamp 1677622389
transform 1 0 4048 0 1 2770
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1677622389
transform 1 0 4056 0 1 2770
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1677622389
transform 1 0 4064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1677622389
transform 1 0 4072 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3608
timestamp 1677622389
transform 1 0 4092 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1677622389
transform 1 0 4132 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_282
timestamp 1677622389
transform 1 0 4080 0 1 2770
box -8 -3 104 105
use FILL  FILL_4829
timestamp 1677622389
transform 1 0 4176 0 1 2770
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1677622389
transform 1 0 4184 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_319
timestamp 1677622389
transform 1 0 4192 0 1 2770
box -9 -3 26 105
use FILL  FILL_4831
timestamp 1677622389
transform 1 0 4208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1677622389
transform 1 0 4216 0 1 2770
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1677622389
transform 1 0 4224 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3610
timestamp 1677622389
transform 1 0 4244 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_284
timestamp 1677622389
transform 1 0 4232 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_320
timestamp 1677622389
transform 1 0 4328 0 1 2770
box -9 -3 26 105
use FILL  FILL_4846
timestamp 1677622389
transform 1 0 4344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1677622389
transform 1 0 4352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1677622389
transform 1 0 4360 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3611
timestamp 1677622389
transform 1 0 4452 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_285
timestamp 1677622389
transform -1 0 4464 0 1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3612
timestamp 1677622389
transform 1 0 4476 0 1 2775
box -3 -3 3 3
use FILL  FILL_4849
timestamp 1677622389
transform 1 0 4464 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_40
timestamp 1677622389
transform 1 0 4472 0 1 2770
box -5 -3 28 105
use FILL  FILL_4850
timestamp 1677622389
transform 1 0 4496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1677622389
transform 1 0 4504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1677622389
transform 1 0 4512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1677622389
transform 1 0 4520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1677622389
transform 1 0 4528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1677622389
transform 1 0 4536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1677622389
transform 1 0 4544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1677622389
transform 1 0 4552 0 1 2770
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1677622389
transform 1 0 4560 0 1 2770
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1677622389
transform 1 0 4568 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_287
timestamp 1677622389
transform -1 0 4672 0 1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3613
timestamp 1677622389
transform 1 0 4692 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1677622389
transform 1 0 4716 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_288
timestamp 1677622389
transform 1 0 4672 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_323
timestamp 1677622389
transform -1 0 4784 0 1 2770
box -9 -3 26 105
use FILL  FILL_4876
timestamp 1677622389
transform 1 0 4784 0 1 2770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_39
timestamp 1677622389
transform 1 0 4819 0 1 2770
box -10 -3 10 3
use M3_M2  M3_M2_3637
timestamp 1677622389
transform 1 0 84 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1677622389
transform 1 0 100 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4069
timestamp 1677622389
transform 1 0 100 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1677622389
transform 1 0 148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1677622389
transform 1 0 180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1677622389
transform 1 0 188 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3689
timestamp 1677622389
transform 1 0 148 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1677622389
transform 1 0 188 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1677622389
transform 1 0 180 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1677622389
transform 1 0 172 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4155
timestamp 1677622389
transform 1 0 204 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3615
timestamp 1677622389
transform 1 0 348 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1677622389
transform 1 0 284 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4070
timestamp 1677622389
transform 1 0 220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1677622389
transform 1 0 228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1677622389
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1677622389
transform 1 0 260 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3660
timestamp 1677622389
transform 1 0 268 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4074
timestamp 1677622389
transform 1 0 284 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3661
timestamp 1677622389
transform 1 0 308 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4156
timestamp 1677622389
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1677622389
transform 1 0 236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1677622389
transform 1 0 252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1677622389
transform 1 0 268 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1677622389
transform 1 0 308 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3691
timestamp 1677622389
transform 1 0 252 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1677622389
transform 1 0 228 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1677622389
transform 1 0 252 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1677622389
transform 1 0 332 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4161
timestamp 1677622389
transform 1 0 364 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1677622389
transform 1 0 388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1677622389
transform 1 0 412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1677622389
transform 1 0 420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1677622389
transform 1 0 436 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3680
timestamp 1677622389
transform 1 0 404 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4163
timestamp 1677622389
transform 1 0 412 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3681
timestamp 1677622389
transform 1 0 420 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4164
timestamp 1677622389
transform 1 0 428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1677622389
transform 1 0 444 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3692
timestamp 1677622389
transform 1 0 412 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1677622389
transform 1 0 492 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1677622389
transform 1 0 516 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4078
timestamp 1677622389
transform 1 0 516 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3662
timestamp 1677622389
transform 1 0 524 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4079
timestamp 1677622389
transform 1 0 532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1677622389
transform 1 0 508 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1677622389
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3694
timestamp 1677622389
transform 1 0 508 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1677622389
transform 1 0 532 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1677622389
transform 1 0 524 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1677622389
transform 1 0 564 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4080
timestamp 1677622389
transform 1 0 596 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3663
timestamp 1677622389
transform 1 0 676 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4168
timestamp 1677622389
transform 1 0 620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1677622389
transform 1 0 676 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1677622389
transform 1 0 692 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3664
timestamp 1677622389
transform 1 0 708 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4082
timestamp 1677622389
transform 1 0 716 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1677622389
transform 1 0 724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1677622389
transform 1 0 692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1677622389
transform 1 0 708 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3747
timestamp 1677622389
transform 1 0 716 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4172
timestamp 1677622389
transform 1 0 732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1677622389
transform 1 0 828 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1677622389
transform 1 0 836 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3665
timestamp 1677622389
transform 1 0 836 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4173
timestamp 1677622389
transform 1 0 964 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1677622389
transform 1 0 1036 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1677622389
transform 1 0 1052 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1677622389
transform 1 0 1044 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3735
timestamp 1677622389
transform 1 0 1044 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1677622389
transform 1 0 1044 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4175
timestamp 1677622389
transform 1 0 1068 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3749
timestamp 1677622389
transform 1 0 1076 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1677622389
transform 1 0 1132 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4086
timestamp 1677622389
transform 1 0 1132 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3642
timestamp 1677622389
transform 1 0 1156 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1677622389
transform 1 0 1156 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4176
timestamp 1677622389
transform 1 0 1156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3667
timestamp 1677622389
transform 1 0 1212 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1677622389
transform 1 0 1228 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4087
timestamp 1677622389
transform 1 0 1252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1677622389
transform 1 0 1172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1677622389
transform 1 0 1212 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1677622389
transform 1 0 1276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1677622389
transform 1 0 1292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1677622389
transform 1 0 1300 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1677622389
transform 1 0 1324 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3750
timestamp 1677622389
transform 1 0 1332 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4252
timestamp 1677622389
transform 1 0 1356 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1677622389
transform 1 0 1364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1677622389
transform 1 0 1388 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3716
timestamp 1677622389
transform 1 0 1436 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4090
timestamp 1677622389
transform 1 0 1460 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1677622389
transform 1 0 1468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1677622389
transform 1 0 1484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1677622389
transform 1 0 1476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1677622389
transform 1 0 1492 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3717
timestamp 1677622389
transform 1 0 1468 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1677622389
transform 1 0 1460 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4093
timestamp 1677622389
transform 1 0 1532 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3643
timestamp 1677622389
transform 1 0 1580 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4094
timestamp 1677622389
transform 1 0 1564 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3669
timestamp 1677622389
transform 1 0 1628 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4184
timestamp 1677622389
transform 1 0 1596 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3752
timestamp 1677622389
transform 1 0 1556 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1677622389
transform 1 0 1652 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4185
timestamp 1677622389
transform 1 0 1668 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1677622389
transform 1 0 1684 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3695
timestamp 1677622389
transform 1 0 1684 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1677622389
transform 1 0 1708 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4096
timestamp 1677622389
transform 1 0 1708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1677622389
transform 1 0 1724 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3696
timestamp 1677622389
transform 1 0 1716 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1677622389
transform 1 0 1756 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4097
timestamp 1677622389
transform 1 0 1756 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3697
timestamp 1677622389
transform 1 0 1740 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1677622389
transform 1 0 1772 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4098
timestamp 1677622389
transform 1 0 1780 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1677622389
transform 1 0 1764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1677622389
transform 1 0 1788 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3671
timestamp 1677622389
transform 1 0 1812 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4099
timestamp 1677622389
transform 1 0 1836 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3672
timestamp 1677622389
transform 1 0 1844 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4189
timestamp 1677622389
transform 1 0 1836 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3753
timestamp 1677622389
transform 1 0 1852 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4100
timestamp 1677622389
transform 1 0 1900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1677622389
transform 1 0 1908 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3673
timestamp 1677622389
transform 1 0 1916 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4190
timestamp 1677622389
transform 1 0 1900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1677622389
transform 1 0 1916 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3718
timestamp 1677622389
transform 1 0 1908 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1677622389
transform 1 0 1900 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4102
timestamp 1677622389
transform 1 0 1940 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1677622389
transform 1 0 1940 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3617
timestamp 1677622389
transform 1 0 2052 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4103
timestamp 1677622389
transform 1 0 1988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1677622389
transform 1 0 2084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1677622389
transform 1 0 2012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1677622389
transform 1 0 2068 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1677622389
transform 1 0 2076 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3719
timestamp 1677622389
transform 1 0 1980 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1677622389
transform 1 0 2084 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1677622389
transform 1 0 2100 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4196
timestamp 1677622389
transform 1 0 2132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1677622389
transform 1 0 2156 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3721
timestamp 1677622389
transform 1 0 2164 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1677622389
transform 1 0 2196 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4197
timestamp 1677622389
transform 1 0 2188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1677622389
transform 1 0 2236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1677622389
transform 1 0 2244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1677622389
transform 1 0 2268 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3722
timestamp 1677622389
transform 1 0 2268 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1677622389
transform 1 0 2316 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4108
timestamp 1677622389
transform 1 0 2316 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3621
timestamp 1677622389
transform 1 0 2340 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4109
timestamp 1677622389
transform 1 0 2340 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3674
timestamp 1677622389
transform 1 0 2364 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4199
timestamp 1677622389
transform 1 0 2364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3622
timestamp 1677622389
transform 1 0 2404 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1677622389
transform 1 0 2388 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1677622389
transform 1 0 2380 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4110
timestamp 1677622389
transform 1 0 2388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1677622389
transform 1 0 2404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1677622389
transform 1 0 2380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1677622389
transform 1 0 2396 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3723
timestamp 1677622389
transform 1 0 2396 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4202
timestamp 1677622389
transform 1 0 2444 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3623
timestamp 1677622389
transform 1 0 2460 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1677622389
transform 1 0 2484 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4112
timestamp 1677622389
transform 1 0 2532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1677622389
transform 1 0 2484 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3724
timestamp 1677622389
transform 1 0 2452 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4204
timestamp 1677622389
transform 1 0 2556 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3647
timestamp 1677622389
transform 1 0 2604 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4113
timestamp 1677622389
transform 1 0 2588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1677622389
transform 1 0 2604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1677622389
transform 1 0 2596 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3682
timestamp 1677622389
transform 1 0 2604 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4115
timestamp 1677622389
transform 1 0 2620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1677622389
transform 1 0 2612 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3683
timestamp 1677622389
transform 1 0 2620 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4207
timestamp 1677622389
transform 1 0 2644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1677622389
transform 1 0 2692 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3755
timestamp 1677622389
transform 1 0 2692 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1677622389
transform 1 0 2772 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4116
timestamp 1677622389
transform 1 0 2708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1677622389
transform 1 0 2740 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3756
timestamp 1677622389
transform 1 0 2716 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1677622389
transform 1 0 2764 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1677622389
transform 1 0 2804 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4068
timestamp 1677622389
transform 1 0 2804 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1677622389
transform 1 0 2812 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3628
timestamp 1677622389
transform 1 0 2828 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4117
timestamp 1677622389
transform 1 0 2836 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3684
timestamp 1677622389
transform 1 0 2836 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4211
timestamp 1677622389
transform 1 0 2844 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3629
timestamp 1677622389
transform 1 0 2868 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1677622389
transform 1 0 2860 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4118
timestamp 1677622389
transform 1 0 2860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1677622389
transform 1 0 2868 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3698
timestamp 1677622389
transform 1 0 2892 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4119
timestamp 1677622389
transform 1 0 2908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1677622389
transform 1 0 2916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1677622389
transform 1 0 2924 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3685
timestamp 1677622389
transform 1 0 2932 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4253
timestamp 1677622389
transform 1 0 2932 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3725
timestamp 1677622389
transform 1 0 2924 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1677622389
transform 1 0 2948 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1677622389
transform 1 0 2956 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4121
timestamp 1677622389
transform 1 0 2964 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1677622389
transform 1 0 2972 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1677622389
transform 1 0 2956 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3686
timestamp 1677622389
transform 1 0 2972 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4254
timestamp 1677622389
transform 1 0 2972 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3726
timestamp 1677622389
transform 1 0 2972 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1677622389
transform 1 0 3012 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4215
timestamp 1677622389
transform 1 0 3012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1677622389
transform 1 0 2996 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1677622389
transform 1 0 3036 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3652
timestamp 1677622389
transform 1 0 3060 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4123
timestamp 1677622389
transform 1 0 3060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1677622389
transform 1 0 3068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1677622389
transform 1 0 3084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1677622389
transform 1 0 3052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1677622389
transform 1 0 3076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1677622389
transform 1 0 3092 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3699
timestamp 1677622389
transform 1 0 3076 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1677622389
transform 1 0 3076 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4126
timestamp 1677622389
transform 1 0 3108 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3728
timestamp 1677622389
transform 1 0 3108 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1677622389
transform 1 0 3140 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4127
timestamp 1677622389
transform 1 0 3148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1677622389
transform 1 0 3140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1677622389
transform 1 0 3156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3700
timestamp 1677622389
transform 1 0 3156 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4128
timestamp 1677622389
transform 1 0 3180 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3654
timestamp 1677622389
transform 1 0 3212 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4129
timestamp 1677622389
transform 1 0 3204 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1677622389
transform 1 0 3212 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3701
timestamp 1677622389
transform 1 0 3220 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1677622389
transform 1 0 3244 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1677622389
transform 1 0 3268 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1677622389
transform 1 0 3308 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4130
timestamp 1677622389
transform 1 0 3276 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1677622389
transform 1 0 3300 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1677622389
transform 1 0 3356 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3758
timestamp 1677622389
transform 1 0 3348 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4256
timestamp 1677622389
transform 1 0 3396 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1677622389
transform 1 0 3388 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3632
timestamp 1677622389
transform 1 0 3420 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4265
timestamp 1677622389
transform 1 0 3412 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3759
timestamp 1677622389
transform 1 0 3396 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4131
timestamp 1677622389
transform 1 0 3436 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3760
timestamp 1677622389
transform 1 0 3436 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1677622389
transform 1 0 3460 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1677622389
transform 1 0 3500 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4132
timestamp 1677622389
transform 1 0 3492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1677622389
transform 1 0 3508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1677622389
transform 1 0 3516 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1677622389
transform 1 0 3476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1677622389
transform 1 0 3468 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3687
timestamp 1677622389
transform 1 0 3484 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4226
timestamp 1677622389
transform 1 0 3500 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1677622389
transform 1 0 3516 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3703
timestamp 1677622389
transform 1 0 3516 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1677622389
transform 1 0 3492 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4135
timestamp 1677622389
transform 1 0 3580 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3704
timestamp 1677622389
transform 1 0 3588 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4136
timestamp 1677622389
transform 1 0 3620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1677622389
transform 1 0 3644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1677622389
transform 1 0 3700 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3705
timestamp 1677622389
transform 1 0 3620 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1677622389
transform 1 0 3644 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4258
timestamp 1677622389
transform 1 0 3740 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1677622389
transform 1 0 3748 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3736
timestamp 1677622389
transform 1 0 3748 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4259
timestamp 1677622389
transform 1 0 3788 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1677622389
transform 1 0 3788 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1677622389
transform 1 0 3788 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1677622389
transform 1 0 3836 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4137
timestamp 1677622389
transform 1 0 3804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1677622389
transform 1 0 3828 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3688
timestamp 1677622389
transform 1 0 3836 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1677622389
transform 1 0 3924 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4231
timestamp 1677622389
transform 1 0 3924 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1677622389
transform 1 0 3932 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3738
timestamp 1677622389
transform 1 0 3932 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1677622389
transform 1 0 3980 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4232
timestamp 1677622389
transform 1 0 3988 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1677622389
transform 1 0 3980 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3729
timestamp 1677622389
transform 1 0 3988 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4261
timestamp 1677622389
transform 1 0 4028 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3739
timestamp 1677622389
transform 1 0 4036 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4233
timestamp 1677622389
transform 1 0 4076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1677622389
transform 1 0 4060 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1677622389
transform 1 0 4076 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1677622389
transform 1 0 4076 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3740
timestamp 1677622389
transform 1 0 4068 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1677622389
transform 1 0 4124 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1677622389
transform 1 0 4196 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4138
timestamp 1677622389
transform 1 0 4132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1677622389
transform 1 0 4180 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3706
timestamp 1677622389
transform 1 0 4180 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1677622389
transform 1 0 4180 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1677622389
transform 1 0 4220 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1677622389
transform 1 0 4236 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4235
timestamp 1677622389
transform 1 0 4252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1677622389
transform 1 0 4300 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3677
timestamp 1677622389
transform 1 0 4308 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4236
timestamp 1677622389
transform 1 0 4308 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3742
timestamp 1677622389
transform 1 0 4316 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1677622389
transform 1 0 4332 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4140
timestamp 1677622389
transform 1 0 4324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1677622389
transform 1 0 4340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1677622389
transform 1 0 4364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1677622389
transform 1 0 4380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1677622389
transform 1 0 4356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1677622389
transform 1 0 4372 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3708
timestamp 1677622389
transform 1 0 4364 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1677622389
transform 1 0 4388 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4240
timestamp 1677622389
transform 1 0 4388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1677622389
transform 1 0 4476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1677622389
transform 1 0 4428 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3709
timestamp 1677622389
transform 1 0 4428 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1677622389
transform 1 0 4436 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1677622389
transform 1 0 4476 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4144
timestamp 1677622389
transform 1 0 4508 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3745
timestamp 1677622389
transform 1 0 4516 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4145
timestamp 1677622389
transform 1 0 4532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1677622389
transform 1 0 4540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1677622389
transform 1 0 4556 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3730
timestamp 1677622389
transform 1 0 4540 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4244
timestamp 1677622389
transform 1 0 4572 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3746
timestamp 1677622389
transform 1 0 4572 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4146
timestamp 1677622389
transform 1 0 4580 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1677622389
transform 1 0 4588 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3710
timestamp 1677622389
transform 1 0 4580 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4148
timestamp 1677622389
transform 1 0 4612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1677622389
transform 1 0 4620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1677622389
transform 1 0 4628 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3658
timestamp 1677622389
transform 1 0 4660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4149
timestamp 1677622389
transform 1 0 4660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1677622389
transform 1 0 4652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1677622389
transform 1 0 4668 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3711
timestamp 1677622389
transform 1 0 4668 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4150
timestamp 1677622389
transform 1 0 4692 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3659
timestamp 1677622389
transform 1 0 4732 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4151
timestamp 1677622389
transform 1 0 4708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1677622389
transform 1 0 4732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1677622389
transform 1 0 4788 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1677622389
transform 1 0 4772 0 1 2715
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_40
timestamp 1677622389
transform 1 0 24 0 1 2670
box -10 -3 10 3
use FILL  FILL_4376
timestamp 1677622389
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1677622389
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1677622389
transform 1 0 88 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_297
timestamp 1677622389
transform -1 0 200 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4394
timestamp 1677622389
transform 1 0 200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1677622389
transform 1 0 208 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_181
timestamp 1677622389
transform -1 0 256 0 -1 2770
box -8 -3 46 105
use INVX2  INVX2_298
timestamp 1677622389
transform 1 0 256 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1677622389
transform 1 0 272 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4396
timestamp 1677622389
transform 1 0 368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1677622389
transform 1 0 376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1677622389
transform 1 0 384 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_299
timestamp 1677622389
transform -1 0 408 0 -1 2770
box -9 -3 26 105
use AOI22X1  AOI22X1_182
timestamp 1677622389
transform 1 0 408 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4399
timestamp 1677622389
transform 1 0 448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1677622389
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1677622389
transform 1 0 464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1677622389
transform 1 0 472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1677622389
transform 1 0 480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1677622389
transform 1 0 488 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_180
timestamp 1677622389
transform 1 0 496 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4406
timestamp 1677622389
transform 1 0 536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1677622389
transform 1 0 544 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3763
timestamp 1677622389
transform 1 0 572 0 1 2675
box -3 -3 3 3
use FILL  FILL_4408
timestamp 1677622389
transform 1 0 552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1677622389
transform 1 0 560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1677622389
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1677622389
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1677622389
transform 1 0 584 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4423
timestamp 1677622389
transform 1 0 680 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_185
timestamp 1677622389
transform 1 0 688 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4428
timestamp 1677622389
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1677622389
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1677622389
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1677622389
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1677622389
transform 1 0 760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1677622389
transform 1 0 768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1677622389
transform 1 0 776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1677622389
transform 1 0 784 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_300
timestamp 1677622389
transform -1 0 808 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4436
timestamp 1677622389
transform 1 0 808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1677622389
transform 1 0 816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1677622389
transform 1 0 824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1677622389
transform 1 0 832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1677622389
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1677622389
transform 1 0 848 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_45
timestamp 1677622389
transform 1 0 856 0 -1 2770
box -8 -3 32 105
use FILL  FILL_4446
timestamp 1677622389
transform 1 0 880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1677622389
transform 1 0 888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1677622389
transform 1 0 896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1677622389
transform 1 0 904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1677622389
transform 1 0 912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1677622389
transform 1 0 920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1677622389
transform 1 0 928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1677622389
transform 1 0 936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1677622389
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1677622389
transform 1 0 952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1677622389
transform 1 0 960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1677622389
transform 1 0 968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1677622389
transform 1 0 976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1677622389
transform 1 0 984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1677622389
transform 1 0 992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1677622389
transform 1 0 1000 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3764
timestamp 1677622389
transform 1 0 1020 0 1 2675
box -3 -3 3 3
use FILL  FILL_4474
timestamp 1677622389
transform 1 0 1008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1677622389
transform 1 0 1016 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_187
timestamp 1677622389
transform 1 0 1024 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4478
timestamp 1677622389
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1677622389
transform 1 0 1072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1677622389
transform 1 0 1080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1677622389
transform 1 0 1088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1677622389
transform 1 0 1096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1677622389
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1677622389
transform 1 0 1112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1677622389
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1677622389
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3765
timestamp 1677622389
transform 1 0 1156 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_301
timestamp 1677622389
transform 1 0 1136 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4501
timestamp 1677622389
transform 1 0 1152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1677622389
transform 1 0 1160 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_267
timestamp 1677622389
transform -1 0 1264 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4503
timestamp 1677622389
transform 1 0 1264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1677622389
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_302
timestamp 1677622389
transform -1 0 1296 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4505
timestamp 1677622389
transform 1 0 1296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1677622389
transform 1 0 1304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1677622389
transform 1 0 1312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1677622389
transform 1 0 1320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1677622389
transform 1 0 1328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1677622389
transform 1 0 1336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1677622389
transform 1 0 1344 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3766
timestamp 1677622389
transform 1 0 1364 0 1 2675
box -3 -3 3 3
use FILL  FILL_4518
timestamp 1677622389
transform 1 0 1352 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_92
timestamp 1677622389
transform -1 0 1392 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4519
timestamp 1677622389
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1677622389
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1677622389
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1677622389
transform 1 0 1416 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3767
timestamp 1677622389
transform 1 0 1436 0 1 2675
box -3 -3 3 3
use FILL  FILL_4527
timestamp 1677622389
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1677622389
transform 1 0 1432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1677622389
transform 1 0 1440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1677622389
transform 1 0 1448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1677622389
transform 1 0 1456 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_182
timestamp 1677622389
transform -1 0 1504 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4537
timestamp 1677622389
transform 1 0 1504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1677622389
transform 1 0 1512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1677622389
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1677622389
transform 1 0 1528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1677622389
transform 1 0 1536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1677622389
transform 1 0 1544 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3768
timestamp 1677622389
transform 1 0 1564 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_268
timestamp 1677622389
transform 1 0 1552 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4556
timestamp 1677622389
transform 1 0 1648 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_303
timestamp 1677622389
transform 1 0 1656 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4560
timestamp 1677622389
transform 1 0 1672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1677622389
transform 1 0 1680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1677622389
transform 1 0 1688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1677622389
transform 1 0 1696 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_36
timestamp 1677622389
transform -1 0 1728 0 -1 2770
box -5 -3 28 105
use FILL  FILL_4569
timestamp 1677622389
transform 1 0 1728 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_37
timestamp 1677622389
transform 1 0 1736 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_38
timestamp 1677622389
transform 1 0 1760 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_39
timestamp 1677622389
transform 1 0 1784 0 -1 2770
box -5 -3 28 105
use FILL  FILL_4570
timestamp 1677622389
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1677622389
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1677622389
transform 1 0 1824 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_305
timestamp 1677622389
transform 1 0 1832 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4576
timestamp 1677622389
transform 1 0 1848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1677622389
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1677622389
transform 1 0 1864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1677622389
transform 1 0 1872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1677622389
transform 1 0 1880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1677622389
transform 1 0 1888 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3769
timestamp 1677622389
transform 1 0 1924 0 1 2675
box -3 -3 3 3
use AOI22X1  AOI22X1_189
timestamp 1677622389
transform 1 0 1896 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4582
timestamp 1677622389
transform 1 0 1936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1677622389
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1677622389
transform 1 0 1952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1677622389
transform 1 0 1960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1677622389
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_271
timestamp 1677622389
transform 1 0 1976 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4596
timestamp 1677622389
transform 1 0 2072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1677622389
transform 1 0 2080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1677622389
transform 1 0 2088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1677622389
transform 1 0 2096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1677622389
transform 1 0 2104 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_191
timestamp 1677622389
transform 1 0 2112 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4603
timestamp 1677622389
transform 1 0 2152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1677622389
transform 1 0 2160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1677622389
transform 1 0 2168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1677622389
transform 1 0 2176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1677622389
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1677622389
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1677622389
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1677622389
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1677622389
transform 1 0 2216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1677622389
transform 1 0 2224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1677622389
transform 1 0 2232 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_307
timestamp 1677622389
transform 1 0 2240 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4620
timestamp 1677622389
transform 1 0 2256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1677622389
transform 1 0 2264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1677622389
transform 1 0 2272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1677622389
transform 1 0 2280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1677622389
transform 1 0 2288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1677622389
transform 1 0 2296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1677622389
transform 1 0 2304 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_308
timestamp 1677622389
transform 1 0 2312 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4627
timestamp 1677622389
transform 1 0 2328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1677622389
transform 1 0 2336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1677622389
transform 1 0 2344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1677622389
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1677622389
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_184
timestamp 1677622389
transform 1 0 2368 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4637
timestamp 1677622389
transform 1 0 2408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1677622389
transform 1 0 2416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1677622389
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1677622389
transform 1 0 2432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1677622389
transform 1 0 2440 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3770
timestamp 1677622389
transform 1 0 2524 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1677622389
transform 1 0 2540 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_275
timestamp 1677622389
transform -1 0 2544 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4646
timestamp 1677622389
transform 1 0 2544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1677622389
transform 1 0 2552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1677622389
transform 1 0 2560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1677622389
transform 1 0 2568 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_194
timestamp 1677622389
transform 1 0 2576 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4655
timestamp 1677622389
transform 1 0 2616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1677622389
transform 1 0 2624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1677622389
transform 1 0 2632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1677622389
transform 1 0 2640 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_310
timestamp 1677622389
transform 1 0 2648 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4663
timestamp 1677622389
transform 1 0 2664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1677622389
transform 1 0 2672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1677622389
transform 1 0 2680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1677622389
transform 1 0 2688 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1677622389
transform 1 0 2696 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4682
timestamp 1677622389
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1677622389
transform 1 0 2800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1677622389
transform 1 0 2808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1677622389
transform 1 0 2816 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_46
timestamp 1677622389
transform 1 0 2824 0 -1 2770
box -8 -3 32 105
use FILL  FILL_4686
timestamp 1677622389
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1677622389
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1677622389
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_95
timestamp 1677622389
transform 1 0 2872 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4692
timestamp 1677622389
transform 1 0 2904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1677622389
transform 1 0 2912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1677622389
transform 1 0 2920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1677622389
transform 1 0 2928 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_96
timestamp 1677622389
transform -1 0 2968 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4701
timestamp 1677622389
transform 1 0 2968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1677622389
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1677622389
transform 1 0 2984 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_98
timestamp 1677622389
transform -1 0 3024 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4707
timestamp 1677622389
transform 1 0 3024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1677622389
transform 1 0 3032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1677622389
transform 1 0 3040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1677622389
transform 1 0 3048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1677622389
transform 1 0 3056 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_186
timestamp 1677622389
transform 1 0 3064 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4717
timestamp 1677622389
transform 1 0 3104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1677622389
transform 1 0 3112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1677622389
transform 1 0 3120 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_187
timestamp 1677622389
transform -1 0 3168 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4723
timestamp 1677622389
transform 1 0 3168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1677622389
transform 1 0 3176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1677622389
transform 1 0 3184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1677622389
transform 1 0 3192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1677622389
transform 1 0 3200 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_313
timestamp 1677622389
transform 1 0 3208 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4728
timestamp 1677622389
transform 1 0 3224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1677622389
transform 1 0 3232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1677622389
transform 1 0 3240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1677622389
transform 1 0 3248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1677622389
transform 1 0 3256 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_278
timestamp 1677622389
transform 1 0 3264 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4743
timestamp 1677622389
transform 1 0 3360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1677622389
transform 1 0 3368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1677622389
transform 1 0 3376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1677622389
transform 1 0 3384 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3772
timestamp 1677622389
transform 1 0 3412 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_25
timestamp 1677622389
transform 1 0 3392 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4753
timestamp 1677622389
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1677622389
transform 1 0 3432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1677622389
transform 1 0 3440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1677622389
transform 1 0 3448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1677622389
transform 1 0 3456 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3773
timestamp 1677622389
transform 1 0 3484 0 1 2675
box -3 -3 3 3
use FILL  FILL_4760
timestamp 1677622389
transform 1 0 3464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1677622389
transform 1 0 3472 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_195
timestamp 1677622389
transform 1 0 3480 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4764
timestamp 1677622389
transform 1 0 3520 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3774
timestamp 1677622389
transform 1 0 3540 0 1 2675
box -3 -3 3 3
use FILL  FILL_4766
timestamp 1677622389
transform 1 0 3528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1677622389
transform 1 0 3536 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3775
timestamp 1677622389
transform 1 0 3556 0 1 2675
box -3 -3 3 3
use FILL  FILL_4770
timestamp 1677622389
transform 1 0 3544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1677622389
transform 1 0 3552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1677622389
transform 1 0 3560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1677622389
transform 1 0 3568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1677622389
transform 1 0 3576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1677622389
transform 1 0 3584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1677622389
transform 1 0 3592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1677622389
transform 1 0 3600 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3776
timestamp 1677622389
transform 1 0 3644 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1677622389
transform 1 0 3692 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_280
timestamp 1677622389
transform 1 0 3608 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4784
timestamp 1677622389
transform 1 0 3704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1677622389
transform 1 0 3712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1677622389
transform 1 0 3720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1677622389
transform 1 0 3728 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3778
timestamp 1677622389
transform 1 0 3764 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_26
timestamp 1677622389
transform -1 0 3768 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4796
timestamp 1677622389
transform 1 0 3768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1677622389
transform 1 0 3776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1677622389
transform 1 0 3784 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1677622389
transform 1 0 3792 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4807
timestamp 1677622389
transform 1 0 3888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1677622389
transform 1 0 3896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1677622389
transform 1 0 3904 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_318
timestamp 1677622389
transform 1 0 3912 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4819
timestamp 1677622389
transform 1 0 3928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1677622389
transform 1 0 3936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1677622389
transform 1 0 3944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1677622389
transform 1 0 3952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1677622389
transform 1 0 3960 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_27
timestamp 1677622389
transform -1 0 4000 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4824
timestamp 1677622389
transform 1 0 4000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1677622389
transform 1 0 4008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1677622389
transform 1 0 4016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1677622389
transform 1 0 4024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1677622389
transform 1 0 4032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1677622389
transform 1 0 4040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1677622389
transform 1 0 4048 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_28
timestamp 1677622389
transform -1 0 4088 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4839
timestamp 1677622389
transform 1 0 4088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1677622389
transform 1 0 4096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1677622389
transform 1 0 4104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1677622389
transform 1 0 4112 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1677622389
transform 1 0 4120 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4843
timestamp 1677622389
transform 1 0 4216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1677622389
transform 1 0 4224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1677622389
transform 1 0 4232 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_321
timestamp 1677622389
transform 1 0 4240 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4852
timestamp 1677622389
transform 1 0 4256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1677622389
transform 1 0 4264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1677622389
transform 1 0 4272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1677622389
transform 1 0 4280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1677622389
transform 1 0 4288 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_322
timestamp 1677622389
transform 1 0 4296 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4857
timestamp 1677622389
transform 1 0 4312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1677622389
transform 1 0 4320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1677622389
transform 1 0 4328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1677622389
transform 1 0 4336 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_191
timestamp 1677622389
transform -1 0 4384 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4861
timestamp 1677622389
transform 1 0 4384 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_286
timestamp 1677622389
transform -1 0 4488 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4862
timestamp 1677622389
transform 1 0 4488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1677622389
transform 1 0 4496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1677622389
transform 1 0 4504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1677622389
transform 1 0 4512 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_197
timestamp 1677622389
transform 1 0 4520 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4874
timestamp 1677622389
transform 1 0 4560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1677622389
transform 1 0 4568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1677622389
transform 1 0 4576 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_324
timestamp 1677622389
transform 1 0 4584 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4879
timestamp 1677622389
transform 1 0 4600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1677622389
transform 1 0 4608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1677622389
transform 1 0 4616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1677622389
transform 1 0 4624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1677622389
transform 1 0 4632 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_192
timestamp 1677622389
transform 1 0 4640 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4884
timestamp 1677622389
transform 1 0 4680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1677622389
transform 1 0 4688 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_289
timestamp 1677622389
transform 1 0 4696 0 -1 2770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_41
timestamp 1677622389
transform 1 0 4843 0 1 2670
box -10 -3 10 3
use M3_M2  M3_M2_3821
timestamp 1677622389
transform 1 0 164 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1677622389
transform 1 0 132 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1677622389
transform 1 0 172 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4285
timestamp 1677622389
transform 1 0 132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1677622389
transform 1 0 164 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1677622389
transform 1 0 172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1677622389
transform 1 0 84 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3956
timestamp 1677622389
transform 1 0 68 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1677622389
transform 1 0 196 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1677622389
transform 1 0 228 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4288
timestamp 1677622389
transform 1 0 180 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3865
timestamp 1677622389
transform 1 0 196 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4289
timestamp 1677622389
transform 1 0 204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1677622389
transform 1 0 228 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3893
timestamp 1677622389
transform 1 0 180 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4395
timestamp 1677622389
transform 1 0 188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1677622389
transform 1 0 196 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1677622389
transform 1 0 212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1677622389
transform 1 0 220 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3894
timestamp 1677622389
transform 1 0 228 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4399
timestamp 1677622389
transform 1 0 236 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3919
timestamp 1677622389
transform 1 0 212 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1677622389
transform 1 0 236 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1677622389
transform 1 0 260 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1677622389
transform 1 0 292 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1677622389
transform 1 0 284 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4291
timestamp 1677622389
transform 1 0 260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1677622389
transform 1 0 276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1677622389
transform 1 0 292 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3866
timestamp 1677622389
transform 1 0 300 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4294
timestamp 1677622389
transform 1 0 308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1677622389
transform 1 0 284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1677622389
transform 1 0 300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1677622389
transform 1 0 316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1677622389
transform 1 0 332 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3957
timestamp 1677622389
transform 1 0 260 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4295
timestamp 1677622389
transform 1 0 348 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3921
timestamp 1677622389
transform 1 0 348 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1677622389
transform 1 0 452 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1677622389
transform 1 0 444 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1677622389
transform 1 0 364 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1677622389
transform 1 0 364 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1677622389
transform 1 0 396 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4296
timestamp 1677622389
transform 1 0 412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1677622389
transform 1 0 364 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3809
timestamp 1677622389
transform 1 0 468 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1677622389
transform 1 0 460 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1677622389
transform 1 0 500 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1677622389
transform 1 0 492 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4297
timestamp 1677622389
transform 1 0 460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1677622389
transform 1 0 468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1677622389
transform 1 0 484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1677622389
transform 1 0 500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1677622389
transform 1 0 452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1677622389
transform 1 0 492 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3922
timestamp 1677622389
transform 1 0 500 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4301
timestamp 1677622389
transform 1 0 516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1677622389
transform 1 0 532 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3779
timestamp 1677622389
transform 1 0 564 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4303
timestamp 1677622389
transform 1 0 564 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3869
timestamp 1677622389
transform 1 0 572 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4407
timestamp 1677622389
transform 1 0 556 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3895
timestamp 1677622389
transform 1 0 564 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4408
timestamp 1677622389
transform 1 0 572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1677622389
transform 1 0 620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1677622389
transform 1 0 668 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3870
timestamp 1677622389
transform 1 0 676 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4409
timestamp 1677622389
transform 1 0 676 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3810
timestamp 1677622389
transform 1 0 692 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4410
timestamp 1677622389
transform 1 0 692 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3871
timestamp 1677622389
transform 1 0 708 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4411
timestamp 1677622389
transform 1 0 724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1677622389
transform 1 0 764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1677622389
transform 1 0 796 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1677622389
transform 1 0 828 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3872
timestamp 1677622389
transform 1 0 828 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4412
timestamp 1677622389
transform 1 0 836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1677622389
transform 1 0 852 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3923
timestamp 1677622389
transform 1 0 860 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1677622389
transform 1 0 924 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4308
timestamp 1677622389
transform 1 0 924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1677622389
transform 1 0 916 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3924
timestamp 1677622389
transform 1 0 932 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4309
timestamp 1677622389
transform 1 0 948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1677622389
transform 1 0 948 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3896
timestamp 1677622389
transform 1 0 956 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4490
timestamp 1677622389
transform 1 0 956 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3794
timestamp 1677622389
transform 1 0 988 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4415
timestamp 1677622389
transform 1 0 1012 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3897
timestamp 1677622389
transform 1 0 1036 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4416
timestamp 1677622389
transform 1 0 1044 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3795
timestamp 1677622389
transform 1 0 1068 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4310
timestamp 1677622389
transform 1 0 1060 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1677622389
transform 1 0 1068 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3898
timestamp 1677622389
transform 1 0 1068 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1677622389
transform 1 0 1060 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4312
timestamp 1677622389
transform 1 0 1100 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3873
timestamp 1677622389
transform 1 0 1108 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4417
timestamp 1677622389
transform 1 0 1100 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3926
timestamp 1677622389
transform 1 0 1100 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4418
timestamp 1677622389
transform 1 0 1108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1677622389
transform 1 0 1124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1677622389
transform 1 0 1156 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1677622389
transform 1 0 1172 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3874
timestamp 1677622389
transform 1 0 1180 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1677622389
transform 1 0 1228 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4270
timestamp 1677622389
transform 1 0 1220 0 1 2655
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1677622389
transform 1 0 1220 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3875
timestamp 1677622389
transform 1 0 1220 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1677622389
transform 1 0 1220 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4419
timestamp 1677622389
transform 1 0 1236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1677622389
transform 1 0 1252 0 1 2655
box -2 -2 2 2
use M3_M2  M3_M2_3811
timestamp 1677622389
transform 1 0 1260 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1677622389
transform 1 0 1260 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4491
timestamp 1677622389
transform 1 0 1276 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1677622389
transform 1 0 1284 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1677622389
transform 1 0 1284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1677622389
transform 1 0 1300 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3928
timestamp 1677622389
transform 1 0 1284 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1677622389
transform 1 0 1308 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4420
timestamp 1677622389
transform 1 0 1348 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3929
timestamp 1677622389
transform 1 0 1348 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4421
timestamp 1677622389
transform 1 0 1372 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1677622389
transform 1 0 1388 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3876
timestamp 1677622389
transform 1 0 1396 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1677622389
transform 1 0 1452 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1677622389
transform 1 0 1476 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1677622389
transform 1 0 1436 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4318
timestamp 1677622389
transform 1 0 1484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1677622389
transform 1 0 1436 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3900
timestamp 1677622389
transform 1 0 1460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1677622389
transform 1 0 1524 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1677622389
transform 1 0 1548 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4319
timestamp 1677622389
transform 1 0 1556 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3812
timestamp 1677622389
transform 1 0 1572 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4320
timestamp 1677622389
transform 1 0 1564 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3930
timestamp 1677622389
transform 1 0 1564 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1677622389
transform 1 0 1620 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4423
timestamp 1677622389
transform 1 0 1628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1677622389
transform 1 0 1652 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1677622389
transform 1 0 1660 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1677622389
transform 1 0 1676 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1677622389
transform 1 0 1692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1677622389
transform 1 0 1668 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1677622389
transform 1 0 1684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1677622389
transform 1 0 1716 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3798
timestamp 1677622389
transform 1 0 1748 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1677622389
transform 1 0 1812 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1677622389
transform 1 0 1828 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4324
timestamp 1677622389
transform 1 0 1780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1677622389
transform 1 0 1828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1677622389
transform 1 0 1748 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3931
timestamp 1677622389
transform 1 0 1780 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4326
timestamp 1677622389
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3901
timestamp 1677622389
transform 1 0 1836 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1677622389
transform 1 0 1852 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1677622389
transform 1 0 1844 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4327
timestamp 1677622389
transform 1 0 1876 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3958
timestamp 1677622389
transform 1 0 1876 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1677622389
transform 1 0 1932 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1677622389
transform 1 0 1924 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1677622389
transform 1 0 1908 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4328
timestamp 1677622389
transform 1 0 1916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1677622389
transform 1 0 1932 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1677622389
transform 1 0 1940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1677622389
transform 1 0 1900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1677622389
transform 1 0 1908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1677622389
transform 1 0 1924 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3959
timestamp 1677622389
transform 1 0 1900 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1677622389
transform 1 0 1940 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4331
timestamp 1677622389
transform 1 0 1972 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3842
timestamp 1677622389
transform 1 0 1996 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4432
timestamp 1677622389
transform 1 0 1988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1677622389
transform 1 0 1996 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1677622389
transform 1 0 2036 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3881
timestamp 1677622389
transform 1 0 2044 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4333
timestamp 1677622389
transform 1 0 2052 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3903
timestamp 1677622389
transform 1 0 2036 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4434
timestamp 1677622389
transform 1 0 2044 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3783
timestamp 1677622389
transform 1 0 2076 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1677622389
transform 1 0 2108 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4435
timestamp 1677622389
transform 1 0 2116 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3933
timestamp 1677622389
transform 1 0 2116 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4436
timestamp 1677622389
transform 1 0 2124 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3800
timestamp 1677622389
transform 1 0 2140 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4437
timestamp 1677622389
transform 1 0 2164 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3934
timestamp 1677622389
transform 1 0 2156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1677622389
transform 1 0 2220 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4334
timestamp 1677622389
transform 1 0 2212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1677622389
transform 1 0 2220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1677622389
transform 1 0 2236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1677622389
transform 1 0 2252 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3814
timestamp 1677622389
transform 1 0 2268 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4338
timestamp 1677622389
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3845
timestamp 1677622389
transform 1 0 2316 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4438
timestamp 1677622389
transform 1 0 2308 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3846
timestamp 1677622389
transform 1 0 2348 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4339
timestamp 1677622389
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1677622389
transform 1 0 2332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1677622389
transform 1 0 2340 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1677622389
transform 1 0 2372 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3904
timestamp 1677622389
transform 1 0 2380 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1677622389
transform 1 0 2420 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4341
timestamp 1677622389
transform 1 0 2412 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3905
timestamp 1677622389
transform 1 0 2404 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4342
timestamp 1677622389
transform 1 0 2452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1677622389
transform 1 0 2468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1677622389
transform 1 0 2444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1677622389
transform 1 0 2460 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3906
timestamp 1677622389
transform 1 0 2468 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4443
timestamp 1677622389
transform 1 0 2476 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3960
timestamp 1677622389
transform 1 0 2460 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1677622389
transform 1 0 2532 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4344
timestamp 1677622389
transform 1 0 2532 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3785
timestamp 1677622389
transform 1 0 2556 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4345
timestamp 1677622389
transform 1 0 2572 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3882
timestamp 1677622389
transform 1 0 2692 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1677622389
transform 1 0 2780 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4346
timestamp 1677622389
transform 1 0 2716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1677622389
transform 1 0 2772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1677622389
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1677622389
transform 1 0 2692 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3935
timestamp 1677622389
transform 1 0 2740 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1677622389
transform 1 0 2756 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4445
timestamp 1677622389
transform 1 0 2804 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3936
timestamp 1677622389
transform 1 0 2804 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4279
timestamp 1677622389
transform 1 0 2844 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1677622389
transform 1 0 2828 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3907
timestamp 1677622389
transform 1 0 2836 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4492
timestamp 1677622389
transform 1 0 2836 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3937
timestamp 1677622389
transform 1 0 2844 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1677622389
transform 1 0 2876 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4447
timestamp 1677622389
transform 1 0 2876 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1677622389
transform 1 0 2884 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3908
timestamp 1677622389
transform 1 0 2892 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1677622389
transform 1 0 2884 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4349
timestamp 1677622389
transform 1 0 2908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1677622389
transform 1 0 2924 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3962
timestamp 1677622389
transform 1 0 2916 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4350
timestamp 1677622389
transform 1 0 2956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1677622389
transform 1 0 2972 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3939
timestamp 1677622389
transform 1 0 2972 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1677622389
transform 1 0 2988 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1677622389
transform 1 0 3036 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4351
timestamp 1677622389
transform 1 0 3036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1677622389
transform 1 0 2988 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3909
timestamp 1677622389
transform 1 0 3036 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1677622389
transform 1 0 3084 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1677622389
transform 1 0 3092 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1677622389
transform 1 0 3124 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1677622389
transform 1 0 3188 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1677622389
transform 1 0 3228 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4352
timestamp 1677622389
transform 1 0 3108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1677622389
transform 1 0 3148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1677622389
transform 1 0 3204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1677622389
transform 1 0 3220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1677622389
transform 1 0 3124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1677622389
transform 1 0 3212 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3941
timestamp 1677622389
transform 1 0 3108 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1677622389
transform 1 0 3124 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1677622389
transform 1 0 3172 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4453
timestamp 1677622389
transform 1 0 3228 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3789
timestamp 1677622389
transform 1 0 3252 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1677622389
transform 1 0 3268 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4356
timestamp 1677622389
transform 1 0 3252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1677622389
transform 1 0 3300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1677622389
transform 1 0 3268 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3910
timestamp 1677622389
transform 1 0 3348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1677622389
transform 1 0 3252 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1677622389
transform 1 0 3284 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1677622389
transform 1 0 3380 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4281
timestamp 1677622389
transform 1 0 3372 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3911
timestamp 1677622389
transform 1 0 3372 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4358
timestamp 1677622389
transform 1 0 3396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1677622389
transform 1 0 3412 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3850
timestamp 1677622389
transform 1 0 3420 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4359
timestamp 1677622389
transform 1 0 3420 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3912
timestamp 1677622389
transform 1 0 3420 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1677622389
transform 1 0 3412 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1677622389
transform 1 0 3444 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4455
timestamp 1677622389
transform 1 0 3444 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3946
timestamp 1677622389
transform 1 0 3444 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4282
timestamp 1677622389
transform 1 0 3460 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3883
timestamp 1677622389
transform 1 0 3460 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1677622389
transform 1 0 3476 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1677622389
transform 1 0 3500 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4360
timestamp 1677622389
transform 1 0 3484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1677622389
transform 1 0 3500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1677622389
transform 1 0 3492 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3913
timestamp 1677622389
transform 1 0 3508 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1677622389
transform 1 0 3524 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1677622389
transform 1 0 3524 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1677622389
transform 1 0 3532 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4457
timestamp 1677622389
transform 1 0 3524 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3853
timestamp 1677622389
transform 1 0 3548 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4362
timestamp 1677622389
transform 1 0 3572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1677622389
transform 1 0 3628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1677622389
transform 1 0 3548 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3914
timestamp 1677622389
transform 1 0 3572 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1677622389
transform 1 0 3548 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1677622389
transform 1 0 3572 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1677622389
transform 1 0 3588 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4364
timestamp 1677622389
transform 1 0 3668 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3819
timestamp 1677622389
transform 1 0 3724 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1677622389
transform 1 0 3700 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4365
timestamp 1677622389
transform 1 0 3692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1677622389
transform 1 0 3708 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3884
timestamp 1677622389
transform 1 0 3716 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4367
timestamp 1677622389
transform 1 0 3724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1677622389
transform 1 0 3700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3793
timestamp 1677622389
transform 1 0 3772 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1677622389
transform 1 0 3796 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1677622389
transform 1 0 3772 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4368
timestamp 1677622389
transform 1 0 3780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1677622389
transform 1 0 3796 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1677622389
transform 1 0 3764 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1677622389
transform 1 0 3772 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1677622389
transform 1 0 3788 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3947
timestamp 1677622389
transform 1 0 3764 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1677622389
transform 1 0 3796 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4370
timestamp 1677622389
transform 1 0 3812 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3948
timestamp 1677622389
transform 1 0 3812 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4371
timestamp 1677622389
transform 1 0 3860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1677622389
transform 1 0 3852 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3915
timestamp 1677622389
transform 1 0 3860 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1677622389
transform 1 0 3876 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1677622389
transform 1 0 3900 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4372
timestamp 1677622389
transform 1 0 3892 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3886
timestamp 1677622389
transform 1 0 3908 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4373
timestamp 1677622389
transform 1 0 3916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1677622389
transform 1 0 3932 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1677622389
transform 1 0 3900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1677622389
transform 1 0 3908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1677622389
transform 1 0 3924 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3916
timestamp 1677622389
transform 1 0 3932 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1677622389
transform 1 0 3908 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1677622389
transform 1 0 3924 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1677622389
transform 1 0 3900 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1677622389
transform 1 0 3948 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4375
timestamp 1677622389
transform 1 0 3948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1677622389
transform 1 0 3956 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1677622389
transform 1 0 3996 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3887
timestamp 1677622389
transform 1 0 4044 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4468
timestamp 1677622389
transform 1 0 4044 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3952
timestamp 1677622389
transform 1 0 3996 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1677622389
transform 1 0 4004 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4273
timestamp 1677622389
transform 1 0 4060 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3803
timestamp 1677622389
transform 1 0 4076 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4283
timestamp 1677622389
transform 1 0 4068 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3828
timestamp 1677622389
transform 1 0 4084 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4274
timestamp 1677622389
transform 1 0 4092 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3820
timestamp 1677622389
transform 1 0 4108 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4469
timestamp 1677622389
transform 1 0 4108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1677622389
transform 1 0 4124 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3917
timestamp 1677622389
transform 1 0 4124 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1677622389
transform 1 0 4140 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4470
timestamp 1677622389
transform 1 0 4132 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1677622389
transform 1 0 4164 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3830
timestamp 1677622389
transform 1 0 4204 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1677622389
transform 1 0 4204 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4378
timestamp 1677622389
transform 1 0 4196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1677622389
transform 1 0 4204 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3804
timestamp 1677622389
transform 1 0 4220 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4379
timestamp 1677622389
transform 1 0 4244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1677622389
transform 1 0 4220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1677622389
transform 1 0 4236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1677622389
transform 1 0 4252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1677622389
transform 1 0 4260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1677622389
transform 1 0 4268 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3859
timestamp 1677622389
transform 1 0 4284 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4381
timestamp 1677622389
transform 1 0 4276 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3860
timestamp 1677622389
transform 1 0 4316 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4382
timestamp 1677622389
transform 1 0 4300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1677622389
transform 1 0 4316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1677622389
transform 1 0 4308 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3861
timestamp 1677622389
transform 1 0 4340 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1677622389
transform 1 0 4380 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1677622389
transform 1 0 4372 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1677622389
transform 1 0 4372 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4384
timestamp 1677622389
transform 1 0 4396 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3889
timestamp 1677622389
transform 1 0 4436 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4385
timestamp 1677622389
transform 1 0 4452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1677622389
transform 1 0 4460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1677622389
transform 1 0 4372 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3970
timestamp 1677622389
transform 1 0 4452 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4478
timestamp 1677622389
transform 1 0 4484 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3831
timestamp 1677622389
transform 1 0 4524 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4387
timestamp 1677622389
transform 1 0 4516 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3863
timestamp 1677622389
transform 1 0 4548 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4388
timestamp 1677622389
transform 1 0 4548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1677622389
transform 1 0 4524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1677622389
transform 1 0 4540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1677622389
transform 1 0 4564 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3953
timestamp 1677622389
transform 1 0 4556 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4482
timestamp 1677622389
transform 1 0 4588 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3806
timestamp 1677622389
transform 1 0 4620 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1677622389
transform 1 0 4612 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1677622389
transform 1 0 4604 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4483
timestamp 1677622389
transform 1 0 4604 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3891
timestamp 1677622389
transform 1 0 4628 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4389
timestamp 1677622389
transform 1 0 4636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1677622389
transform 1 0 4620 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1677622389
transform 1 0 4652 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3864
timestamp 1677622389
transform 1 0 4700 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4391
timestamp 1677622389
transform 1 0 4684 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3892
timestamp 1677622389
transform 1 0 4692 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4392
timestamp 1677622389
transform 1 0 4700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1677622389
transform 1 0 4676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1677622389
transform 1 0 4692 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3954
timestamp 1677622389
transform 1 0 4684 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4393
timestamp 1677622389
transform 1 0 4724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1677622389
transform 1 0 4716 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3955
timestamp 1677622389
transform 1 0 4724 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4488
timestamp 1677622389
transform 1 0 4780 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3918
timestamp 1677622389
transform 1 0 4804 0 1 2605
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_42
timestamp 1677622389
transform 1 0 48 0 1 2570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_290
timestamp 1677622389
transform 1 0 72 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_325
timestamp 1677622389
transform -1 0 184 0 1 2570
box -9 -3 26 105
use AOI22X1  AOI22X1_198
timestamp 1677622389
transform -1 0 224 0 1 2570
box -8 -3 46 105
use INVX2  INVX2_326
timestamp 1677622389
transform -1 0 240 0 1 2570
box -9 -3 26 105
use FILL  FILL_4886
timestamp 1677622389
transform 1 0 240 0 1 2570
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1677622389
transform 1 0 248 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_200
timestamp 1677622389
transform 1 0 256 0 1 2570
box -8 -3 46 105
use M3_M2  M3_M2_3971
timestamp 1677622389
transform 1 0 308 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_193
timestamp 1677622389
transform -1 0 336 0 1 2570
box -8 -3 46 105
use FILL  FILL_4904
timestamp 1677622389
transform 1 0 336 0 1 2570
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1677622389
transform 1 0 344 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_291
timestamp 1677622389
transform 1 0 352 0 1 2570
box -8 -3 104 105
use FILL  FILL_4906
timestamp 1677622389
transform 1 0 448 0 1 2570
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1677622389
transform 1 0 456 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_202
timestamp 1677622389
transform 1 0 464 0 1 2570
box -8 -3 46 105
use M3_M2  M3_M2_3972
timestamp 1677622389
transform 1 0 516 0 1 2575
box -3 -3 3 3
use FILL  FILL_4923
timestamp 1677622389
transform 1 0 504 0 1 2570
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1677622389
transform 1 0 512 0 1 2570
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1677622389
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1677622389
transform 1 0 528 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_194
timestamp 1677622389
transform 1 0 536 0 1 2570
box -8 -3 46 105
use FILL  FILL_4934
timestamp 1677622389
transform 1 0 576 0 1 2570
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1677622389
transform 1 0 584 0 1 2570
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1677622389
transform 1 0 592 0 1 2570
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1677622389
transform 1 0 600 0 1 2570
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1677622389
transform 1 0 608 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_332
timestamp 1677622389
transform -1 0 632 0 1 2570
box -9 -3 26 105
use FILL  FILL_4948
timestamp 1677622389
transform 1 0 632 0 1 2570
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1677622389
transform 1 0 640 0 1 2570
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1677622389
transform 1 0 648 0 1 2570
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1677622389
transform 1 0 656 0 1 2570
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1677622389
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1677622389
transform 1 0 672 0 1 2570
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1677622389
transform 1 0 680 0 1 2570
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1677622389
transform 1 0 688 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_333
timestamp 1677622389
transform 1 0 696 0 1 2570
box -9 -3 26 105
use FILL  FILL_4956
timestamp 1677622389
transform 1 0 712 0 1 2570
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1677622389
transform 1 0 720 0 1 2570
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1677622389
transform 1 0 728 0 1 2570
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1677622389
transform 1 0 736 0 1 2570
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1677622389
transform 1 0 744 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_99
timestamp 1677622389
transform 1 0 752 0 1 2570
box -8 -3 34 105
use FILL  FILL_4967
timestamp 1677622389
transform 1 0 784 0 1 2570
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1677622389
transform 1 0 792 0 1 2570
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1677622389
transform 1 0 800 0 1 2570
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1677622389
transform 1 0 808 0 1 2570
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1677622389
transform 1 0 816 0 1 2570
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1677622389
transform 1 0 824 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_48
timestamp 1677622389
transform 1 0 832 0 1 2570
box -8 -3 32 105
use FILL  FILL_4978
timestamp 1677622389
transform 1 0 856 0 1 2570
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1677622389
transform 1 0 864 0 1 2570
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1677622389
transform 1 0 872 0 1 2570
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1677622389
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1677622389
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1677622389
transform 1 0 896 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_204
timestamp 1677622389
transform 1 0 904 0 1 2570
box -8 -3 46 105
use FILL  FILL_4991
timestamp 1677622389
transform 1 0 944 0 1 2570
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1677622389
transform 1 0 952 0 1 2570
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1677622389
transform 1 0 960 0 1 2570
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1677622389
transform 1 0 968 0 1 2570
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1677622389
transform 1 0 976 0 1 2570
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1677622389
transform 1 0 984 0 1 2570
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1677622389
transform 1 0 992 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_50
timestamp 1677622389
transform 1 0 1000 0 1 2570
box -8 -3 32 105
use FILL  FILL_5003
timestamp 1677622389
transform 1 0 1024 0 1 2570
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1677622389
transform 1 0 1032 0 1 2570
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1677622389
transform 1 0 1040 0 1 2570
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1677622389
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1677622389
transform 1 0 1056 0 1 2570
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1677622389
transform 1 0 1064 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_101
timestamp 1677622389
transform 1 0 1072 0 1 2570
box -8 -3 34 105
use FILL  FILL_5017
timestamp 1677622389
transform 1 0 1104 0 1 2570
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1677622389
transform 1 0 1112 0 1 2570
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1677622389
transform 1 0 1120 0 1 2570
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1677622389
transform 1 0 1128 0 1 2570
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1677622389
transform 1 0 1136 0 1 2570
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1677622389
transform 1 0 1144 0 1 2570
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1677622389
transform 1 0 1152 0 1 2570
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1677622389
transform 1 0 1160 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_102
timestamp 1677622389
transform -1 0 1200 0 1 2570
box -8 -3 34 105
use FILL  FILL_5032
timestamp 1677622389
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1677622389
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1677622389
transform 1 0 1216 0 1 2570
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1677622389
transform 1 0 1224 0 1 2570
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1677622389
transform 1 0 1232 0 1 2570
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1677622389
transform 1 0 1240 0 1 2570
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1677622389
transform 1 0 1248 0 1 2570
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1677622389
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1677622389
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1677622389
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_103
timestamp 1677622389
transform -1 0 1312 0 1 2570
box -8 -3 34 105
use FILL  FILL_5052
timestamp 1677622389
transform 1 0 1312 0 1 2570
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1677622389
transform 1 0 1320 0 1 2570
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1677622389
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1677622389
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1677622389
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1677622389
transform 1 0 1352 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_335
timestamp 1677622389
transform -1 0 1376 0 1 2570
box -9 -3 26 105
use FILL  FILL_5062
timestamp 1677622389
transform 1 0 1376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1677622389
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1677622389
transform 1 0 1392 0 1 2570
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1677622389
transform 1 0 1400 0 1 2570
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1677622389
transform 1 0 1408 0 1 2570
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1677622389
transform 1 0 1416 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_293
timestamp 1677622389
transform 1 0 1424 0 1 2570
box -8 -3 104 105
use FILL  FILL_5073
timestamp 1677622389
transform 1 0 1520 0 1 2570
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1677622389
transform 1 0 1528 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_337
timestamp 1677622389
transform 1 0 1536 0 1 2570
box -9 -3 26 105
use FILL  FILL_5084
timestamp 1677622389
transform 1 0 1552 0 1 2570
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1677622389
transform 1 0 1560 0 1 2570
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1677622389
transform 1 0 1568 0 1 2570
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1677622389
transform 1 0 1576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1677622389
transform 1 0 1584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1677622389
transform 1 0 1592 0 1 2570
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1677622389
transform 1 0 1600 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_339
timestamp 1677622389
transform -1 0 1624 0 1 2570
box -9 -3 26 105
use FILL  FILL_5097
timestamp 1677622389
transform 1 0 1624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1677622389
transform 1 0 1632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1677622389
transform 1 0 1640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1677622389
transform 1 0 1648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1677622389
transform 1 0 1656 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_196
timestamp 1677622389
transform -1 0 1704 0 1 2570
box -8 -3 46 105
use FILL  FILL_5102
timestamp 1677622389
transform 1 0 1704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1677622389
transform 1 0 1712 0 1 2570
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1677622389
transform 1 0 1720 0 1 2570
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1677622389
transform 1 0 1728 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3973
timestamp 1677622389
transform 1 0 1836 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_295
timestamp 1677622389
transform 1 0 1736 0 1 2570
box -8 -3 104 105
use FILL  FILL_5111
timestamp 1677622389
transform 1 0 1832 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3974
timestamp 1677622389
transform 1 0 1852 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_340
timestamp 1677622389
transform -1 0 1856 0 1 2570
box -9 -3 26 105
use FILL  FILL_5112
timestamp 1677622389
transform 1 0 1856 0 1 2570
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1677622389
transform 1 0 1864 0 1 2570
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1677622389
transform 1 0 1872 0 1 2570
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1677622389
transform 1 0 1880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1677622389
transform 1 0 1888 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_207
timestamp 1677622389
transform -1 0 1936 0 1 2570
box -8 -3 46 105
use FILL  FILL_5122
timestamp 1677622389
transform 1 0 1936 0 1 2570
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1677622389
transform 1 0 1944 0 1 2570
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1677622389
transform 1 0 1952 0 1 2570
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1677622389
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1677622389
transform 1 0 1968 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_343
timestamp 1677622389
transform -1 0 1992 0 1 2570
box -9 -3 26 105
use FILL  FILL_5133
timestamp 1677622389
transform 1 0 1992 0 1 2570
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1677622389
transform 1 0 2000 0 1 2570
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1677622389
transform 1 0 2008 0 1 2570
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1677622389
transform 1 0 2016 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_197
timestamp 1677622389
transform -1 0 2064 0 1 2570
box -8 -3 46 105
use FILL  FILL_5137
timestamp 1677622389
transform 1 0 2064 0 1 2570
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1677622389
transform 1 0 2072 0 1 2570
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1677622389
transform 1 0 2080 0 1 2570
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1677622389
transform 1 0 2088 0 1 2570
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1677622389
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1677622389
transform 1 0 2104 0 1 2570
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1677622389
transform 1 0 2112 0 1 2570
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1677622389
transform 1 0 2120 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_345
timestamp 1677622389
transform 1 0 2128 0 1 2570
box -9 -3 26 105
use FILL  FILL_5152
timestamp 1677622389
transform 1 0 2144 0 1 2570
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1677622389
transform 1 0 2152 0 1 2570
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1677622389
transform 1 0 2160 0 1 2570
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1677622389
transform 1 0 2168 0 1 2570
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1677622389
transform 1 0 2176 0 1 2570
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1677622389
transform 1 0 2184 0 1 2570
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1677622389
transform 1 0 2192 0 1 2570
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1677622389
transform 1 0 2200 0 1 2570
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1677622389
transform 1 0 2208 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_208
timestamp 1677622389
transform 1 0 2216 0 1 2570
box -8 -3 46 105
use FILL  FILL_5162
timestamp 1677622389
transform 1 0 2256 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3975
timestamp 1677622389
transform 1 0 2276 0 1 2575
box -3 -3 3 3
use FILL  FILL_5163
timestamp 1677622389
transform 1 0 2264 0 1 2570
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1677622389
transform 1 0 2272 0 1 2570
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1677622389
transform 1 0 2280 0 1 2570
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1677622389
transform 1 0 2288 0 1 2570
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1677622389
transform 1 0 2296 0 1 2570
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1677622389
transform 1 0 2304 0 1 2570
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1677622389
transform 1 0 2312 0 1 2570
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1677622389
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3976
timestamp 1677622389
transform 1 0 2364 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_209
timestamp 1677622389
transform 1 0 2328 0 1 2570
box -8 -3 46 105
use FILL  FILL_5174
timestamp 1677622389
transform 1 0 2368 0 1 2570
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1677622389
transform 1 0 2376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1677622389
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1677622389
transform 1 0 2392 0 1 2570
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1677622389
transform 1 0 2400 0 1 2570
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1677622389
transform 1 0 2408 0 1 2570
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1677622389
transform 1 0 2416 0 1 2570
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1677622389
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1677622389
transform 1 0 2432 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_198
timestamp 1677622389
transform -1 0 2480 0 1 2570
box -8 -3 46 105
use FILL  FILL_5188
timestamp 1677622389
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1677622389
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1677622389
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1677622389
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1677622389
transform 1 0 2512 0 1 2570
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1677622389
transform 1 0 2520 0 1 2570
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1677622389
transform 1 0 2528 0 1 2570
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1677622389
transform 1 0 2536 0 1 2570
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1677622389
transform 1 0 2544 0 1 2570
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1677622389
transform 1 0 2552 0 1 2570
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1677622389
transform 1 0 2560 0 1 2570
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1677622389
transform 1 0 2568 0 1 2570
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1677622389
transform 1 0 2576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1677622389
transform 1 0 2584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1677622389
transform 1 0 2592 0 1 2570
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1677622389
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1677622389
transform 1 0 2608 0 1 2570
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1677622389
transform 1 0 2616 0 1 2570
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1677622389
transform 1 0 2624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1677622389
transform 1 0 2632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1677622389
transform 1 0 2640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1677622389
transform 1 0 2648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1677622389
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1677622389
transform 1 0 2664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1677622389
transform 1 0 2672 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_300
timestamp 1677622389
transform 1 0 2680 0 1 2570
box -8 -3 104 105
use FILL  FILL_5230
timestamp 1677622389
transform 1 0 2776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1677622389
transform 1 0 2784 0 1 2570
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1677622389
transform 1 0 2792 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_104
timestamp 1677622389
transform 1 0 2800 0 1 2570
box -8 -3 34 105
use FILL  FILL_5236
timestamp 1677622389
transform 1 0 2832 0 1 2570
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1677622389
transform 1 0 2840 0 1 2570
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1677622389
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1677622389
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_52
timestamp 1677622389
transform 1 0 2864 0 1 2570
box -8 -3 32 105
use FILL  FILL_5244
timestamp 1677622389
transform 1 0 2888 0 1 2570
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1677622389
transform 1 0 2896 0 1 2570
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1677622389
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1677622389
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_106
timestamp 1677622389
transform -1 0 2952 0 1 2570
box -8 -3 34 105
use FILL  FILL_5252
timestamp 1677622389
transform 1 0 2952 0 1 2570
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1677622389
transform 1 0 2960 0 1 2570
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1677622389
transform 1 0 2968 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_302
timestamp 1677622389
transform 1 0 2976 0 1 2570
box -8 -3 104 105
use FILL  FILL_5255
timestamp 1677622389
transform 1 0 3072 0 1 2570
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1677622389
transform 1 0 3080 0 1 2570
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1677622389
transform 1 0 3088 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_348
timestamp 1677622389
transform 1 0 3096 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_303
timestamp 1677622389
transform 1 0 3112 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_349
timestamp 1677622389
transform 1 0 3208 0 1 2570
box -9 -3 26 105
use BUFX2  BUFX2_42
timestamp 1677622389
transform -1 0 3248 0 1 2570
box -5 -3 28 105
use FILL  FILL_5271
timestamp 1677622389
transform 1 0 3248 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_305
timestamp 1677622389
transform 1 0 3256 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_351
timestamp 1677622389
transform 1 0 3352 0 1 2570
box -9 -3 26 105
use FILL  FILL_5278
timestamp 1677622389
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1677622389
transform 1 0 3376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1677622389
transform 1 0 3384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1677622389
transform 1 0 3392 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_29
timestamp 1677622389
transform -1 0 3432 0 1 2570
box -8 -3 40 105
use FILL  FILL_5290
timestamp 1677622389
transform 1 0 3432 0 1 2570
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1677622389
transform 1 0 3440 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3977
timestamp 1677622389
transform 1 0 3460 0 1 2575
box -3 -3 3 3
use FILL  FILL_5292
timestamp 1677622389
transform 1 0 3448 0 1 2570
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1677622389
transform 1 0 3456 0 1 2570
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1677622389
transform 1 0 3464 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_201
timestamp 1677622389
transform 1 0 3472 0 1 2570
box -8 -3 46 105
use FILL  FILL_5299
timestamp 1677622389
transform 1 0 3512 0 1 2570
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1677622389
transform 1 0 3520 0 1 2570
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1677622389
transform 1 0 3528 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_306
timestamp 1677622389
transform 1 0 3536 0 1 2570
box -8 -3 104 105
use FILL  FILL_5305
timestamp 1677622389
transform 1 0 3632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1677622389
transform 1 0 3640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1677622389
transform 1 0 3648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1677622389
transform 1 0 3656 0 1 2570
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1677622389
transform 1 0 3664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1677622389
transform 1 0 3672 0 1 2570
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1677622389
transform 1 0 3680 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_211
timestamp 1677622389
transform -1 0 3728 0 1 2570
box -8 -3 46 105
use FILL  FILL_5326
timestamp 1677622389
transform 1 0 3728 0 1 2570
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1677622389
transform 1 0 3736 0 1 2570
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1677622389
transform 1 0 3744 0 1 2570
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1677622389
transform 1 0 3752 0 1 2570
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1677622389
transform 1 0 3760 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3978
timestamp 1677622389
transform 1 0 3804 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_203
timestamp 1677622389
transform 1 0 3768 0 1 2570
box -8 -3 46 105
use FILL  FILL_5336
timestamp 1677622389
transform 1 0 3808 0 1 2570
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1677622389
transform 1 0 3816 0 1 2570
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1677622389
transform 1 0 3824 0 1 2570
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1677622389
transform 1 0 3832 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3979
timestamp 1677622389
transform 1 0 3852 0 1 2575
box -3 -3 3 3
use FILL  FILL_5340
timestamp 1677622389
transform 1 0 3840 0 1 2570
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1677622389
transform 1 0 3848 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_354
timestamp 1677622389
transform -1 0 3872 0 1 2570
box -9 -3 26 105
use FILL  FILL_5342
timestamp 1677622389
transform 1 0 3872 0 1 2570
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1677622389
transform 1 0 3880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1677622389
transform 1 0 3888 0 1 2570
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1677622389
transform 1 0 3896 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_204
timestamp 1677622389
transform 1 0 3904 0 1 2570
box -8 -3 46 105
use FILL  FILL_5349
timestamp 1677622389
transform 1 0 3944 0 1 2570
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1677622389
transform 1 0 3952 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_308
timestamp 1677622389
transform -1 0 4056 0 1 2570
box -8 -3 104 105
use FILL  FILL_5351
timestamp 1677622389
transform 1 0 4056 0 1 2570
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1677622389
transform 1 0 4064 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_30
timestamp 1677622389
transform 1 0 4072 0 1 2570
box -8 -3 40 105
use FILL  FILL_5353
timestamp 1677622389
transform 1 0 4104 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3980
timestamp 1677622389
transform 1 0 4124 0 1 2575
box -3 -3 3 3
use FILL  FILL_5354
timestamp 1677622389
transform 1 0 4112 0 1 2570
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1677622389
transform 1 0 4120 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_50
timestamp 1677622389
transform -1 0 4152 0 1 2570
box -5 -3 28 105
use FILL  FILL_5356
timestamp 1677622389
transform 1 0 4152 0 1 2570
box -8 -3 16 105
use FILL  FILL_5357
timestamp 1677622389
transform 1 0 4160 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_51
timestamp 1677622389
transform 1 0 4168 0 1 2570
box -5 -3 28 105
use FILL  FILL_5358
timestamp 1677622389
transform 1 0 4192 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3981
timestamp 1677622389
transform 1 0 4212 0 1 2575
box -3 -3 3 3
use FILL  FILL_5367
timestamp 1677622389
transform 1 0 4200 0 1 2570
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1677622389
transform 1 0 4208 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3982
timestamp 1677622389
transform 1 0 4252 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_206
timestamp 1677622389
transform 1 0 4216 0 1 2570
box -8 -3 46 105
use FILL  FILL_5370
timestamp 1677622389
transform 1 0 4256 0 1 2570
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1677622389
transform 1 0 4264 0 1 2570
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1677622389
transform 1 0 4272 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_212
timestamp 1677622389
transform -1 0 4320 0 1 2570
box -8 -3 46 105
use M3_M2  M3_M2_3983
timestamp 1677622389
transform 1 0 4332 0 1 2575
box -3 -3 3 3
use FILL  FILL_5376
timestamp 1677622389
transform 1 0 4320 0 1 2570
box -8 -3 16 105
use FILL  FILL_5377
timestamp 1677622389
transform 1 0 4328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5378
timestamp 1677622389
transform 1 0 4336 0 1 2570
box -8 -3 16 105
use FILL  FILL_5383
timestamp 1677622389
transform 1 0 4344 0 1 2570
box -8 -3 16 105
use FILL  FILL_5385
timestamp 1677622389
transform 1 0 4352 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3984
timestamp 1677622389
transform 1 0 4428 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_311
timestamp 1677622389
transform 1 0 4360 0 1 2570
box -8 -3 104 105
use BUFX2  BUFX2_52
timestamp 1677622389
transform 1 0 4456 0 1 2570
box -5 -3 28 105
use FILL  FILL_5387
timestamp 1677622389
transform 1 0 4480 0 1 2570
box -8 -3 16 105
use FILL  FILL_5393
timestamp 1677622389
transform 1 0 4488 0 1 2570
box -8 -3 16 105
use FILL  FILL_5395
timestamp 1677622389
transform 1 0 4496 0 1 2570
box -8 -3 16 105
use FILL  FILL_5397
timestamp 1677622389
transform 1 0 4504 0 1 2570
box -8 -3 16 105
use FILL  FILL_5399
timestamp 1677622389
transform 1 0 4512 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3985
timestamp 1677622389
transform 1 0 4540 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_208
timestamp 1677622389
transform 1 0 4520 0 1 2570
box -8 -3 46 105
use FILL  FILL_5400
timestamp 1677622389
transform 1 0 4560 0 1 2570
box -8 -3 16 105
use FILL  FILL_5401
timestamp 1677622389
transform 1 0 4568 0 1 2570
box -8 -3 16 105
use FILL  FILL_5402
timestamp 1677622389
transform 1 0 4576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5403
timestamp 1677622389
transform 1 0 4584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5404
timestamp 1677622389
transform 1 0 4592 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3986
timestamp 1677622389
transform 1 0 4612 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_358
timestamp 1677622389
transform 1 0 4600 0 1 2570
box -9 -3 26 105
use FILL  FILL_5405
timestamp 1677622389
transform 1 0 4616 0 1 2570
box -8 -3 16 105
use FILL  FILL_5406
timestamp 1677622389
transform 1 0 4624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5407
timestamp 1677622389
transform 1 0 4632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5408
timestamp 1677622389
transform 1 0 4640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5409
timestamp 1677622389
transform 1 0 4648 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_209
timestamp 1677622389
transform 1 0 4656 0 1 2570
box -8 -3 46 105
use FILL  FILL_5410
timestamp 1677622389
transform 1 0 4696 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_359
timestamp 1677622389
transform -1 0 4720 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_360
timestamp 1677622389
transform -1 0 4736 0 1 2570
box -9 -3 26 105
use FILL  FILL_5411
timestamp 1677622389
transform 1 0 4736 0 1 2570
box -8 -3 16 105
use FILL  FILL_5412
timestamp 1677622389
transform 1 0 4744 0 1 2570
box -8 -3 16 105
use FILL  FILL_5413
timestamp 1677622389
transform 1 0 4752 0 1 2570
box -8 -3 16 105
use FILL  FILL_5414
timestamp 1677622389
transform 1 0 4760 0 1 2570
box -8 -3 16 105
use FILL  FILL_5415
timestamp 1677622389
transform 1 0 4768 0 1 2570
box -8 -3 16 105
use FILL  FILL_5416
timestamp 1677622389
transform 1 0 4776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5417
timestamp 1677622389
transform 1 0 4784 0 1 2570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_43
timestamp 1677622389
transform 1 0 4819 0 1 2570
box -10 -3 10 3
use M2_M1  M2_M1_4585
timestamp 1677622389
transform 1 0 116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1677622389
transform 1 0 164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1677622389
transform 1 0 172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1677622389
transform 1 0 196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1677622389
transform 1 0 156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1677622389
transform 1 0 180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1677622389
transform 1 0 212 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4037
timestamp 1677622389
transform 1 0 220 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4588
timestamp 1677622389
transform 1 0 244 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4111
timestamp 1677622389
transform 1 0 244 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4589
timestamp 1677622389
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3991
timestamp 1677622389
transform 1 0 316 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1677622389
transform 1 0 316 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1677622389
transform 1 0 332 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1677622389
transform 1 0 356 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4502
timestamp 1677622389
transform 1 0 316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1677622389
transform 1 0 324 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4038
timestamp 1677622389
transform 1 0 348 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4504
timestamp 1677622389
transform 1 0 356 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1677622389
transform 1 0 316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1677622389
transform 1 0 332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1677622389
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4081
timestamp 1677622389
transform 1 0 316 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1677622389
transform 1 0 348 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4593
timestamp 1677622389
transform 1 0 372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1677622389
transform 1 0 380 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4082
timestamp 1677622389
transform 1 0 380 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1677622389
transform 1 0 404 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1677622389
transform 1 0 412 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4505
timestamp 1677622389
transform 1 0 428 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4017
timestamp 1677622389
transform 1 0 444 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4506
timestamp 1677622389
transform 1 0 444 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4040
timestamp 1677622389
transform 1 0 452 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4595
timestamp 1677622389
transform 1 0 436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1677622389
transform 1 0 444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1677622389
transform 1 0 452 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4083
timestamp 1677622389
transform 1 0 428 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1677622389
transform 1 0 452 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1677622389
transform 1 0 468 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4507
timestamp 1677622389
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4018
timestamp 1677622389
transform 1 0 596 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1677622389
transform 1 0 644 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4508
timestamp 1677622389
transform 1 0 644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1677622389
transform 1 0 732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1677622389
transform 1 0 668 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1677622389
transform 1 0 724 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4141
timestamp 1677622389
transform 1 0 644 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4510
timestamp 1677622389
transform 1 0 748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1677622389
transform 1 0 748 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4113
timestamp 1677622389
transform 1 0 748 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1677622389
transform 1 0 796 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1677622389
transform 1 0 780 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1677622389
transform 1 0 796 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4601
timestamp 1677622389
transform 1 0 780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1677622389
transform 1 0 796 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4085
timestamp 1677622389
transform 1 0 780 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1677622389
transform 1 0 772 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1677622389
transform 1 0 828 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4511
timestamp 1677622389
transform 1 0 828 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4115
timestamp 1677622389
transform 1 0 820 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4512
timestamp 1677622389
transform 1 0 836 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4043
timestamp 1677622389
transform 1 0 844 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1677622389
transform 1 0 836 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4493
timestamp 1677622389
transform 1 0 860 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1677622389
transform 1 0 884 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4044
timestamp 1677622389
transform 1 0 900 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1677622389
transform 1 0 908 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1677622389
transform 1 0 972 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4513
timestamp 1677622389
transform 1 0 956 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4045
timestamp 1677622389
transform 1 0 964 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4514
timestamp 1677622389
transform 1 0 972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1677622389
transform 1 0 964 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4046
timestamp 1677622389
transform 1 0 988 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4515
timestamp 1677622389
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1677622389
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1677622389
transform 1 0 1012 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4116
timestamp 1677622389
transform 1 0 1020 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1677622389
transform 1 0 1012 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1677622389
transform 1 0 1060 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4685
timestamp 1677622389
transform 1 0 1060 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_3995
timestamp 1677622389
transform 1 0 1092 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4517
timestamp 1677622389
transform 1 0 1076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1677622389
transform 1 0 1084 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4066
timestamp 1677622389
transform 1 0 1092 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4518
timestamp 1677622389
transform 1 0 1108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1677622389
transform 1 0 1100 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4087
timestamp 1677622389
transform 1 0 1084 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1677622389
transform 1 0 1116 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4608
timestamp 1677622389
transform 1 0 1132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1677622389
transform 1 0 1196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1677622389
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1677622389
transform 1 0 1220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1677622389
transform 1 0 1204 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4089
timestamp 1677622389
transform 1 0 1204 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1677622389
transform 1 0 1236 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4610
timestamp 1677622389
transform 1 0 1252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1677622389
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1677622389
transform 1 0 1300 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4156
timestamp 1677622389
transform 1 0 1284 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4612
timestamp 1677622389
transform 1 0 1340 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3996
timestamp 1677622389
transform 1 0 1356 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4686
timestamp 1677622389
transform 1 0 1348 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4157
timestamp 1677622389
transform 1 0 1340 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4523
timestamp 1677622389
transform 1 0 1372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1677622389
transform 1 0 1428 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4142
timestamp 1677622389
transform 1 0 1468 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1677622389
transform 1 0 1492 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1677622389
transform 1 0 1532 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4525
timestamp 1677622389
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1677622389
transform 1 0 1508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1677622389
transform 1 0 1524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1677622389
transform 1 0 1532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1677622389
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4090
timestamp 1677622389
transform 1 0 1532 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1677622389
transform 1 0 1500 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1677622389
transform 1 0 1524 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4614
timestamp 1677622389
transform 1 0 1548 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4091
timestamp 1677622389
transform 1 0 1548 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1677622389
transform 1 0 1540 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1677622389
transform 1 0 1532 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1677622389
transform 1 0 1564 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1677622389
transform 1 0 1572 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4615
timestamp 1677622389
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1677622389
transform 1 0 1596 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4092
timestamp 1677622389
transform 1 0 1596 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1677622389
transform 1 0 1612 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1677622389
transform 1 0 1612 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4617
timestamp 1677622389
transform 1 0 1628 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3997
timestamp 1677622389
transform 1 0 1724 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1677622389
transform 1 0 1692 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4529
timestamp 1677622389
transform 1 0 1716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1677622389
transform 1 0 1684 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3998
timestamp 1677622389
transform 1 0 1780 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4530
timestamp 1677622389
transform 1 0 1756 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3999
timestamp 1677622389
transform 1 0 1852 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4531
timestamp 1677622389
transform 1 0 1844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1677622389
transform 1 0 1804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1677622389
transform 1 0 1836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1677622389
transform 1 0 1844 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4094
timestamp 1677622389
transform 1 0 1804 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1677622389
transform 1 0 1844 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1677622389
transform 1 0 1852 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4622
timestamp 1677622389
transform 1 0 1900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1677622389
transform 1 0 1908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1677622389
transform 1 0 1916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1677622389
transform 1 0 1956 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4119
timestamp 1677622389
transform 1 0 1956 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4623
timestamp 1677622389
transform 1 0 1980 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4096
timestamp 1677622389
transform 1 0 1980 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4535
timestamp 1677622389
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4052
timestamp 1677622389
transform 1 0 2020 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1677622389
transform 1 0 2076 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4624
timestamp 1677622389
transform 1 0 2020 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4097
timestamp 1677622389
transform 1 0 2020 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1677622389
transform 1 0 2060 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4625
timestamp 1677622389
transform 1 0 2084 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4121
timestamp 1677622389
transform 1 0 2084 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4626
timestamp 1677622389
transform 1 0 2100 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4023
timestamp 1677622389
transform 1 0 2140 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4536
timestamp 1677622389
transform 1 0 2140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1677622389
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4000
timestamp 1677622389
transform 1 0 2172 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1677622389
transform 1 0 2260 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1677622389
transform 1 0 2244 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4537
timestamp 1677622389
transform 1 0 2244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1677622389
transform 1 0 2260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1677622389
transform 1 0 2212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1677622389
transform 1 0 2276 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1677622389
transform 1 0 2268 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4098
timestamp 1677622389
transform 1 0 2268 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1677622389
transform 1 0 2252 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1677622389
transform 1 0 2276 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4698
timestamp 1677622389
transform 1 0 2276 0 1 2485
box -2 -2 2 2
use M3_M2  M3_M2_4002
timestamp 1677622389
transform 1 0 2348 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1677622389
transform 1 0 2300 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1677622389
transform 1 0 2332 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4539
timestamp 1677622389
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4003
timestamp 1677622389
transform 1 0 2388 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4540
timestamp 1677622389
transform 1 0 2388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1677622389
transform 1 0 2332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1677622389
transform 1 0 2380 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4099
timestamp 1677622389
transform 1 0 2332 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1677622389
transform 1 0 2316 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1677622389
transform 1 0 2388 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4632
timestamp 1677622389
transform 1 0 2404 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4123
timestamp 1677622389
transform 1 0 2420 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1677622389
transform 1 0 2444 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1677622389
transform 1 0 2476 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1677622389
transform 1 0 2468 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4541
timestamp 1677622389
transform 1 0 2444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1677622389
transform 1 0 2460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1677622389
transform 1 0 2452 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4124
timestamp 1677622389
transform 1 0 2444 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4634
timestamp 1677622389
transform 1 0 2468 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4005
timestamp 1677622389
transform 1 0 2564 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4543
timestamp 1677622389
transform 1 0 2548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1677622389
transform 1 0 2564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1677622389
transform 1 0 2572 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4067
timestamp 1677622389
transform 1 0 2540 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4635
timestamp 1677622389
transform 1 0 2556 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4068
timestamp 1677622389
transform 1 0 2564 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4636
timestamp 1677622389
transform 1 0 2572 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4100
timestamp 1677622389
transform 1 0 2548 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1677622389
transform 1 0 2596 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1677622389
transform 1 0 2588 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4637
timestamp 1677622389
transform 1 0 2612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1677622389
transform 1 0 2652 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4102
timestamp 1677622389
transform 1 0 2652 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4495
timestamp 1677622389
transform 1 0 2756 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1677622389
transform 1 0 2668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1677622389
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4069
timestamp 1677622389
transform 1 0 2740 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4547
timestamp 1677622389
transform 1 0 2764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1677622389
transform 1 0 2748 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4103
timestamp 1677622389
transform 1 0 2692 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4641
timestamp 1677622389
transform 1 0 2780 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4007
timestamp 1677622389
transform 1 0 2812 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4496
timestamp 1677622389
transform 1 0 2820 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1677622389
transform 1 0 2828 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3988
timestamp 1677622389
transform 1 0 2876 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4497
timestamp 1677622389
transform 1 0 2876 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1677622389
transform 1 0 2892 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4070
timestamp 1677622389
transform 1 0 2892 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4687
timestamp 1677622389
transform 1 0 2892 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4125
timestamp 1677622389
transform 1 0 2892 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4550
timestamp 1677622389
transform 1 0 2916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1677622389
transform 1 0 2924 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4071
timestamp 1677622389
transform 1 0 2908 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4642
timestamp 1677622389
transform 1 0 2916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1677622389
transform 1 0 2932 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4126
timestamp 1677622389
transform 1 0 2924 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4689
timestamp 1677622389
transform 1 0 2956 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1677622389
transform 1 0 2980 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4072
timestamp 1677622389
transform 1 0 3020 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1677622389
transform 1 0 3036 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1677622389
transform 1 0 3068 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4552
timestamp 1677622389
transform 1 0 3036 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1677622389
transform 1 0 3044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1677622389
transform 1 0 3060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1677622389
transform 1 0 3076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1677622389
transform 1 0 3052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1677622389
transform 1 0 3068 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4127
timestamp 1677622389
transform 1 0 3060 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1677622389
transform 1 0 3068 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1677622389
transform 1 0 3092 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4556
timestamp 1677622389
transform 1 0 3108 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4008
timestamp 1677622389
transform 1 0 3212 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4557
timestamp 1677622389
transform 1 0 3132 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4073
timestamp 1677622389
transform 1 0 3132 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4646
timestamp 1677622389
transform 1 0 3156 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4074
timestamp 1677622389
transform 1 0 3196 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1677622389
transform 1 0 3156 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1677622389
transform 1 0 3236 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4647
timestamp 1677622389
transform 1 0 3244 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4129
timestamp 1677622389
transform 1 0 3252 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1677622389
transform 1 0 3244 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4648
timestamp 1677622389
transform 1 0 3268 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4030
timestamp 1677622389
transform 1 0 3284 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4558
timestamp 1677622389
transform 1 0 3284 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4130
timestamp 1677622389
transform 1 0 3276 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4649
timestamp 1677622389
transform 1 0 3292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1677622389
transform 1 0 3356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4131
timestamp 1677622389
transform 1 0 3364 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4559
timestamp 1677622389
transform 1 0 3380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1677622389
transform 1 0 3380 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4055
timestamp 1677622389
transform 1 0 3396 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1677622389
transform 1 0 3420 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4560
timestamp 1677622389
transform 1 0 3420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1677622389
transform 1 0 3404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1677622389
transform 1 0 3428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1677622389
transform 1 0 3460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1677622389
transform 1 0 3460 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4105
timestamp 1677622389
transform 1 0 3460 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1677622389
transform 1 0 3452 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4562
timestamp 1677622389
transform 1 0 3508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1677622389
transform 1 0 3524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1677622389
transform 1 0 3484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1677622389
transform 1 0 3492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1677622389
transform 1 0 3516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1677622389
transform 1 0 3532 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4075
timestamp 1677622389
transform 1 0 3564 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1677622389
transform 1 0 3556 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4564
timestamp 1677622389
transform 1 0 3628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1677622389
transform 1 0 3636 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4076
timestamp 1677622389
transform 1 0 3636 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1677622389
transform 1 0 3652 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1677622389
transform 1 0 3676 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4659
timestamp 1677622389
transform 1 0 3668 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1677622389
transform 1 0 3676 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4032
timestamp 1677622389
transform 1 0 3724 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4566
timestamp 1677622389
transform 1 0 3716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1677622389
transform 1 0 3740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1677622389
transform 1 0 3724 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4077
timestamp 1677622389
transform 1 0 3740 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1677622389
transform 1 0 3788 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1677622389
transform 1 0 3820 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1677622389
transform 1 0 3796 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1677622389
transform 1 0 3828 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4568
timestamp 1677622389
transform 1 0 3796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1677622389
transform 1 0 3820 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4056
timestamp 1677622389
transform 1 0 3884 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4663
timestamp 1677622389
transform 1 0 3900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1677622389
transform 1 0 3924 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4078
timestamp 1677622389
transform 1 0 3924 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4664
timestamp 1677622389
transform 1 0 3948 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4079
timestamp 1677622389
transform 1 0 3988 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4665
timestamp 1677622389
transform 1 0 4004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1677622389
transform 1 0 4012 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4057
timestamp 1677622389
transform 1 0 4084 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4570
timestamp 1677622389
transform 1 0 4108 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4080
timestamp 1677622389
transform 1 0 4044 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4667
timestamp 1677622389
transform 1 0 4084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1677622389
transform 1 0 4124 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4058
timestamp 1677622389
transform 1 0 4148 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4572
timestamp 1677622389
transform 1 0 4156 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4059
timestamp 1677622389
transform 1 0 4164 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4573
timestamp 1677622389
transform 1 0 4172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1677622389
transform 1 0 4148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1677622389
transform 1 0 4180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1677622389
transform 1 0 4196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1677622389
transform 1 0 4188 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4134
timestamp 1677622389
transform 1 0 4196 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4691
timestamp 1677622389
transform 1 0 4244 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1677622389
transform 1 0 4228 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_4159
timestamp 1677622389
transform 1 0 4236 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4671
timestamp 1677622389
transform 1 0 4292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1677622389
transform 1 0 4300 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1677622389
transform 1 0 4284 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_4150
timestamp 1677622389
transform 1 0 4292 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1677622389
transform 1 0 4324 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4574
timestamp 1677622389
transform 1 0 4324 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4107
timestamp 1677622389
transform 1 0 4316 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4672
timestamp 1677622389
transform 1 0 4340 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4135
timestamp 1677622389
transform 1 0 4332 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4575
timestamp 1677622389
transform 1 0 4348 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4060
timestamp 1677622389
transform 1 0 4356 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1677622389
transform 1 0 4348 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1677622389
transform 1 0 4396 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4576
timestamp 1677622389
transform 1 0 4380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1677622389
transform 1 0 4396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1677622389
transform 1 0 4372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1677622389
transform 1 0 4388 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4061
timestamp 1677622389
transform 1 0 4412 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4675
timestamp 1677622389
transform 1 0 4404 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4137
timestamp 1677622389
transform 1 0 4396 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4676
timestamp 1677622389
transform 1 0 4420 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4108
timestamp 1677622389
transform 1 0 4412 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4693
timestamp 1677622389
transform 1 0 4436 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4138
timestamp 1677622389
transform 1 0 4436 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4578
timestamp 1677622389
transform 1 0 4444 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4012
timestamp 1677622389
transform 1 0 4460 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4677
timestamp 1677622389
transform 1 0 4460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1677622389
transform 1 0 4452 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1677622389
transform 1 0 4484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1677622389
transform 1 0 4476 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1677622389
transform 1 0 4524 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4062
timestamp 1677622389
transform 1 0 4548 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4581
timestamp 1677622389
transform 1 0 4556 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4063
timestamp 1677622389
transform 1 0 4564 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4582
timestamp 1677622389
transform 1 0 4572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1677622389
transform 1 0 4588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1677622389
transform 1 0 4532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1677622389
transform 1 0 4548 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4109
timestamp 1677622389
transform 1 0 4524 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1677622389
transform 1 0 4532 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4680
timestamp 1677622389
transform 1 0 4564 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4110
timestamp 1677622389
transform 1 0 4564 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4681
timestamp 1677622389
transform 1 0 4612 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4139
timestamp 1677622389
transform 1 0 4580 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1677622389
transform 1 0 4684 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1677622389
transform 1 0 4676 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1677622389
transform 1 0 4588 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1677622389
transform 1 0 4668 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4682
timestamp 1677622389
transform 1 0 4684 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4036
timestamp 1677622389
transform 1 0 4716 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4584
timestamp 1677622389
transform 1 0 4700 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4065
timestamp 1677622389
transform 1 0 4724 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4683
timestamp 1677622389
transform 1 0 4724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1677622389
transform 1 0 4780 0 1 2525
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_44
timestamp 1677622389
transform 1 0 24 0 1 2470
box -10 -3 10 3
use FILL  FILL_4887
timestamp 1677622389
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1677622389
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1677622389
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1677622389
transform 1 0 96 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1677622389
transform 1 0 104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1677622389
transform 1 0 112 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_327
timestamp 1677622389
transform -1 0 136 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4893
timestamp 1677622389
transform 1 0 136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1677622389
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1677622389
transform 1 0 152 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_199
timestamp 1677622389
transform -1 0 200 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4896
timestamp 1677622389
transform 1 0 200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1677622389
transform 1 0 208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1677622389
transform 1 0 216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1677622389
transform 1 0 224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1677622389
transform 1 0 232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1677622389
transform 1 0 240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1677622389
transform 1 0 248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1677622389
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1677622389
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_328
timestamp 1677622389
transform -1 0 288 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4909
timestamp 1677622389
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1677622389
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1677622389
transform 1 0 304 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_201
timestamp 1677622389
transform -1 0 352 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4912
timestamp 1677622389
transform 1 0 352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1677622389
transform 1 0 360 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_329
timestamp 1677622389
transform -1 0 384 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4914
timestamp 1677622389
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1677622389
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1677622389
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1677622389
transform 1 0 408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1677622389
transform 1 0 416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1677622389
transform 1 0 424 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_330
timestamp 1677622389
transform -1 0 448 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4920
timestamp 1677622389
transform 1 0 448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1677622389
transform 1 0 456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1677622389
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_331
timestamp 1677622389
transform -1 0 488 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4925
timestamp 1677622389
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1677622389
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1677622389
transform 1 0 504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1677622389
transform 1 0 512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1677622389
transform 1 0 520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1677622389
transform 1 0 528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1677622389
transform 1 0 536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1677622389
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1677622389
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1677622389
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4160
timestamp 1677622389
transform 1 0 580 0 1 2475
box -3 -3 3 3
use FILL  FILL_4939
timestamp 1677622389
transform 1 0 568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1677622389
transform 1 0 576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1677622389
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1677622389
transform 1 0 592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1677622389
transform 1 0 600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1677622389
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1677622389
transform 1 0 616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1677622389
transform 1 0 624 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1677622389
transform 1 0 632 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4962
timestamp 1677622389
transform 1 0 728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1677622389
transform 1 0 736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1677622389
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1677622389
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_203
timestamp 1677622389
transform 1 0 760 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4971
timestamp 1677622389
transform 1 0 800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1677622389
transform 1 0 808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1677622389
transform 1 0 816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1677622389
transform 1 0 824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1677622389
transform 1 0 832 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4161
timestamp 1677622389
transform 1 0 860 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_334
timestamp 1677622389
transform 1 0 840 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4980
timestamp 1677622389
transform 1 0 856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1677622389
transform 1 0 864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1677622389
transform 1 0 872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1677622389
transform 1 0 880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1677622389
transform 1 0 888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1677622389
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_49
timestamp 1677622389
transform 1 0 904 0 -1 2570
box -8 -3 32 105
use FILL  FILL_4992
timestamp 1677622389
transform 1 0 928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1677622389
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1677622389
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1677622389
transform 1 0 952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1677622389
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_100
timestamp 1677622389
transform 1 0 968 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5004
timestamp 1677622389
transform 1 0 1000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1677622389
transform 1 0 1008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1677622389
transform 1 0 1016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1677622389
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1677622389
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1677622389
transform 1 0 1040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1677622389
transform 1 0 1048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1677622389
transform 1 0 1056 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_205
timestamp 1677622389
transform 1 0 1064 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5018
timestamp 1677622389
transform 1 0 1104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1677622389
transform 1 0 1112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1677622389
transform 1 0 1120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1677622389
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1677622389
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1677622389
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1677622389
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1677622389
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1677622389
transform 1 0 1168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1677622389
transform 1 0 1176 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_206
timestamp 1677622389
transform 1 0 1184 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5039
timestamp 1677622389
transform 1 0 1224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1677622389
transform 1 0 1232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1677622389
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1677622389
transform 1 0 1248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1677622389
transform 1 0 1256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1677622389
transform 1 0 1264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1677622389
transform 1 0 1272 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1677622389
transform -1 0 1312 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5053
timestamp 1677622389
transform 1 0 1312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1677622389
transform 1 0 1320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1677622389
transform 1 0 1328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1677622389
transform 1 0 1336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1677622389
transform 1 0 1344 0 -1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1677622389
transform -1 0 1376 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5064
timestamp 1677622389
transform 1 0 1376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1677622389
transform 1 0 1384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1677622389
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1677622389
transform 1 0 1400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1677622389
transform 1 0 1408 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_336
timestamp 1677622389
transform -1 0 1432 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5076
timestamp 1677622389
transform 1 0 1432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1677622389
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1677622389
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1677622389
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1677622389
transform 1 0 1464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1677622389
transform 1 0 1472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1677622389
transform 1 0 1480 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_195
timestamp 1677622389
transform -1 0 1528 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5083
timestamp 1677622389
transform 1 0 1528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1677622389
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1677622389
transform 1 0 1544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1677622389
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1677622389
transform 1 0 1560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1677622389
transform 1 0 1568 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_338
timestamp 1677622389
transform 1 0 1576 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5095
timestamp 1677622389
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1677622389
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1677622389
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1677622389
transform 1 0 1616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1677622389
transform 1 0 1624 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_294
timestamp 1677622389
transform -1 0 1728 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5110
timestamp 1677622389
transform 1 0 1728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1677622389
transform 1 0 1736 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_296
timestamp 1677622389
transform 1 0 1744 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5114
timestamp 1677622389
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1677622389
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1677622389
transform 1 0 1856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1677622389
transform 1 0 1864 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_341
timestamp 1677622389
transform 1 0 1872 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5123
timestamp 1677622389
transform 1 0 1888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1677622389
transform 1 0 1896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1677622389
transform 1 0 1904 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_342
timestamp 1677622389
transform 1 0 1912 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5126
timestamp 1677622389
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1677622389
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1677622389
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_344
timestamp 1677622389
transform 1 0 1952 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5140
timestamp 1677622389
transform 1 0 1968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1677622389
transform 1 0 1976 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4162
timestamp 1677622389
transform 1 0 2044 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_297
timestamp 1677622389
transform 1 0 1984 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5142
timestamp 1677622389
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1677622389
transform 1 0 2088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1677622389
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1677622389
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1677622389
transform 1 0 2112 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_41
timestamp 1677622389
transform 1 0 2120 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5153
timestamp 1677622389
transform 1 0 2144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1677622389
transform 1 0 2152 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_298
timestamp 1677622389
transform -1 0 2256 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_346
timestamp 1677622389
transform 1 0 2256 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5166
timestamp 1677622389
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1677622389
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1677622389
transform 1 0 2288 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5177
timestamp 1677622389
transform 1 0 2384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1677622389
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1677622389
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1677622389
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1677622389
transform 1 0 2416 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4163
timestamp 1677622389
transform 1 0 2468 0 1 2475
box -3 -3 3 3
use OAI22X1  OAI22X1_199
timestamp 1677622389
transform 1 0 2424 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5189
timestamp 1677622389
transform 1 0 2464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1677622389
transform 1 0 2472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1677622389
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1677622389
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1677622389
transform 1 0 2496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1677622389
transform 1 0 2504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1677622389
transform 1 0 2512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1677622389
transform 1 0 2520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1677622389
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_210
timestamp 1677622389
transform 1 0 2536 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5210
timestamp 1677622389
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1677622389
transform 1 0 2584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1677622389
transform 1 0 2592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1677622389
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_347
timestamp 1677622389
transform 1 0 2608 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5220
timestamp 1677622389
transform 1 0 2624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1677622389
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4164
timestamp 1677622389
transform 1 0 2652 0 1 2475
box -3 -3 3 3
use FILL  FILL_5224
timestamp 1677622389
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1677622389
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_301
timestamp 1677622389
transform 1 0 2656 0 -1 2570
box -8 -3 104 105
use M3_M2  M3_M2_4165
timestamp 1677622389
transform 1 0 2764 0 1 2475
box -3 -3 3 3
use NOR2X1  NOR2X1_51
timestamp 1677622389
transform 1 0 2752 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5231
timestamp 1677622389
transform 1 0 2776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1677622389
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1677622389
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1677622389
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1677622389
transform 1 0 2808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1677622389
transform 1 0 2816 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_105
timestamp 1677622389
transform 1 0 2824 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5243
timestamp 1677622389
transform 1 0 2856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1677622389
transform 1 0 2864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1677622389
transform 1 0 2872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1677622389
transform 1 0 2880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1677622389
transform 1 0 2888 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_53
timestamp 1677622389
transform 1 0 2896 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5257
timestamp 1677622389
transform 1 0 2920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1677622389
transform 1 0 2928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1677622389
transform 1 0 2936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1677622389
transform 1 0 2944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1677622389
transform 1 0 2952 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_107
timestamp 1677622389
transform -1 0 2992 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5262
timestamp 1677622389
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1677622389
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1677622389
transform 1 0 3008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1677622389
transform 1 0 3016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1677622389
transform 1 0 3024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1677622389
transform 1 0 3032 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4166
timestamp 1677622389
transform 1 0 3052 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1677622389
transform 1 0 3084 0 1 2475
box -3 -3 3 3
use OAI22X1  OAI22X1_200
timestamp 1677622389
transform 1 0 3040 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5268
timestamp 1677622389
transform 1 0 3080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1677622389
transform 1 0 3088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1677622389
transform 1 0 3096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1677622389
transform 1 0 3104 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4168
timestamp 1677622389
transform 1 0 3124 0 1 2475
box -3 -3 3 3
use FILL  FILL_5274
timestamp 1677622389
transform 1 0 3112 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4169
timestamp 1677622389
transform 1 0 3164 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_304
timestamp 1677622389
transform 1 0 3120 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5275
timestamp 1677622389
transform 1 0 3216 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_350
timestamp 1677622389
transform 1 0 3224 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5276
timestamp 1677622389
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1677622389
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1677622389
transform 1 0 3256 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_43
timestamp 1677622389
transform 1 0 3264 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5281
timestamp 1677622389
transform 1 0 3288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1677622389
transform 1 0 3296 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_44
timestamp 1677622389
transform 1 0 3304 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5283
timestamp 1677622389
transform 1 0 3328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1677622389
transform 1 0 3336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1677622389
transform 1 0 3344 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_45
timestamp 1677622389
transform 1 0 3352 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5286
timestamp 1677622389
transform 1 0 3376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1677622389
transform 1 0 3384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1677622389
transform 1 0 3392 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_46
timestamp 1677622389
transform 1 0 3400 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_47
timestamp 1677622389
transform 1 0 3424 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5294
timestamp 1677622389
transform 1 0 3448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1677622389
transform 1 0 3456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1677622389
transform 1 0 3464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1677622389
transform 1 0 3472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1677622389
transform 1 0 3480 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_202
timestamp 1677622389
transform 1 0 3488 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5304
timestamp 1677622389
transform 1 0 3528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1677622389
transform 1 0 3536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1677622389
transform 1 0 3544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1677622389
transform 1 0 3552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1677622389
transform 1 0 3560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1677622389
transform 1 0 3568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1677622389
transform 1 0 3576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1677622389
transform 1 0 3584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1677622389
transform 1 0 3592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1677622389
transform 1 0 3600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1677622389
transform 1 0 3608 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_352
timestamp 1677622389
transform -1 0 3632 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5316
timestamp 1677622389
transform 1 0 3632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1677622389
transform 1 0 3640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1677622389
transform 1 0 3648 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_353
timestamp 1677622389
transform 1 0 3656 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5324
timestamp 1677622389
transform 1 0 3672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1677622389
transform 1 0 3680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1677622389
transform 1 0 3688 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_48
timestamp 1677622389
transform 1 0 3696 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_49
timestamp 1677622389
transform 1 0 3720 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5331
timestamp 1677622389
transform 1 0 3744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1677622389
transform 1 0 3752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1677622389
transform 1 0 3760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1677622389
transform 1 0 3768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1677622389
transform 1 0 3776 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1677622389
transform 1 0 3784 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5346
timestamp 1677622389
transform 1 0 3880 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_355
timestamp 1677622389
transform 1 0 3888 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5359
timestamp 1677622389
transform 1 0 3904 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_309
timestamp 1677622389
transform 1 0 3912 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5360
timestamp 1677622389
transform 1 0 4008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1677622389
transform 1 0 4016 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_310
timestamp 1677622389
transform -1 0 4120 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5362
timestamp 1677622389
transform 1 0 4120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1677622389
transform 1 0 4128 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_205
timestamp 1677622389
transform -1 0 4176 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5364
timestamp 1677622389
transform 1 0 4176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1677622389
transform 1 0 4184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1677622389
transform 1 0 4192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1677622389
transform 1 0 4200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1677622389
transform 1 0 4208 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_31
timestamp 1677622389
transform -1 0 4248 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5372
timestamp 1677622389
transform 1 0 4248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1677622389
transform 1 0 4256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5379
timestamp 1677622389
transform 1 0 4264 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_32
timestamp 1677622389
transform -1 0 4304 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5380
timestamp 1677622389
transform 1 0 4304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5381
timestamp 1677622389
transform 1 0 4312 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_356
timestamp 1677622389
transform 1 0 4320 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5382
timestamp 1677622389
transform 1 0 4336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5384
timestamp 1677622389
transform 1 0 4344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5386
timestamp 1677622389
transform 1 0 4352 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_207
timestamp 1677622389
transform 1 0 4360 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5388
timestamp 1677622389
transform 1 0 4400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5389
timestamp 1677622389
transform 1 0 4408 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_357
timestamp 1677622389
transform -1 0 4432 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5390
timestamp 1677622389
transform 1 0 4432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5391
timestamp 1677622389
transform 1 0 4440 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_33
timestamp 1677622389
transform 1 0 4448 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5392
timestamp 1677622389
transform 1 0 4480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5394
timestamp 1677622389
transform 1 0 4488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5396
timestamp 1677622389
transform 1 0 4496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5398
timestamp 1677622389
transform 1 0 4504 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_213
timestamp 1677622389
transform 1 0 4512 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5418
timestamp 1677622389
transform 1 0 4552 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_361
timestamp 1677622389
transform -1 0 4576 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_312
timestamp 1677622389
transform 1 0 4576 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5419
timestamp 1677622389
transform 1 0 4672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5420
timestamp 1677622389
transform 1 0 4680 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_313
timestamp 1677622389
transform 1 0 4688 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5421
timestamp 1677622389
transform 1 0 4784 0 -1 2570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_45
timestamp 1677622389
transform 1 0 4843 0 1 2470
box -10 -3 10 3
use M3_M2  M3_M2_4178
timestamp 1677622389
transform 1 0 156 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1677622389
transform 1 0 172 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1677622389
transform 1 0 164 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1677622389
transform 1 0 84 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4719
timestamp 1677622389
transform 1 0 116 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4246
timestamp 1677622389
transform 1 0 156 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4720
timestamp 1677622389
transform 1 0 164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1677622389
transform 1 0 180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1677622389
transform 1 0 84 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4335
timestamp 1677622389
transform 1 0 132 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4825
timestamp 1677622389
transform 1 0 188 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4336
timestamp 1677622389
transform 1 0 180 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4722
timestamp 1677622389
transform 1 0 260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1677622389
transform 1 0 228 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4289
timestamp 1677622389
transform 1 0 228 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4723
timestamp 1677622389
transform 1 0 324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1677622389
transform 1 0 372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1677622389
transform 1 0 340 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4290
timestamp 1677622389
transform 1 0 372 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4725
timestamp 1677622389
transform 1 0 436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1677622389
transform 1 0 452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1677622389
transform 1 0 468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1677622389
transform 1 0 476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1677622389
transform 1 0 436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1677622389
transform 1 0 460 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4291
timestamp 1677622389
transform 1 0 436 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4830
timestamp 1677622389
transform 1 0 484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1677622389
transform 1 0 500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1677622389
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1677622389
transform 1 0 508 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4337
timestamp 1677622389
transform 1 0 508 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4731
timestamp 1677622389
transform 1 0 532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1677622389
transform 1 0 532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1677622389
transform 1 0 588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1677622389
transform 1 0 564 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1677622389
transform 1 0 580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4292
timestamp 1677622389
transform 1 0 564 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1677622389
transform 1 0 604 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4835
timestamp 1677622389
transform 1 0 604 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1677622389
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4293
timestamp 1677622389
transform 1 0 612 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1677622389
transform 1 0 628 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4733
timestamp 1677622389
transform 1 0 628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1677622389
transform 1 0 644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1677622389
transform 1 0 644 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4294
timestamp 1677622389
transform 1 0 644 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4735
timestamp 1677622389
transform 1 0 660 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4170
timestamp 1677622389
transform 1 0 692 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1677622389
transform 1 0 716 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4736
timestamp 1677622389
transform 1 0 700 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1677622389
transform 1 0 716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1677622389
transform 1 0 692 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1677622389
transform 1 0 708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1677622389
transform 1 0 724 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4171
timestamp 1677622389
transform 1 0 732 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4738
timestamp 1677622389
transform 1 0 756 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4216
timestamp 1677622389
transform 1 0 772 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1677622389
transform 1 0 796 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4841
timestamp 1677622389
transform 1 0 796 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1677622389
transform 1 0 828 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4247
timestamp 1677622389
transform 1 0 828 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4739
timestamp 1677622389
transform 1 0 884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1677622389
transform 1 0 844 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4338
timestamp 1677622389
transform 1 0 860 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4740
timestamp 1677622389
transform 1 0 956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1677622389
transform 1 0 972 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4295
timestamp 1677622389
transform 1 0 964 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1677622389
transform 1 0 996 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4741
timestamp 1677622389
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1677622389
transform 1 0 1012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1677622389
transform 1 0 988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1677622389
transform 1 0 1012 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4296
timestamp 1677622389
transform 1 0 1012 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4906
timestamp 1677622389
transform 1 0 1036 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1677622389
transform 1 0 1084 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4261
timestamp 1677622389
transform 1 0 1076 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1677622389
transform 1 0 1076 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4744
timestamp 1677622389
transform 1 0 1108 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4262
timestamp 1677622389
transform 1 0 1108 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1677622389
transform 1 0 1116 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4845
timestamp 1677622389
transform 1 0 1132 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4298
timestamp 1677622389
transform 1 0 1132 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4846
timestamp 1677622389
transform 1 0 1156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1677622389
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4299
timestamp 1677622389
transform 1 0 1196 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4706
timestamp 1677622389
transform 1 0 1212 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4300
timestamp 1677622389
transform 1 0 1212 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4707
timestamp 1677622389
transform 1 0 1244 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1677622389
transform 1 0 1252 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1677622389
transform 1 0 1236 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4263
timestamp 1677622389
transform 1 0 1236 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4709
timestamp 1677622389
transform 1 0 1284 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4248
timestamp 1677622389
transform 1 0 1276 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4907
timestamp 1677622389
transform 1 0 1276 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4218
timestamp 1677622389
transform 1 0 1300 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4847
timestamp 1677622389
transform 1 0 1300 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4264
timestamp 1677622389
transform 1 0 1308 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1677622389
transform 1 0 1300 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1677622389
transform 1 0 1348 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4747
timestamp 1677622389
transform 1 0 1340 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4265
timestamp 1677622389
transform 1 0 1340 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1677622389
transform 1 0 1324 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1677622389
transform 1 0 1364 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1677622389
transform 1 0 1372 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4848
timestamp 1677622389
transform 1 0 1372 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4172
timestamp 1677622389
transform 1 0 1436 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1677622389
transform 1 0 1412 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1677622389
transform 1 0 1444 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4748
timestamp 1677622389
transform 1 0 1444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1677622389
transform 1 0 1396 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4266
timestamp 1677622389
transform 1 0 1420 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1677622389
transform 1 0 1460 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1677622389
transform 1 0 1492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1677622389
transform 1 0 1508 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1677622389
transform 1 0 1508 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1677622389
transform 1 0 1524 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4749
timestamp 1677622389
transform 1 0 1516 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4268
timestamp 1677622389
transform 1 0 1508 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1677622389
transform 1 0 1548 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1677622389
transform 1 0 1572 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4850
timestamp 1677622389
transform 1 0 1580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4223
timestamp 1677622389
transform 1 0 1596 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4750
timestamp 1677622389
transform 1 0 1596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1677622389
transform 1 0 1612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1677622389
transform 1 0 1604 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4303
timestamp 1677622389
transform 1 0 1612 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1677622389
transform 1 0 1668 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1677622389
transform 1 0 1716 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4752
timestamp 1677622389
transform 1 0 1676 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1677622389
transform 1 0 1724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1677622389
transform 1 0 1668 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4269
timestamp 1677622389
transform 1 0 1676 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4853
timestamp 1677622389
transform 1 0 1756 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4304
timestamp 1677622389
transform 1 0 1716 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1677622389
transform 1 0 1804 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1677622389
transform 1 0 1804 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4754
timestamp 1677622389
transform 1 0 1812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1677622389
transform 1 0 1828 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4305
timestamp 1677622389
transform 1 0 1804 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4854
timestamp 1677622389
transform 1 0 1820 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4306
timestamp 1677622389
transform 1 0 1836 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4855
timestamp 1677622389
transform 1 0 1852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1677622389
transform 1 0 1852 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1677622389
transform 1 0 1860 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1677622389
transform 1 0 1884 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4195
timestamp 1677622389
transform 1 0 1908 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4711
timestamp 1677622389
transform 1 0 1908 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1677622389
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4270
timestamp 1677622389
transform 1 0 1900 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1677622389
transform 1 0 1948 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4757
timestamp 1677622389
transform 1 0 1940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1677622389
transform 1 0 1956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1677622389
transform 1 0 1948 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1677622389
transform 1 0 1964 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4307
timestamp 1677622389
transform 1 0 1932 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1677622389
transform 1 0 1972 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1677622389
transform 1 0 1964 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4911
timestamp 1677622389
transform 1 0 1996 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1677622389
transform 1 0 2028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1677622389
transform 1 0 2020 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4180
timestamp 1677622389
transform 1 0 2052 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4760
timestamp 1677622389
transform 1 0 2044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1677622389
transform 1 0 2060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1677622389
transform 1 0 2052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1677622389
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1677622389
transform 1 0 2092 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4272
timestamp 1677622389
transform 1 0 2092 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1677622389
transform 1 0 2116 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4860
timestamp 1677622389
transform 1 0 2116 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4181
timestamp 1677622389
transform 1 0 2164 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1677622389
transform 1 0 2156 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4763
timestamp 1677622389
transform 1 0 2156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1677622389
transform 1 0 2172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1677622389
transform 1 0 2188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1677622389
transform 1 0 2156 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4273
timestamp 1677622389
transform 1 0 2172 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4862
timestamp 1677622389
transform 1 0 2188 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4198
timestamp 1677622389
transform 1 0 2220 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1677622389
transform 1 0 2212 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4766
timestamp 1677622389
transform 1 0 2276 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4182
timestamp 1677622389
transform 1 0 2300 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1677622389
transform 1 0 2340 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4767
timestamp 1677622389
transform 1 0 2316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1677622389
transform 1 0 2332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1677622389
transform 1 0 2308 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4275
timestamp 1677622389
transform 1 0 2316 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1677622389
transform 1 0 2332 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1677622389
transform 1 0 2348 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1677622389
transform 1 0 2364 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4913
timestamp 1677622389
transform 1 0 2356 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4199
timestamp 1677622389
transform 1 0 2388 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4769
timestamp 1677622389
transform 1 0 2380 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4225
timestamp 1677622389
transform 1 0 2396 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1677622389
transform 1 0 2396 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1677622389
transform 1 0 2420 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1677622389
transform 1 0 2436 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4864
timestamp 1677622389
transform 1 0 2452 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4185
timestamp 1677622389
transform 1 0 2476 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1677622389
transform 1 0 2468 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4914
timestamp 1677622389
transform 1 0 2476 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1677622389
transform 1 0 2556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1677622389
transform 1 0 2572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1677622389
transform 1 0 2580 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4277
timestamp 1677622389
transform 1 0 2572 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4865
timestamp 1677622389
transform 1 0 2588 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4313
timestamp 1677622389
transform 1 0 2580 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1677622389
transform 1 0 2644 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4773
timestamp 1677622389
transform 1 0 2644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1677622389
transform 1 0 2660 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4278
timestamp 1677622389
transform 1 0 2636 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1677622389
transform 1 0 2660 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4866
timestamp 1677622389
transform 1 0 2708 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4227
timestamp 1677622389
transform 1 0 2716 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4867
timestamp 1677622389
transform 1 0 2716 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4228
timestamp 1677622389
transform 1 0 2748 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4775
timestamp 1677622389
transform 1 0 2748 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4229
timestamp 1677622389
transform 1 0 2788 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4776
timestamp 1677622389
transform 1 0 2788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1677622389
transform 1 0 2844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1677622389
transform 1 0 2764 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4314
timestamp 1677622389
transform 1 0 2764 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1677622389
transform 1 0 2812 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4910
timestamp 1677622389
transform 1 0 2860 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1677622389
transform 1 0 2892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1677622389
transform 1 0 2884 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4316
timestamp 1677622389
transform 1 0 2884 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1677622389
transform 1 0 2996 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4779
timestamp 1677622389
transform 1 0 2940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1677622389
transform 1 0 2996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1677622389
transform 1 0 3020 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4317
timestamp 1677622389
transform 1 0 2940 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4781
timestamp 1677622389
transform 1 0 3044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1677622389
transform 1 0 3036 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4318
timestamp 1677622389
transform 1 0 3036 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1677622389
transform 1 0 3076 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4782
timestamp 1677622389
transform 1 0 3052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1677622389
transform 1 0 3068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1677622389
transform 1 0 3084 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4253
timestamp 1677622389
transform 1 0 3092 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4872
timestamp 1677622389
transform 1 0 3060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1677622389
transform 1 0 3076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1677622389
transform 1 0 3092 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4319
timestamp 1677622389
transform 1 0 3060 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4875
timestamp 1677622389
transform 1 0 3108 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4320
timestamp 1677622389
transform 1 0 3108 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1677622389
transform 1 0 3164 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1677622389
transform 1 0 3180 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4876
timestamp 1677622389
transform 1 0 3172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1677622389
transform 1 0 3188 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4321
timestamp 1677622389
transform 1 0 3180 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4877
timestamp 1677622389
transform 1 0 3236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1677622389
transform 1 0 3244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4322
timestamp 1677622389
transform 1 0 3244 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1677622389
transform 1 0 3260 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4712
timestamp 1677622389
transform 1 0 3292 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1677622389
transform 1 0 3284 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4186
timestamp 1677622389
transform 1 0 3324 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1677622389
transform 1 0 3308 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4699
timestamp 1677622389
transform 1 0 3316 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1677622389
transform 1 0 3348 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1677622389
transform 1 0 3380 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1677622389
transform 1 0 3364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1677622389
transform 1 0 3372 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4254
timestamp 1677622389
transform 1 0 3372 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4715
timestamp 1677622389
transform 1 0 3396 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4255
timestamp 1677622389
transform 1 0 3396 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4702
timestamp 1677622389
transform 1 0 3444 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4234
timestamp 1677622389
transform 1 0 3452 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4787
timestamp 1677622389
transform 1 0 3452 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4280
timestamp 1677622389
transform 1 0 3444 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4788
timestamp 1677622389
transform 1 0 3476 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4208
timestamp 1677622389
transform 1 0 3500 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4716
timestamp 1677622389
transform 1 0 3500 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4200
timestamp 1677622389
transform 1 0 3516 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1677622389
transform 1 0 3540 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1677622389
transform 1 0 3524 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4789
timestamp 1677622389
transform 1 0 3524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1677622389
transform 1 0 3540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1677622389
transform 1 0 3508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1677622389
transform 1 0 3532 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4187
timestamp 1677622389
transform 1 0 3556 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4881
timestamp 1677622389
transform 1 0 3556 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4202
timestamp 1677622389
transform 1 0 3572 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4791
timestamp 1677622389
transform 1 0 3580 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4324
timestamp 1677622389
transform 1 0 3580 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1677622389
transform 1 0 3604 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4792
timestamp 1677622389
transform 1 0 3596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1677622389
transform 1 0 3612 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4281
timestamp 1677622389
transform 1 0 3596 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4882
timestamp 1677622389
transform 1 0 3604 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1677622389
transform 1 0 3628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1677622389
transform 1 0 3644 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4282
timestamp 1677622389
transform 1 0 3660 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1677622389
transform 1 0 3732 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1677622389
transform 1 0 3716 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4795
timestamp 1677622389
transform 1 0 3732 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4257
timestamp 1677622389
transform 1 0 3780 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4884
timestamp 1677622389
transform 1 0 3780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1677622389
transform 1 0 3796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1677622389
transform 1 0 3820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1677622389
transform 1 0 3844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1677622389
transform 1 0 3836 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4209
timestamp 1677622389
transform 1 0 3876 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4799
timestamp 1677622389
transform 1 0 3876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1677622389
transform 1 0 3892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1677622389
transform 1 0 3900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1677622389
transform 1 0 3860 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4325
timestamp 1677622389
transform 1 0 3860 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1677622389
transform 1 0 3892 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1677622389
transform 1 0 3932 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1677622389
transform 1 0 3924 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1677622389
transform 1 0 3956 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4802
timestamp 1677622389
transform 1 0 3956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1677622389
transform 1 0 3924 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1677622389
transform 1 0 3932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1677622389
transform 1 0 3948 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4284
timestamp 1677622389
transform 1 0 3956 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1677622389
transform 1 0 3940 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1677622389
transform 1 0 3980 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4803
timestamp 1677622389
transform 1 0 3972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1677622389
transform 1 0 3980 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4239
timestamp 1677622389
transform 1 0 4004 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4804
timestamp 1677622389
transform 1 0 3996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1677622389
transform 1 0 4004 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4176
timestamp 1677622389
transform 1 0 4108 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1677622389
transform 1 0 4100 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4806
timestamp 1677622389
transform 1 0 4020 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1677622389
transform 1 0 4052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1677622389
transform 1 0 4012 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1677622389
transform 1 0 4100 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4327
timestamp 1677622389
transform 1 0 4052 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1677622389
transform 1 0 4116 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1677622389
transform 1 0 4140 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1677622389
transform 1 0 4172 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1677622389
transform 1 0 4148 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4808
timestamp 1677622389
transform 1 0 4148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1677622389
transform 1 0 4164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1677622389
transform 1 0 4180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1677622389
transform 1 0 4140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1677622389
transform 1 0 4156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1677622389
transform 1 0 4172 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4241
timestamp 1677622389
transform 1 0 4220 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4811
timestamp 1677622389
transform 1 0 4220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1677622389
transform 1 0 4196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1677622389
transform 1 0 4212 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4285
timestamp 1677622389
transform 1 0 4220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1677622389
transform 1 0 4244 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4812
timestamp 1677622389
transform 1 0 4268 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4258
timestamp 1677622389
transform 1 0 4276 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4898
timestamp 1677622389
transform 1 0 4228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1677622389
transform 1 0 4244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4286
timestamp 1677622389
transform 1 0 4268 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1677622389
transform 1 0 4228 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1677622389
transform 1 0 4260 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1677622389
transform 1 0 4340 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4813
timestamp 1677622389
transform 1 0 4340 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4259
timestamp 1677622389
transform 1 0 4364 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4814
timestamp 1677622389
transform 1 0 4372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1677622389
transform 1 0 4396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1677622389
transform 1 0 4412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1677622389
transform 1 0 4420 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4205
timestamp 1677622389
transform 1 0 4460 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4703
timestamp 1677622389
transform 1 0 4460 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1677622389
transform 1 0 4452 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1677622389
transform 1 0 4468 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4340
timestamp 1677622389
transform 1 0 4460 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4718
timestamp 1677622389
transform 1 0 4508 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4243
timestamp 1677622389
transform 1 0 4532 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4818
timestamp 1677622389
transform 1 0 4516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1677622389
transform 1 0 4508 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4331
timestamp 1677622389
transform 1 0 4508 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1677622389
transform 1 0 4524 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4819
timestamp 1677622389
transform 1 0 4540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1677622389
transform 1 0 4532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1677622389
transform 1 0 4572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1677622389
transform 1 0 4580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4244
timestamp 1677622389
transform 1 0 4620 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4821
timestamp 1677622389
transform 1 0 4620 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4287
timestamp 1677622389
transform 1 0 4644 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4904
timestamp 1677622389
transform 1 0 4668 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4332
timestamp 1677622389
transform 1 0 4604 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1677622389
transform 1 0 4668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1677622389
transform 1 0 4604 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1677622389
transform 1 0 4636 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4822
timestamp 1677622389
transform 1 0 4724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1677622389
transform 1 0 4780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1677622389
transform 1 0 4700 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4288
timestamp 1677622389
transform 1 0 4724 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1677622389
transform 1 0 4740 0 1 2395
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_46
timestamp 1677622389
transform 1 0 48 0 1 2370
box -10 -3 10 3
use M3_M2  M3_M2_4343
timestamp 1677622389
transform 1 0 164 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1677622389
transform 1 0 180 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_314
timestamp 1677622389
transform 1 0 72 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_362
timestamp 1677622389
transform -1 0 184 0 1 2370
box -9 -3 26 105
use FILL  FILL_5422
timestamp 1677622389
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5423
timestamp 1677622389
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5424
timestamp 1677622389
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5425
timestamp 1677622389
transform 1 0 208 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_315
timestamp 1677622389
transform 1 0 216 0 1 2370
box -8 -3 104 105
use FILL  FILL_5426
timestamp 1677622389
transform 1 0 312 0 1 2370
box -8 -3 16 105
use FILL  FILL_5427
timestamp 1677622389
transform 1 0 320 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_316
timestamp 1677622389
transform 1 0 328 0 1 2370
box -8 -3 104 105
use FILL  FILL_5428
timestamp 1677622389
transform 1 0 424 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_214
timestamp 1677622389
transform -1 0 472 0 1 2370
box -8 -3 46 105
use FILL  FILL_5429
timestamp 1677622389
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_5430
timestamp 1677622389
transform 1 0 480 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4345
timestamp 1677622389
transform 1 0 532 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_210
timestamp 1677622389
transform 1 0 488 0 1 2370
box -8 -3 46 105
use FILL  FILL_5431
timestamp 1677622389
transform 1 0 528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5435
timestamp 1677622389
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5436
timestamp 1677622389
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5437
timestamp 1677622389
transform 1 0 552 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_211
timestamp 1677622389
transform 1 0 560 0 1 2370
box -8 -3 46 105
use FILL  FILL_5439
timestamp 1677622389
transform 1 0 600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5440
timestamp 1677622389
transform 1 0 608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5441
timestamp 1677622389
transform 1 0 616 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_366
timestamp 1677622389
transform 1 0 624 0 1 2370
box -9 -3 26 105
use FILL  FILL_5442
timestamp 1677622389
transform 1 0 640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5443
timestamp 1677622389
transform 1 0 648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5444
timestamp 1677622389
transform 1 0 656 0 1 2370
box -8 -3 16 105
use FILL  FILL_5445
timestamp 1677622389
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5446
timestamp 1677622389
transform 1 0 672 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_218
timestamp 1677622389
transform 1 0 680 0 1 2370
box -8 -3 46 105
use FILL  FILL_5447
timestamp 1677622389
transform 1 0 720 0 1 2370
box -8 -3 16 105
use FILL  FILL_5448
timestamp 1677622389
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_5449
timestamp 1677622389
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_5456
timestamp 1677622389
transform 1 0 744 0 1 2370
box -8 -3 16 105
use FILL  FILL_5458
timestamp 1677622389
transform 1 0 752 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_108
timestamp 1677622389
transform 1 0 760 0 1 2370
box -8 -3 34 105
use FILL  FILL_5460
timestamp 1677622389
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5466
timestamp 1677622389
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_5468
timestamp 1677622389
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_5470
timestamp 1677622389
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_5472
timestamp 1677622389
transform 1 0 824 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_321
timestamp 1677622389
transform 1 0 832 0 1 2370
box -8 -3 104 105
use FILL  FILL_5473
timestamp 1677622389
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_5481
timestamp 1677622389
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5483
timestamp 1677622389
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5485
timestamp 1677622389
transform 1 0 952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5487
timestamp 1677622389
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5489
timestamp 1677622389
transform 1 0 968 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_220
timestamp 1677622389
transform 1 0 976 0 1 2370
box -8 -3 46 105
use FILL  FILL_5491
timestamp 1677622389
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5492
timestamp 1677622389
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5495
timestamp 1677622389
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_5497
timestamp 1677622389
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use FILL  FILL_5499
timestamp 1677622389
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_5501
timestamp 1677622389
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_5503
timestamp 1677622389
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_5505
timestamp 1677622389
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_5507
timestamp 1677622389
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_222
timestamp 1677622389
transform 1 0 1088 0 1 2370
box -8 -3 46 105
use FILL  FILL_5509
timestamp 1677622389
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_5510
timestamp 1677622389
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use FILL  FILL_5511
timestamp 1677622389
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5512
timestamp 1677622389
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5517
timestamp 1677622389
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_5519
timestamp 1677622389
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_5521
timestamp 1677622389
transform 1 0 1176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5523
timestamp 1677622389
transform 1 0 1184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5525
timestamp 1677622389
transform 1 0 1192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5527
timestamp 1677622389
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_110
timestamp 1677622389
transform -1 0 1240 0 1 2370
box -8 -3 34 105
use FILL  FILL_5528
timestamp 1677622389
transform 1 0 1240 0 1 2370
box -8 -3 16 105
use FILL  FILL_5532
timestamp 1677622389
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_5534
timestamp 1677622389
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_5536
timestamp 1677622389
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5538
timestamp 1677622389
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_5540
timestamp 1677622389
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5542
timestamp 1677622389
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_5544
timestamp 1677622389
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_5546
timestamp 1677622389
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_111
timestamp 1677622389
transform -1 0 1344 0 1 2370
box -8 -3 34 105
use FILL  FILL_5547
timestamp 1677622389
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4346
timestamp 1677622389
transform 1 0 1364 0 1 2375
box -3 -3 3 3
use FILL  FILL_5552
timestamp 1677622389
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5554
timestamp 1677622389
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_5556
timestamp 1677622389
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4347
timestamp 1677622389
transform 1 0 1396 0 1 2375
box -3 -3 3 3
use FILL  FILL_5558
timestamp 1677622389
transform 1 0 1376 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_322
timestamp 1677622389
transform 1 0 1384 0 1 2370
box -8 -3 104 105
use FILL  FILL_5560
timestamp 1677622389
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5574
timestamp 1677622389
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5576
timestamp 1677622389
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_368
timestamp 1677622389
transform 1 0 1504 0 1 2370
box -9 -3 26 105
use FILL  FILL_5578
timestamp 1677622389
transform 1 0 1520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5582
timestamp 1677622389
transform 1 0 1528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5584
timestamp 1677622389
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5585
timestamp 1677622389
transform 1 0 1544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5586
timestamp 1677622389
transform 1 0 1552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5587
timestamp 1677622389
transform 1 0 1560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5590
timestamp 1677622389
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5591
timestamp 1677622389
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_212
timestamp 1677622389
transform -1 0 1624 0 1 2370
box -8 -3 46 105
use FILL  FILL_5592
timestamp 1677622389
transform 1 0 1624 0 1 2370
box -8 -3 16 105
use FILL  FILL_5593
timestamp 1677622389
transform 1 0 1632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5594
timestamp 1677622389
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5595
timestamp 1677622389
transform 1 0 1648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5596
timestamp 1677622389
transform 1 0 1656 0 1 2370
box -8 -3 16 105
use FILL  FILL_5597
timestamp 1677622389
transform 1 0 1664 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_323
timestamp 1677622389
transform -1 0 1768 0 1 2370
box -8 -3 104 105
use FILL  FILL_5598
timestamp 1677622389
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use FILL  FILL_5611
timestamp 1677622389
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5613
timestamp 1677622389
transform 1 0 1784 0 1 2370
box -8 -3 16 105
use FILL  FILL_5614
timestamp 1677622389
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5615
timestamp 1677622389
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4348
timestamp 1677622389
transform 1 0 1820 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_224
timestamp 1677622389
transform 1 0 1808 0 1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4349
timestamp 1677622389
transform 1 0 1860 0 1 2375
box -3 -3 3 3
use FILL  FILL_5616
timestamp 1677622389
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_5617
timestamp 1677622389
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5618
timestamp 1677622389
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_5619
timestamp 1677622389
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use FILL  FILL_5620
timestamp 1677622389
transform 1 0 1880 0 1 2370
box -8 -3 16 105
use FILL  FILL_5621
timestamp 1677622389
transform 1 0 1888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5629
timestamp 1677622389
transform 1 0 1896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5631
timestamp 1677622389
transform 1 0 1904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5633
timestamp 1677622389
transform 1 0 1912 0 1 2370
box -8 -3 16 105
use FILL  FILL_5635
timestamp 1677622389
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_213
timestamp 1677622389
transform -1 0 1968 0 1 2370
box -8 -3 46 105
use FILL  FILL_5636
timestamp 1677622389
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use FILL  FILL_5637
timestamp 1677622389
transform 1 0 1976 0 1 2370
box -8 -3 16 105
use FILL  FILL_5638
timestamp 1677622389
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_5639
timestamp 1677622389
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use FILL  FILL_5640
timestamp 1677622389
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_5641
timestamp 1677622389
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5642
timestamp 1677622389
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5643
timestamp 1677622389
transform 1 0 2024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5644
timestamp 1677622389
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_226
timestamp 1677622389
transform 1 0 2040 0 1 2370
box -8 -3 46 105
use FILL  FILL_5648
timestamp 1677622389
transform 1 0 2080 0 1 2370
box -8 -3 16 105
use FILL  FILL_5649
timestamp 1677622389
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_5650
timestamp 1677622389
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5651
timestamp 1677622389
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5658
timestamp 1677622389
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5660
timestamp 1677622389
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5661
timestamp 1677622389
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use FILL  FILL_5662
timestamp 1677622389
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4350
timestamp 1677622389
transform 1 0 2156 0 1 2375
box -3 -3 3 3
use FILL  FILL_5663
timestamp 1677622389
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_227
timestamp 1677622389
transform 1 0 2152 0 1 2370
box -8 -3 46 105
use FILL  FILL_5664
timestamp 1677622389
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5668
timestamp 1677622389
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5670
timestamp 1677622389
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5672
timestamp 1677622389
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use FILL  FILL_5674
timestamp 1677622389
transform 1 0 2224 0 1 2370
box -8 -3 16 105
use FILL  FILL_5676
timestamp 1677622389
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_5678
timestamp 1677622389
transform 1 0 2240 0 1 2370
box -8 -3 16 105
use FILL  FILL_5679
timestamp 1677622389
transform 1 0 2248 0 1 2370
box -8 -3 16 105
use FILL  FILL_5680
timestamp 1677622389
transform 1 0 2256 0 1 2370
box -8 -3 16 105
use FILL  FILL_5682
timestamp 1677622389
transform 1 0 2264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5684
timestamp 1677622389
transform 1 0 2272 0 1 2370
box -8 -3 16 105
use FILL  FILL_5686
timestamp 1677622389
transform 1 0 2280 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4351
timestamp 1677622389
transform 1 0 2300 0 1 2375
box -3 -3 3 3
use FILL  FILL_5688
timestamp 1677622389
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_229
timestamp 1677622389
transform 1 0 2296 0 1 2370
box -8 -3 46 105
use FILL  FILL_5689
timestamp 1677622389
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5693
timestamp 1677622389
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5695
timestamp 1677622389
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5697
timestamp 1677622389
transform 1 0 2360 0 1 2370
box -8 -3 16 105
use FILL  FILL_5699
timestamp 1677622389
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use FILL  FILL_5701
timestamp 1677622389
transform 1 0 2376 0 1 2370
box -8 -3 16 105
use FILL  FILL_5703
timestamp 1677622389
transform 1 0 2384 0 1 2370
box -8 -3 16 105
use FILL  FILL_5704
timestamp 1677622389
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_5705
timestamp 1677622389
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use FILL  FILL_5706
timestamp 1677622389
transform 1 0 2408 0 1 2370
box -8 -3 16 105
use FILL  FILL_5707
timestamp 1677622389
transform 1 0 2416 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4352
timestamp 1677622389
transform 1 0 2436 0 1 2375
box -3 -3 3 3
use FILL  FILL_5708
timestamp 1677622389
transform 1 0 2424 0 1 2370
box -8 -3 16 105
use FILL  FILL_5709
timestamp 1677622389
transform 1 0 2432 0 1 2370
box -8 -3 16 105
use FILL  FILL_5712
timestamp 1677622389
transform 1 0 2440 0 1 2370
box -8 -3 16 105
use FILL  FILL_5714
timestamp 1677622389
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_5716
timestamp 1677622389
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_5718
timestamp 1677622389
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_5719
timestamp 1677622389
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use FILL  FILL_5720
timestamp 1677622389
transform 1 0 2480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5722
timestamp 1677622389
transform 1 0 2488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5724
timestamp 1677622389
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_375
timestamp 1677622389
transform 1 0 2504 0 1 2370
box -9 -3 26 105
use FILL  FILL_5726
timestamp 1677622389
transform 1 0 2520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5730
timestamp 1677622389
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5731
timestamp 1677622389
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5732
timestamp 1677622389
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5733
timestamp 1677622389
transform 1 0 2552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5734
timestamp 1677622389
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_376
timestamp 1677622389
transform -1 0 2584 0 1 2370
box -9 -3 26 105
use FILL  FILL_5735
timestamp 1677622389
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_5736
timestamp 1677622389
transform 1 0 2592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5737
timestamp 1677622389
transform 1 0 2600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5738
timestamp 1677622389
transform 1 0 2608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5739
timestamp 1677622389
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_231
timestamp 1677622389
transform 1 0 2624 0 1 2370
box -8 -3 46 105
use FILL  FILL_5740
timestamp 1677622389
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5741
timestamp 1677622389
transform 1 0 2672 0 1 2370
box -8 -3 16 105
use FILL  FILL_5742
timestamp 1677622389
transform 1 0 2680 0 1 2370
box -8 -3 16 105
use FILL  FILL_5743
timestamp 1677622389
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use FILL  FILL_5744
timestamp 1677622389
transform 1 0 2696 0 1 2370
box -8 -3 16 105
use FILL  FILL_5745
timestamp 1677622389
transform 1 0 2704 0 1 2370
box -8 -3 16 105
use FILL  FILL_5746
timestamp 1677622389
transform 1 0 2712 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_377
timestamp 1677622389
transform 1 0 2720 0 1 2370
box -9 -3 26 105
use FILL  FILL_5747
timestamp 1677622389
transform 1 0 2736 0 1 2370
box -8 -3 16 105
use FILL  FILL_5748
timestamp 1677622389
transform 1 0 2744 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_328
timestamp 1677622389
transform 1 0 2752 0 1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4353
timestamp 1677622389
transform 1 0 2860 0 1 2375
box -3 -3 3 3
use FILL  FILL_5753
timestamp 1677622389
transform 1 0 2848 0 1 2370
box -8 -3 16 105
use FILL  FILL_5763
timestamp 1677622389
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5765
timestamp 1677622389
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1677622389
transform 1 0 2872 0 1 2370
box -8 -3 32 105
use FILL  FILL_5766
timestamp 1677622389
transform 1 0 2896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5768
timestamp 1677622389
transform 1 0 2904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5770
timestamp 1677622389
transform 1 0 2912 0 1 2370
box -8 -3 16 105
use FILL  FILL_5772
timestamp 1677622389
transform 1 0 2920 0 1 2370
box -8 -3 16 105
use FILL  FILL_5774
timestamp 1677622389
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_329
timestamp 1677622389
transform -1 0 3032 0 1 2370
box -8 -3 104 105
use FILL  FILL_5775
timestamp 1677622389
transform 1 0 3032 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_378
timestamp 1677622389
transform 1 0 3040 0 1 2370
box -9 -3 26 105
use OAI22X1  OAI22X1_214
timestamp 1677622389
transform -1 0 3096 0 1 2370
box -8 -3 46 105
use FILL  FILL_5776
timestamp 1677622389
transform 1 0 3096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5790
timestamp 1677622389
transform 1 0 3104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5792
timestamp 1677622389
transform 1 0 3112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5793
timestamp 1677622389
transform 1 0 3120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5794
timestamp 1677622389
transform 1 0 3128 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_379
timestamp 1677622389
transform 1 0 3136 0 1 2370
box -9 -3 26 105
use FILL  FILL_5795
timestamp 1677622389
transform 1 0 3152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5796
timestamp 1677622389
transform 1 0 3160 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_55
timestamp 1677622389
transform -1 0 3192 0 1 2370
box -5 -3 28 105
use FILL  FILL_5797
timestamp 1677622389
transform 1 0 3192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5798
timestamp 1677622389
transform 1 0 3200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5799
timestamp 1677622389
transform 1 0 3208 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_56
timestamp 1677622389
transform 1 0 3216 0 1 2370
box -5 -3 28 105
use FILL  FILL_5800
timestamp 1677622389
transform 1 0 3240 0 1 2370
box -8 -3 16 105
use FILL  FILL_5801
timestamp 1677622389
transform 1 0 3248 0 1 2370
box -8 -3 16 105
use FILL  FILL_5802
timestamp 1677622389
transform 1 0 3256 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_57
timestamp 1677622389
transform -1 0 3288 0 1 2370
box -5 -3 28 105
use FILL  FILL_5803
timestamp 1677622389
transform 1 0 3288 0 1 2370
box -8 -3 16 105
use FILL  FILL_5804
timestamp 1677622389
transform 1 0 3296 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_34
timestamp 1677622389
transform -1 0 3336 0 1 2370
box -8 -3 40 105
use FILL  FILL_5805
timestamp 1677622389
transform 1 0 3336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5813
timestamp 1677622389
transform 1 0 3344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5814
timestamp 1677622389
transform 1 0 3352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5815
timestamp 1677622389
transform 1 0 3360 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_35
timestamp 1677622389
transform -1 0 3400 0 1 2370
box -8 -3 40 105
use FILL  FILL_5816
timestamp 1677622389
transform 1 0 3400 0 1 2370
box -8 -3 16 105
use FILL  FILL_5817
timestamp 1677622389
transform 1 0 3408 0 1 2370
box -8 -3 16 105
use FILL  FILL_5818
timestamp 1677622389
transform 1 0 3416 0 1 2370
box -8 -3 16 105
use FILL  FILL_5819
timestamp 1677622389
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_36
timestamp 1677622389
transform -1 0 3464 0 1 2370
box -8 -3 40 105
use FILL  FILL_5820
timestamp 1677622389
transform 1 0 3464 0 1 2370
box -8 -3 16 105
use FILL  FILL_5830
timestamp 1677622389
transform 1 0 3472 0 1 2370
box -8 -3 16 105
use FILL  FILL_5832
timestamp 1677622389
transform 1 0 3480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5834
timestamp 1677622389
transform 1 0 3488 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4354
timestamp 1677622389
transform 1 0 3508 0 1 2375
box -3 -3 3 3
use FILL  FILL_5835
timestamp 1677622389
transform 1 0 3496 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_232
timestamp 1677622389
transform 1 0 3504 0 1 2370
box -8 -3 46 105
use FILL  FILL_5836
timestamp 1677622389
transform 1 0 3544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5840
timestamp 1677622389
transform 1 0 3552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5842
timestamp 1677622389
transform 1 0 3560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5844
timestamp 1677622389
transform 1 0 3568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5845
timestamp 1677622389
transform 1 0 3576 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4355
timestamp 1677622389
transform 1 0 3612 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1677622389
transform 1 0 3628 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_218
timestamp 1677622389
transform 1 0 3584 0 1 2370
box -8 -3 46 105
use FILL  FILL_5846
timestamp 1677622389
transform 1 0 3624 0 1 2370
box -8 -3 16 105
use FILL  FILL_5847
timestamp 1677622389
transform 1 0 3632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5848
timestamp 1677622389
transform 1 0 3640 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_381
timestamp 1677622389
transform -1 0 3664 0 1 2370
box -9 -3 26 105
use FILL  FILL_5849
timestamp 1677622389
transform 1 0 3664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5851
timestamp 1677622389
transform 1 0 3672 0 1 2370
box -8 -3 16 105
use FILL  FILL_5852
timestamp 1677622389
transform 1 0 3680 0 1 2370
box -8 -3 16 105
use FILL  FILL_5853
timestamp 1677622389
transform 1 0 3688 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_332
timestamp 1677622389
transform -1 0 3792 0 1 2370
box -8 -3 104 105
use FILL  FILL_5854
timestamp 1677622389
transform 1 0 3792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5855
timestamp 1677622389
transform 1 0 3800 0 1 2370
box -8 -3 16 105
use FILL  FILL_5859
timestamp 1677622389
transform 1 0 3808 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_60
timestamp 1677622389
transform 1 0 3816 0 1 2370
box -5 -3 28 105
use FILL  FILL_5861
timestamp 1677622389
transform 1 0 3840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5862
timestamp 1677622389
transform 1 0 3848 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_233
timestamp 1677622389
transform 1 0 3856 0 1 2370
box -8 -3 46 105
use FILL  FILL_5863
timestamp 1677622389
transform 1 0 3896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5870
timestamp 1677622389
transform 1 0 3904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5872
timestamp 1677622389
transform 1 0 3912 0 1 2370
box -8 -3 16 105
use FILL  FILL_5874
timestamp 1677622389
transform 1 0 3920 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_219
timestamp 1677622389
transform 1 0 3928 0 1 2370
box -8 -3 46 105
use FILL  FILL_5875
timestamp 1677622389
transform 1 0 3968 0 1 2370
box -8 -3 16 105
use FILL  FILL_5878
timestamp 1677622389
transform 1 0 3976 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_383
timestamp 1677622389
transform -1 0 4000 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_384
timestamp 1677622389
transform -1 0 4016 0 1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_334
timestamp 1677622389
transform -1 0 4112 0 1 2370
box -8 -3 104 105
use FILL  FILL_5879
timestamp 1677622389
transform 1 0 4112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5896
timestamp 1677622389
transform 1 0 4120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5897
timestamp 1677622389
transform 1 0 4128 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4357
timestamp 1677622389
transform 1 0 4148 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_221
timestamp 1677622389
transform 1 0 4136 0 1 2370
box -8 -3 46 105
use FILL  FILL_5898
timestamp 1677622389
transform 1 0 4176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5899
timestamp 1677622389
transform 1 0 4184 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_222
timestamp 1677622389
transform 1 0 4192 0 1 2370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_335
timestamp 1677622389
transform 1 0 4232 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_386
timestamp 1677622389
transform 1 0 4328 0 1 2370
box -9 -3 26 105
use FILL  FILL_5900
timestamp 1677622389
transform 1 0 4344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5911
timestamp 1677622389
transform 1 0 4352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5913
timestamp 1677622389
transform 1 0 4360 0 1 2370
box -8 -3 16 105
use FILL  FILL_5914
timestamp 1677622389
transform 1 0 4368 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_235
timestamp 1677622389
transform -1 0 4416 0 1 2370
box -8 -3 46 105
use FILL  FILL_5915
timestamp 1677622389
transform 1 0 4416 0 1 2370
box -8 -3 16 105
use FILL  FILL_5919
timestamp 1677622389
transform 1 0 4424 0 1 2370
box -8 -3 16 105
use FILL  FILL_5921
timestamp 1677622389
transform 1 0 4432 0 1 2370
box -8 -3 16 105
use FILL  FILL_5923
timestamp 1677622389
transform 1 0 4440 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_37
timestamp 1677622389
transform -1 0 4480 0 1 2370
box -8 -3 40 105
use FILL  FILL_5924
timestamp 1677622389
transform 1 0 4480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5927
timestamp 1677622389
transform 1 0 4488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5929
timestamp 1677622389
transform 1 0 4496 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4358
timestamp 1677622389
transform 1 0 4516 0 1 2375
box -3 -3 3 3
use FILL  FILL_5931
timestamp 1677622389
transform 1 0 4504 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4359
timestamp 1677622389
transform 1 0 4556 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_224
timestamp 1677622389
transform 1 0 4512 0 1 2370
box -8 -3 46 105
use FILL  FILL_5932
timestamp 1677622389
transform 1 0 4552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5933
timestamp 1677622389
transform 1 0 4560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5934
timestamp 1677622389
transform 1 0 4568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5935
timestamp 1677622389
transform 1 0 4576 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_337
timestamp 1677622389
transform -1 0 4680 0 1 2370
box -8 -3 104 105
use FILL  FILL_5936
timestamp 1677622389
transform 1 0 4680 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_338
timestamp 1677622389
transform 1 0 4688 0 1 2370
box -8 -3 104 105
use FILL  FILL_5943
timestamp 1677622389
transform 1 0 4784 0 1 2370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_47
timestamp 1677622389
transform 1 0 4819 0 1 2370
box -10 -3 10 3
use M2_M1  M2_M1_4916
timestamp 1677622389
transform 1 0 84 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1677622389
transform 1 0 180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1677622389
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4395
timestamp 1677622389
transform 1 0 220 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1677622389
transform 1 0 252 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4919
timestamp 1677622389
transform 1 0 220 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4379
timestamp 1677622389
transform 1 0 316 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1677622389
transform 1 0 412 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1677622389
transform 1 0 332 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4920
timestamp 1677622389
transform 1 0 316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1677622389
transform 1 0 332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1677622389
transform 1 0 132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1677622389
transform 1 0 164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1677622389
transform 1 0 172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1677622389
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1677622389
transform 1 0 204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1677622389
transform 1 0 268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1677622389
transform 1 0 300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1677622389
transform 1 0 308 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4465
timestamp 1677622389
transform 1 0 268 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1677622389
transform 1 0 308 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1677622389
transform 1 0 204 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1677622389
transform 1 0 300 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1677622389
transform 1 0 452 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1677622389
transform 1 0 436 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4922
timestamp 1677622389
transform 1 0 436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1677622389
transform 1 0 444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1677622389
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1677622389
transform 1 0 380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1677622389
transform 1 0 412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1677622389
transform 1 0 420 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1677622389
transform 1 0 436 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4467
timestamp 1677622389
transform 1 0 380 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1677622389
transform 1 0 420 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1677622389
transform 1 0 444 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1677622389
transform 1 0 484 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1677622389
transform 1 0 492 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4925
timestamp 1677622389
transform 1 0 484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1677622389
transform 1 0 500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1677622389
transform 1 0 452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1677622389
transform 1 0 468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1677622389
transform 1 0 492 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4502
timestamp 1677622389
transform 1 0 460 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1677622389
transform 1 0 436 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1677622389
transform 1 0 500 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5015
timestamp 1677622389
transform 1 0 508 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4469
timestamp 1677622389
transform 1 0 492 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1677622389
transform 1 0 516 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1677622389
transform 1 0 508 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4927
timestamp 1677622389
transform 1 0 540 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4471
timestamp 1677622389
transform 1 0 540 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4928
timestamp 1677622389
transform 1 0 604 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4381
timestamp 1677622389
transform 1 0 636 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1677622389
transform 1 0 724 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4929
timestamp 1677622389
transform 1 0 636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1677622389
transform 1 0 588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1677622389
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1677622389
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1677622389
transform 1 0 628 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4503
timestamp 1677622389
transform 1 0 588 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1677622389
transform 1 0 612 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1677622389
transform 1 0 596 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1677622389
transform 1 0 724 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4930
timestamp 1677622389
transform 1 0 724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1677622389
transform 1 0 676 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4504
timestamp 1677622389
transform 1 0 676 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1677622389
transform 1 0 692 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1677622389
transform 1 0 708 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1677622389
transform 1 0 716 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1677622389
transform 1 0 756 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1677622389
transform 1 0 748 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5021
timestamp 1677622389
transform 1 0 780 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4521
timestamp 1677622389
transform 1 0 796 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1677622389
transform 1 0 852 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1677622389
transform 1 0 828 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1677622389
transform 1 0 844 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1677622389
transform 1 0 820 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5022
timestamp 1677622389
transform 1 0 836 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4474
timestamp 1677622389
transform 1 0 836 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5103
timestamp 1677622389
transform 1 0 852 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1677622389
transform 1 0 860 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4403
timestamp 1677622389
transform 1 0 884 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4931
timestamp 1677622389
transform 1 0 884 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4404
timestamp 1677622389
transform 1 0 924 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5023
timestamp 1677622389
transform 1 0 924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1677622389
transform 1 0 996 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1677622389
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1677622389
transform 1 0 1020 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4522
timestamp 1677622389
transform 1 0 1004 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4933
timestamp 1677622389
transform 1 0 1052 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1677622389
transform 1 0 1100 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4383
timestamp 1677622389
transform 1 0 1140 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4935
timestamp 1677622389
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1677622389
transform 1 0 1116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1677622389
transform 1 0 1132 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4363
timestamp 1677622389
transform 1 0 1156 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1677622389
transform 1 0 1156 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5028
timestamp 1677622389
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1677622389
transform 1 0 1180 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4364
timestamp 1677622389
transform 1 0 1284 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4936
timestamp 1677622389
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1677622389
transform 1 0 1300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1677622389
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1677622389
transform 1 0 1348 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4365
timestamp 1677622389
transform 1 0 1388 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5032
timestamp 1677622389
transform 1 0 1548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1677622389
transform 1 0 1660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1677622389
transform 1 0 1612 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4366
timestamp 1677622389
transform 1 0 1676 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1677622389
transform 1 0 1676 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5034
timestamp 1677622389
transform 1 0 1708 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4425
timestamp 1677622389
transform 1 0 1724 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1677622389
transform 1 0 1740 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5035
timestamp 1677622389
transform 1 0 1740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1677622389
transform 1 0 1756 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4530
timestamp 1677622389
transform 1 0 1772 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1677622389
transform 1 0 1788 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1677622389
transform 1 0 1812 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4940
timestamp 1677622389
transform 1 0 1820 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4476
timestamp 1677622389
transform 1 0 1820 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1677622389
transform 1 0 1844 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4941
timestamp 1677622389
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1677622389
transform 1 0 1852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1677622389
transform 1 0 1868 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4477
timestamp 1677622389
transform 1 0 1868 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1677622389
transform 1 0 1884 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1677622389
transform 1 0 1852 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4942
timestamp 1677622389
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4429
timestamp 1677622389
transform 1 0 1908 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5038
timestamp 1677622389
transform 1 0 1908 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4532
timestamp 1677622389
transform 1 0 1916 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5039
timestamp 1677622389
transform 1 0 1932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1677622389
transform 1 0 2020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1677622389
transform 1 0 1996 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4367
timestamp 1677622389
transform 1 0 2036 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4944
timestamp 1677622389
transform 1 0 2036 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4406
timestamp 1677622389
transform 1 0 2068 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5041
timestamp 1677622389
transform 1 0 2100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1677622389
transform 1 0 2124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1677622389
transform 1 0 2140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1677622389
transform 1 0 2156 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4430
timestamp 1677622389
transform 1 0 2180 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1677622389
transform 1 0 2140 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5043
timestamp 1677622389
transform 1 0 2148 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4448
timestamp 1677622389
transform 1 0 2156 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5044
timestamp 1677622389
transform 1 0 2164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1677622389
transform 1 0 2180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1677622389
transform 1 0 2196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1677622389
transform 1 0 2212 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4407
timestamp 1677622389
transform 1 0 2252 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5046
timestamp 1677622389
transform 1 0 2244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1677622389
transform 1 0 2300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1677622389
transform 1 0 2316 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4533
timestamp 1677622389
transform 1 0 2308 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1677622389
transform 1 0 2356 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1677622389
transform 1 0 2348 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1677622389
transform 1 0 2380 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5049
timestamp 1677622389
transform 1 0 2372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1677622389
transform 1 0 2380 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4449
timestamp 1677622389
transform 1 0 2388 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4949
timestamp 1677622389
transform 1 0 2404 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4432
timestamp 1677622389
transform 1 0 2412 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4950
timestamp 1677622389
transform 1 0 2420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1677622389
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4507
timestamp 1677622389
transform 1 0 2396 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1677622389
transform 1 0 2412 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4951
timestamp 1677622389
transform 1 0 2436 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4508
timestamp 1677622389
transform 1 0 2436 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1677622389
transform 1 0 2452 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1677622389
transform 1 0 2460 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5052
timestamp 1677622389
transform 1 0 2468 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4434
timestamp 1677622389
transform 1 0 2508 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5053
timestamp 1677622389
transform 1 0 2500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1677622389
transform 1 0 2508 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4450
timestamp 1677622389
transform 1 0 2532 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1677622389
transform 1 0 2532 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4952
timestamp 1677622389
transform 1 0 2620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1677622389
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4451
timestamp 1677622389
transform 1 0 2580 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1677622389
transform 1 0 2620 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1677622389
transform 1 0 2620 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1677622389
transform 1 0 2684 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1677622389
transform 1 0 2708 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4953
timestamp 1677622389
transform 1 0 2660 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4435
timestamp 1677622389
transform 1 0 2684 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5056
timestamp 1677622389
transform 1 0 2692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1677622389
transform 1 0 2740 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4510
timestamp 1677622389
transform 1 0 2740 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4954
timestamp 1677622389
transform 1 0 2780 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4436
timestamp 1677622389
transform 1 0 2788 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5058
timestamp 1677622389
transform 1 0 2788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1677622389
transform 1 0 2820 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4511
timestamp 1677622389
transform 1 0 2820 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1677622389
transform 1 0 2844 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5059
timestamp 1677622389
transform 1 0 2844 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4437
timestamp 1677622389
transform 1 0 2868 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5060
timestamp 1677622389
transform 1 0 2868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1677622389
transform 1 0 2860 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1677622389
transform 1 0 2892 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4512
timestamp 1677622389
transform 1 0 2908 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1677622389
transform 1 0 2932 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5061
timestamp 1677622389
transform 1 0 2972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1677622389
transform 1 0 2956 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4483
timestamp 1677622389
transform 1 0 2972 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1677622389
transform 1 0 2956 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4957
timestamp 1677622389
transform 1 0 3036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1677622389
transform 1 0 3044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1677622389
transform 1 0 3060 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1677622389
transform 1 0 3052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1677622389
transform 1 0 3068 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4385
timestamp 1677622389
transform 1 0 3092 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4960
timestamp 1677622389
transform 1 0 3092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1677622389
transform 1 0 3084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1677622389
transform 1 0 3108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1677622389
transform 1 0 3124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1677622389
transform 1 0 3148 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4452
timestamp 1677622389
transform 1 0 3148 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4963
timestamp 1677622389
transform 1 0 3164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1677622389
transform 1 0 3156 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4453
timestamp 1677622389
transform 1 0 3164 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5067
timestamp 1677622389
transform 1 0 3180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1677622389
transform 1 0 3196 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4484
timestamp 1677622389
transform 1 0 3196 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1677622389
transform 1 0 3228 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4964
timestamp 1677622389
transform 1 0 3228 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4485
timestamp 1677622389
transform 1 0 3228 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1677622389
transform 1 0 3284 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1677622389
transform 1 0 3300 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4965
timestamp 1677622389
transform 1 0 3252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1677622389
transform 1 0 3300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1677622389
transform 1 0 3364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1677622389
transform 1 0 3356 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4454
timestamp 1677622389
transform 1 0 3364 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1677622389
transform 1 0 3356 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1677622389
transform 1 0 3380 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1677622389
transform 1 0 3420 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4967
timestamp 1677622389
transform 1 0 3404 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4438
timestamp 1677622389
transform 1 0 3412 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1677622389
transform 1 0 3444 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4968
timestamp 1677622389
transform 1 0 3420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1677622389
transform 1 0 3436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1677622389
transform 1 0 3444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1677622389
transform 1 0 3412 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4487
timestamp 1677622389
transform 1 0 3412 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1677622389
transform 1 0 3516 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1677622389
transform 1 0 3508 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4971
timestamp 1677622389
transform 1 0 3492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1677622389
transform 1 0 3508 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4439
timestamp 1677622389
transform 1 0 3516 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4973
timestamp 1677622389
transform 1 0 3524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1677622389
transform 1 0 3500 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4455
timestamp 1677622389
transform 1 0 3508 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5073
timestamp 1677622389
transform 1 0 3516 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4488
timestamp 1677622389
transform 1 0 3492 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1677622389
transform 1 0 3516 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1677622389
transform 1 0 3532 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1677622389
transform 1 0 3556 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1677622389
transform 1 0 3604 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4974
timestamp 1677622389
transform 1 0 3580 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4456
timestamp 1677622389
transform 1 0 3580 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5074
timestamp 1677622389
transform 1 0 3604 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4457
timestamp 1677622389
transform 1 0 3644 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1677622389
transform 1 0 3604 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1677622389
transform 1 0 3668 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5075
timestamp 1677622389
transform 1 0 3684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4490
timestamp 1677622389
transform 1 0 3692 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1677622389
transform 1 0 3684 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1677622389
transform 1 0 3740 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4975
timestamp 1677622389
transform 1 0 3716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1677622389
transform 1 0 3740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1677622389
transform 1 0 3796 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4491
timestamp 1677622389
transform 1 0 3740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1677622389
transform 1 0 3772 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1677622389
transform 1 0 3796 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1677622389
transform 1 0 3844 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4976
timestamp 1677622389
transform 1 0 3836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1677622389
transform 1 0 3828 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1677622389
transform 1 0 3852 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4458
timestamp 1677622389
transform 1 0 3852 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1677622389
transform 1 0 3892 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5079
timestamp 1677622389
transform 1 0 3860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1677622389
transform 1 0 3876 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4459
timestamp 1677622389
transform 1 0 3884 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1677622389
transform 1 0 3876 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1677622389
transform 1 0 3932 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1677622389
transform 1 0 3956 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4978
timestamp 1677622389
transform 1 0 3916 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1677622389
transform 1 0 3924 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4440
timestamp 1677622389
transform 1 0 3932 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4980
timestamp 1677622389
transform 1 0 3940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1677622389
transform 1 0 3956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1677622389
transform 1 0 3924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1677622389
transform 1 0 3932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1677622389
transform 1 0 3948 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4492
timestamp 1677622389
transform 1 0 3916 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1677622389
transform 1 0 3948 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5084
timestamp 1677622389
transform 1 0 3964 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4494
timestamp 1677622389
transform 1 0 3964 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1677622389
transform 1 0 3980 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1677622389
transform 1 0 3996 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4982
timestamp 1677622389
transform 1 0 4020 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4374
timestamp 1677622389
transform 1 0 4100 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1677622389
transform 1 0 4108 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1677622389
transform 1 0 4132 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1677622389
transform 1 0 4172 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1677622389
transform 1 0 4172 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1677622389
transform 1 0 4132 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1677622389
transform 1 0 4148 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1677622389
transform 1 0 4196 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4983
timestamp 1677622389
transform 1 0 4132 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4441
timestamp 1677622389
transform 1 0 4180 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1677622389
transform 1 0 4132 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5085
timestamp 1677622389
transform 1 0 4156 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4495
timestamp 1677622389
transform 1 0 4164 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1677622389
transform 1 0 4244 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1677622389
transform 1 0 4252 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5086
timestamp 1677622389
transform 1 0 4244 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4496
timestamp 1677622389
transform 1 0 4244 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4984
timestamp 1677622389
transform 1 0 4260 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4391
timestamp 1677622389
transform 1 0 4308 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4985
timestamp 1677622389
transform 1 0 4292 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4442
timestamp 1677622389
transform 1 0 4300 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5087
timestamp 1677622389
transform 1 0 4284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1677622389
transform 1 0 4300 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4497
timestamp 1677622389
transform 1 0 4284 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1677622389
transform 1 0 4332 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4986
timestamp 1677622389
transform 1 0 4340 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4540
timestamp 1677622389
transform 1 0 4348 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4987
timestamp 1677622389
transform 1 0 4364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1677622389
transform 1 0 4372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1677622389
transform 1 0 4388 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4498
timestamp 1677622389
transform 1 0 4364 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4988
timestamp 1677622389
transform 1 0 4420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1677622389
transform 1 0 4412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1677622389
transform 1 0 4412 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1677622389
transform 1 0 4428 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1677622389
transform 1 0 4460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1677622389
transform 1 0 4484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1677622389
transform 1 0 4476 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4516
timestamp 1677622389
transform 1 0 4460 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1677622389
transform 1 0 4548 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1677622389
transform 1 0 4540 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4989
timestamp 1677622389
transform 1 0 4516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1677622389
transform 1 0 4540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1677622389
transform 1 0 4548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1677622389
transform 1 0 4564 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4461
timestamp 1677622389
transform 1 0 4516 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1677622389
transform 1 0 4572 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4993
timestamp 1677622389
transform 1 0 4580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1677622389
transform 1 0 4524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1677622389
transform 1 0 4548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1677622389
transform 1 0 4556 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4517
timestamp 1677622389
transform 1 0 4532 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1677622389
transform 1 0 4564 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5097
timestamp 1677622389
transform 1 0 4572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1677622389
transform 1 0 4588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1677622389
transform 1 0 4604 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4377
timestamp 1677622389
transform 1 0 4628 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1677622389
transform 1 0 4628 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1677622389
transform 1 0 4660 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1677622389
transform 1 0 4652 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4994
timestamp 1677622389
transform 1 0 4620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1677622389
transform 1 0 4628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1677622389
transform 1 0 4644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1677622389
transform 1 0 4660 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4463
timestamp 1677622389
transform 1 0 4620 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1677622389
transform 1 0 4620 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5100
timestamp 1677622389
transform 1 0 4636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1677622389
transform 1 0 4652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1677622389
transform 1 0 4668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1677622389
transform 1 0 4676 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4444
timestamp 1677622389
transform 1 0 4700 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1677622389
transform 1 0 4756 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4999
timestamp 1677622389
transform 1 0 4780 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4500
timestamp 1677622389
transform 1 0 4796 0 1 2315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_48
timestamp 1677622389
transform 1 0 24 0 1 2270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_317
timestamp 1677622389
transform 1 0 72 0 -1 2370
box -8 -3 104 105
use AOI22X1  AOI22X1_215
timestamp 1677622389
transform -1 0 208 0 -1 2370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_318
timestamp 1677622389
transform 1 0 208 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_363
timestamp 1677622389
transform -1 0 320 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_319
timestamp 1677622389
transform 1 0 320 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_364
timestamp 1677622389
transform -1 0 432 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_216
timestamp 1677622389
transform 1 0 432 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1677622389
transform -1 0 512 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5432
timestamp 1677622389
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5433
timestamp 1677622389
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5434
timestamp 1677622389
transform 1 0 528 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_365
timestamp 1677622389
transform 1 0 536 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5438
timestamp 1677622389
transform 1 0 552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5450
timestamp 1677622389
transform 1 0 560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5451
timestamp 1677622389
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5452
timestamp 1677622389
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5453
timestamp 1677622389
transform 1 0 584 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_219
timestamp 1677622389
transform 1 0 592 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5454
timestamp 1677622389
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_320
timestamp 1677622389
transform -1 0 736 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5455
timestamp 1677622389
transform 1 0 736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5457
timestamp 1677622389
transform 1 0 744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5459
timestamp 1677622389
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5461
timestamp 1677622389
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5462
timestamp 1677622389
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5463
timestamp 1677622389
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5464
timestamp 1677622389
transform 1 0 784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5465
timestamp 1677622389
transform 1 0 792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5467
timestamp 1677622389
transform 1 0 800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5469
timestamp 1677622389
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5471
timestamp 1677622389
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_109
timestamp 1677622389
transform 1 0 824 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5474
timestamp 1677622389
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5475
timestamp 1677622389
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5476
timestamp 1677622389
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5477
timestamp 1677622389
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5478
timestamp 1677622389
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_54
timestamp 1677622389
transform 1 0 896 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5479
timestamp 1677622389
transform 1 0 920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5480
timestamp 1677622389
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5482
timestamp 1677622389
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5484
timestamp 1677622389
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5486
timestamp 1677622389
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5488
timestamp 1677622389
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5490
timestamp 1677622389
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5493
timestamp 1677622389
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_221
timestamp 1677622389
transform 1 0 984 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5494
timestamp 1677622389
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5496
timestamp 1677622389
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5498
timestamp 1677622389
transform 1 0 1040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5500
timestamp 1677622389
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5502
timestamp 1677622389
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5504
timestamp 1677622389
transform 1 0 1064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5506
timestamp 1677622389
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5508
timestamp 1677622389
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5513
timestamp 1677622389
transform 1 0 1088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5514
timestamp 1677622389
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5515
timestamp 1677622389
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_223
timestamp 1677622389
transform 1 0 1112 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5516
timestamp 1677622389
transform 1 0 1152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5518
timestamp 1677622389
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5520
timestamp 1677622389
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5522
timestamp 1677622389
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5524
timestamp 1677622389
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5526
timestamp 1677622389
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5529
timestamp 1677622389
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_53
timestamp 1677622389
transform 1 0 1208 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5530
timestamp 1677622389
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5531
timestamp 1677622389
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5533
timestamp 1677622389
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5535
timestamp 1677622389
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5537
timestamp 1677622389
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5539
timestamp 1677622389
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5541
timestamp 1677622389
transform 1 0 1280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5543
timestamp 1677622389
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5545
timestamp 1677622389
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5548
timestamp 1677622389
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_367
timestamp 1677622389
transform -1 0 1328 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5549
timestamp 1677622389
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5550
timestamp 1677622389
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5551
timestamp 1677622389
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5553
timestamp 1677622389
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5555
timestamp 1677622389
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5557
timestamp 1677622389
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5559
timestamp 1677622389
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5561
timestamp 1677622389
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5562
timestamp 1677622389
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5563
timestamp 1677622389
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5564
timestamp 1677622389
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5565
timestamp 1677622389
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5566
timestamp 1677622389
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5567
timestamp 1677622389
transform 1 0 1432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5568
timestamp 1677622389
transform 1 0 1440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5569
timestamp 1677622389
transform 1 0 1448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5570
timestamp 1677622389
transform 1 0 1456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5571
timestamp 1677622389
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5572
timestamp 1677622389
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5573
timestamp 1677622389
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5575
timestamp 1677622389
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5577
timestamp 1677622389
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4541
timestamp 1677622389
transform 1 0 1516 0 1 2275
box -3 -3 3 3
use FILL  FILL_5579
timestamp 1677622389
transform 1 0 1504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5580
timestamp 1677622389
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5581
timestamp 1677622389
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5583
timestamp 1677622389
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5588
timestamp 1677622389
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_369
timestamp 1677622389
transform -1 0 1560 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5589
timestamp 1677622389
transform 1 0 1560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5599
timestamp 1677622389
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_324
timestamp 1677622389
transform -1 0 1672 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5600
timestamp 1677622389
transform 1 0 1672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5601
timestamp 1677622389
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5602
timestamp 1677622389
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5603
timestamp 1677622389
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5604
timestamp 1677622389
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4542
timestamp 1677622389
transform 1 0 1724 0 1 2275
box -3 -3 3 3
use FILL  FILL_5605
timestamp 1677622389
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5606
timestamp 1677622389
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_370
timestamp 1677622389
transform -1 0 1744 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5607
timestamp 1677622389
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5608
timestamp 1677622389
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4543
timestamp 1677622389
transform 1 0 1772 0 1 2275
box -3 -3 3 3
use FILL  FILL_5609
timestamp 1677622389
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5610
timestamp 1677622389
transform 1 0 1768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5612
timestamp 1677622389
transform 1 0 1776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5622
timestamp 1677622389
transform 1 0 1784 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_371
timestamp 1677622389
transform -1 0 1808 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5623
timestamp 1677622389
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5624
timestamp 1677622389
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5625
timestamp 1677622389
transform 1 0 1824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5626
timestamp 1677622389
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5627
timestamp 1677622389
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_225
timestamp 1677622389
transform 1 0 1848 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5628
timestamp 1677622389
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5630
timestamp 1677622389
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5632
timestamp 1677622389
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5634
timestamp 1677622389
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5645
timestamp 1677622389
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5646
timestamp 1677622389
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_325
timestamp 1677622389
transform -1 0 2032 0 -1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4544
timestamp 1677622389
transform 1 0 2044 0 1 2275
box -3 -3 3 3
use FILL  FILL_5647
timestamp 1677622389
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5652
timestamp 1677622389
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5653
timestamp 1677622389
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4545
timestamp 1677622389
transform 1 0 2068 0 1 2275
box -3 -3 3 3
use FILL  FILL_5654
timestamp 1677622389
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5655
timestamp 1677622389
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5656
timestamp 1677622389
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_54
timestamp 1677622389
transform -1 0 2104 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5657
timestamp 1677622389
transform 1 0 2104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5659
timestamp 1677622389
transform 1 0 2112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5665
timestamp 1677622389
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_372
timestamp 1677622389
transform -1 0 2144 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_228
timestamp 1677622389
transform 1 0 2144 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5666
timestamp 1677622389
transform 1 0 2184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5667
timestamp 1677622389
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5669
timestamp 1677622389
transform 1 0 2200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5671
timestamp 1677622389
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5673
timestamp 1677622389
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5675
timestamp 1677622389
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5677
timestamp 1677622389
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_373
timestamp 1677622389
transform 1 0 2240 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5681
timestamp 1677622389
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5683
timestamp 1677622389
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5685
timestamp 1677622389
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5687
timestamp 1677622389
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5690
timestamp 1677622389
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use AND2X2  AND2X2_12
timestamp 1677622389
transform -1 0 2328 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5691
timestamp 1677622389
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5692
timestamp 1677622389
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5694
timestamp 1677622389
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5696
timestamp 1677622389
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5698
timestamp 1677622389
transform 1 0 2360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5700
timestamp 1677622389
transform 1 0 2368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5702
timestamp 1677622389
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5710
timestamp 1677622389
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_230
timestamp 1677622389
transform -1 0 2432 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5711
timestamp 1677622389
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5713
timestamp 1677622389
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5715
timestamp 1677622389
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5717
timestamp 1677622389
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_374
timestamp 1677622389
transform 1 0 2464 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5721
timestamp 1677622389
transform 1 0 2480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5723
timestamp 1677622389
transform 1 0 2488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5725
timestamp 1677622389
transform 1 0 2496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5727
timestamp 1677622389
transform 1 0 2504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5728
timestamp 1677622389
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5729
timestamp 1677622389
transform 1 0 2520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5749
timestamp 1677622389
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4546
timestamp 1677622389
transform 1 0 2548 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_326
timestamp 1677622389
transform -1 0 2632 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5750
timestamp 1677622389
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5751
timestamp 1677622389
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_327
timestamp 1677622389
transform 1 0 2648 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5752
timestamp 1677622389
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5754
timestamp 1677622389
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5755
timestamp 1677622389
transform 1 0 2760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5756
timestamp 1677622389
transform 1 0 2768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5757
timestamp 1677622389
transform 1 0 2776 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_112
timestamp 1677622389
transform 1 0 2784 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5758
timestamp 1677622389
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5759
timestamp 1677622389
transform 1 0 2824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5760
timestamp 1677622389
transform 1 0 2832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5761
timestamp 1677622389
transform 1 0 2840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5762
timestamp 1677622389
transform 1 0 2848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5764
timestamp 1677622389
transform 1 0 2856 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_113
timestamp 1677622389
transform 1 0 2864 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5767
timestamp 1677622389
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5769
timestamp 1677622389
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5771
timestamp 1677622389
transform 1 0 2912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5773
timestamp 1677622389
transform 1 0 2920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5777
timestamp 1677622389
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5778
timestamp 1677622389
transform 1 0 2936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5779
timestamp 1677622389
transform 1 0 2944 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1677622389
transform -1 0 2984 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5780
timestamp 1677622389
transform 1 0 2984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5781
timestamp 1677622389
transform 1 0 2992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5782
timestamp 1677622389
transform 1 0 3000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5783
timestamp 1677622389
transform 1 0 3008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5784
timestamp 1677622389
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5785
timestamp 1677622389
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5786
timestamp 1677622389
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_215
timestamp 1677622389
transform -1 0 3080 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5787
timestamp 1677622389
transform 1 0 3080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5788
timestamp 1677622389
transform 1 0 3088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5789
timestamp 1677622389
transform 1 0 3096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5791
timestamp 1677622389
transform 1 0 3104 0 -1 2370
box -8 -3 16 105
use AND2X2  AND2X2_13
timestamp 1677622389
transform 1 0 3112 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5806
timestamp 1677622389
transform 1 0 3144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5807
timestamp 1677622389
transform 1 0 3152 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_58
timestamp 1677622389
transform -1 0 3184 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5808
timestamp 1677622389
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_59
timestamp 1677622389
transform 1 0 3192 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5809
timestamp 1677622389
transform 1 0 3216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5810
timestamp 1677622389
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5811
timestamp 1677622389
transform 1 0 3232 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_330
timestamp 1677622389
transform 1 0 3240 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5812
timestamp 1677622389
transform 1 0 3336 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_380
timestamp 1677622389
transform 1 0 3344 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5821
timestamp 1677622389
transform 1 0 3360 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4547
timestamp 1677622389
transform 1 0 3380 0 1 2275
box -3 -3 3 3
use FILL  FILL_5822
timestamp 1677622389
transform 1 0 3368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5823
timestamp 1677622389
transform 1 0 3376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5824
timestamp 1677622389
transform 1 0 3384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5825
timestamp 1677622389
transform 1 0 3392 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_216
timestamp 1677622389
transform -1 0 3440 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5826
timestamp 1677622389
transform 1 0 3440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5827
timestamp 1677622389
transform 1 0 3448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5828
timestamp 1677622389
transform 1 0 3456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5829
timestamp 1677622389
transform 1 0 3464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5831
timestamp 1677622389
transform 1 0 3472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5833
timestamp 1677622389
transform 1 0 3480 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_217
timestamp 1677622389
transform 1 0 3488 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5837
timestamp 1677622389
transform 1 0 3528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5838
timestamp 1677622389
transform 1 0 3536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5839
timestamp 1677622389
transform 1 0 3544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5841
timestamp 1677622389
transform 1 0 3552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5843
timestamp 1677622389
transform 1 0 3560 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_331
timestamp 1677622389
transform 1 0 3568 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5850
timestamp 1677622389
transform 1 0 3664 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_382
timestamp 1677622389
transform 1 0 3672 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5856
timestamp 1677622389
transform 1 0 3688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5857
timestamp 1677622389
transform 1 0 3696 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4548
timestamp 1677622389
transform 1 0 3788 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_333
timestamp 1677622389
transform 1 0 3704 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5858
timestamp 1677622389
transform 1 0 3800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5860
timestamp 1677622389
transform 1 0 3808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5864
timestamp 1677622389
transform 1 0 3816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5865
timestamp 1677622389
transform 1 0 3824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5866
timestamp 1677622389
transform 1 0 3832 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_234
timestamp 1677622389
transform 1 0 3840 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5867
timestamp 1677622389
transform 1 0 3880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5868
timestamp 1677622389
transform 1 0 3888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5869
timestamp 1677622389
transform 1 0 3896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5871
timestamp 1677622389
transform 1 0 3904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5873
timestamp 1677622389
transform 1 0 3912 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_220
timestamp 1677622389
transform 1 0 3920 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5876
timestamp 1677622389
transform 1 0 3960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5877
timestamp 1677622389
transform 1 0 3968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5880
timestamp 1677622389
transform 1 0 3976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5881
timestamp 1677622389
transform 1 0 3984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5882
timestamp 1677622389
transform 1 0 3992 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_385
timestamp 1677622389
transform -1 0 4016 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5883
timestamp 1677622389
transform 1 0 4016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5884
timestamp 1677622389
transform 1 0 4024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5885
timestamp 1677622389
transform 1 0 4032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5886
timestamp 1677622389
transform 1 0 4040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5887
timestamp 1677622389
transform 1 0 4048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5888
timestamp 1677622389
transform 1 0 4056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5889
timestamp 1677622389
transform 1 0 4064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5890
timestamp 1677622389
transform 1 0 4072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5891
timestamp 1677622389
transform 1 0 4080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5892
timestamp 1677622389
transform 1 0 4088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5893
timestamp 1677622389
transform 1 0 4096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5894
timestamp 1677622389
transform 1 0 4104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5895
timestamp 1677622389
transform 1 0 4112 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_336
timestamp 1677622389
transform 1 0 4120 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5901
timestamp 1677622389
transform 1 0 4216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5902
timestamp 1677622389
transform 1 0 4224 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_387
timestamp 1677622389
transform 1 0 4232 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5903
timestamp 1677622389
transform 1 0 4248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5904
timestamp 1677622389
transform 1 0 4256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5905
timestamp 1677622389
transform 1 0 4264 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_223
timestamp 1677622389
transform -1 0 4312 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5906
timestamp 1677622389
transform 1 0 4312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5907
timestamp 1677622389
transform 1 0 4320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5908
timestamp 1677622389
transform 1 0 4328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5909
timestamp 1677622389
transform 1 0 4336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5910
timestamp 1677622389
transform 1 0 4344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5912
timestamp 1677622389
transform 1 0 4352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5916
timestamp 1677622389
transform 1 0 4360 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_236
timestamp 1677622389
transform -1 0 4408 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5917
timestamp 1677622389
transform 1 0 4408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5918
timestamp 1677622389
transform 1 0 4416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5920
timestamp 1677622389
transform 1 0 4424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5922
timestamp 1677622389
transform 1 0 4432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5925
timestamp 1677622389
transform 1 0 4440 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_38
timestamp 1677622389
transform 1 0 4448 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5926
timestamp 1677622389
transform 1 0 4480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5928
timestamp 1677622389
transform 1 0 4488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5930
timestamp 1677622389
transform 1 0 4496 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_237
timestamp 1677622389
transform 1 0 4504 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_225
timestamp 1677622389
transform 1 0 4544 0 -1 2370
box -8 -3 46 105
use INVX2  INVX2_388
timestamp 1677622389
transform -1 0 4600 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5937
timestamp 1677622389
transform 1 0 4600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5938
timestamp 1677622389
transform 1 0 4608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5939
timestamp 1677622389
transform 1 0 4616 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_226
timestamp 1677622389
transform 1 0 4624 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5940
timestamp 1677622389
transform 1 0 4664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5941
timestamp 1677622389
transform 1 0 4672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5942
timestamp 1677622389
transform 1 0 4680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5944
timestamp 1677622389
transform 1 0 4688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5945
timestamp 1677622389
transform 1 0 4696 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_389
timestamp 1677622389
transform -1 0 4720 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5946
timestamp 1677622389
transform 1 0 4720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5947
timestamp 1677622389
transform 1 0 4728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5948
timestamp 1677622389
transform 1 0 4736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5949
timestamp 1677622389
transform 1 0 4744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5950
timestamp 1677622389
transform 1 0 4752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5951
timestamp 1677622389
transform 1 0 4760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5952
timestamp 1677622389
transform 1 0 4768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5953
timestamp 1677622389
transform 1 0 4776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5954
timestamp 1677622389
transform 1 0 4784 0 -1 2370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_49
timestamp 1677622389
transform 1 0 4843 0 1 2270
box -10 -3 10 3
use M3_M2  M3_M2_4580
timestamp 1677622389
transform 1 0 164 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1677622389
transform 1 0 132 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1677622389
transform 1 0 172 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1677622389
transform 1 0 84 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5125
timestamp 1677622389
transform 1 0 132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1677622389
transform 1 0 164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1677622389
transform 1 0 172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1677622389
transform 1 0 84 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4581
timestamp 1677622389
transform 1 0 196 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5128
timestamp 1677622389
transform 1 0 180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1677622389
transform 1 0 204 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4629
timestamp 1677622389
transform 1 0 236 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5130
timestamp 1677622389
transform 1 0 276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1677622389
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1677622389
transform 1 0 196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1677622389
transform 1 0 212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1677622389
transform 1 0 220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1677622389
transform 1 0 236 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4662
timestamp 1677622389
transform 1 0 180 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1677622389
transform 1 0 236 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5131
timestamp 1677622389
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4630
timestamp 1677622389
transform 1 0 332 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5230
timestamp 1677622389
transform 1 0 372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1677622389
transform 1 0 404 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4562
timestamp 1677622389
transform 1 0 428 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5132
timestamp 1677622389
transform 1 0 420 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4640
timestamp 1677622389
transform 1 0 420 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1677622389
transform 1 0 468 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1677622389
transform 1 0 468 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1677622389
transform 1 0 524 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1677622389
transform 1 0 500 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1677622389
transform 1 0 540 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5133
timestamp 1677622389
transform 1 0 468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1677622389
transform 1 0 476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1677622389
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1677622389
transform 1 0 508 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1677622389
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1677622389
transform 1 0 460 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4631
timestamp 1677622389
transform 1 0 588 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5138
timestamp 1677622389
transform 1 0 604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1677622389
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1677622389
transform 1 0 500 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1677622389
transform 1 0 588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4664
timestamp 1677622389
transform 1 0 484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1677622389
transform 1 0 548 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1677622389
transform 1 0 628 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1677622389
transform 1 0 636 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1677622389
transform 1 0 620 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1677622389
transform 1 0 660 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1677622389
transform 1 0 660 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5139
timestamp 1677622389
transform 1 0 660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1677622389
transform 1 0 628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1677622389
transform 1 0 636 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4642
timestamp 1677622389
transform 1 0 652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1677622389
transform 1 0 660 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5315
timestamp 1677622389
transform 1 0 668 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1677622389
transform 1 0 708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1677622389
transform 1 0 716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1677622389
transform 1 0 732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1677622389
transform 1 0 756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1677622389
transform 1 0 772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1677622389
transform 1 0 748 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4643
timestamp 1677622389
transform 1 0 756 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5240
timestamp 1677622389
transform 1 0 780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1677622389
transform 1 0 852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1677622389
transform 1 0 828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1677622389
transform 1 0 932 0 1 2245
box -2 -2 2 2
use M3_M2  M3_M2_4583
timestamp 1677622389
transform 1 0 932 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1677622389
transform 1 0 924 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5145
timestamp 1677622389
transform 1 0 940 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4666
timestamp 1677622389
transform 1 0 940 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5110
timestamp 1677622389
transform 1 0 956 0 1 2245
box -2 -2 2 2
use M3_M2  M3_M2_4584
timestamp 1677622389
transform 1 0 964 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5146
timestamp 1677622389
transform 1 0 980 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4634
timestamp 1677622389
transform 1 0 996 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5242
timestamp 1677622389
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1677622389
transform 1 0 972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1677622389
transform 1 0 996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1677622389
transform 1 0 1004 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4667
timestamp 1677622389
transform 1 0 996 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5147
timestamp 1677622389
transform 1 0 1020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1677622389
transform 1 0 1012 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4697
timestamp 1677622389
transform 1 0 1012 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5246
timestamp 1677622389
transform 1 0 1060 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4668
timestamp 1677622389
transform 1 0 1060 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1677622389
transform 1 0 1124 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5148
timestamp 1677622389
transform 1 0 1140 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4669
timestamp 1677622389
transform 1 0 1140 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5149
timestamp 1677622389
transform 1 0 1156 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4606
timestamp 1677622389
transform 1 0 1180 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5247
timestamp 1677622389
transform 1 0 1180 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4670
timestamp 1677622389
transform 1 0 1180 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1677622389
transform 1 0 1244 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5120
timestamp 1677622389
transform 1 0 1252 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4585
timestamp 1677622389
transform 1 0 1284 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1677622389
transform 1 0 1300 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5150
timestamp 1677622389
transform 1 0 1308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1677622389
transform 1 0 1300 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4586
timestamp 1677622389
transform 1 0 1428 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5151
timestamp 1677622389
transform 1 0 1348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1677622389
transform 1 0 1404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1677622389
transform 1 0 1428 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4671
timestamp 1677622389
transform 1 0 1404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1677622389
transform 1 0 1444 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1677622389
transform 1 0 1468 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5250
timestamp 1677622389
transform 1 0 1468 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4608
timestamp 1677622389
transform 1 0 1484 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5153
timestamp 1677622389
transform 1 0 1484 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4644
timestamp 1677622389
transform 1 0 1484 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5251
timestamp 1677622389
transform 1 0 1492 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4672
timestamp 1677622389
transform 1 0 1492 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5154
timestamp 1677622389
transform 1 0 1516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1677622389
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4555
timestamp 1677622389
transform 1 0 1580 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1677622389
transform 1 0 1620 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1677622389
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5155
timestamp 1677622389
transform 1 0 1556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1677622389
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4645
timestamp 1677622389
transform 1 0 1596 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5253
timestamp 1677622389
transform 1 0 1636 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4549
timestamp 1677622389
transform 1 0 1668 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1677622389
transform 1 0 1660 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5254
timestamp 1677622389
transform 1 0 1692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1677622389
transform 1 0 1708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1677622389
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1677622389
transform 1 0 1716 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1677622389
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1677622389
transform 1 0 1900 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4587
timestamp 1677622389
transform 1 0 1940 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1677622389
transform 1 0 1932 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5159
timestamp 1677622389
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1677622389
transform 1 0 1948 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4612
timestamp 1677622389
transform 1 0 1964 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5258
timestamp 1677622389
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1677622389
transform 1 0 1956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1677622389
transform 1 0 1996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1677622389
transform 1 0 2052 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4699
timestamp 1677622389
transform 1 0 2076 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1677622389
transform 1 0 2204 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1677622389
transform 1 0 2188 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1677622389
transform 1 0 2228 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5162
timestamp 1677622389
transform 1 0 2092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1677622389
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1677622389
transform 1 0 2188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1677622389
transform 1 0 2244 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4646
timestamp 1677622389
transform 1 0 2092 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5261
timestamp 1677622389
transform 1 0 2172 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4647
timestamp 1677622389
transform 1 0 2188 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5262
timestamp 1677622389
transform 1 0 2268 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4673
timestamp 1677622389
transform 1 0 2172 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1677622389
transform 1 0 2268 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1677622389
transform 1 0 2220 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1677622389
transform 1 0 2252 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1677622389
transform 1 0 2292 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1677622389
transform 1 0 2300 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1677622389
transform 1 0 2372 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1677622389
transform 1 0 2404 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5166
timestamp 1677622389
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1677622389
transform 1 0 2396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1677622389
transform 1 0 2388 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4648
timestamp 1677622389
transform 1 0 2396 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5264
timestamp 1677622389
transform 1 0 2404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1677622389
transform 1 0 2428 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4649
timestamp 1677622389
transform 1 0 2428 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5317
timestamp 1677622389
transform 1 0 2428 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4702
timestamp 1677622389
transform 1 0 2444 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1677622389
transform 1 0 2492 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5169
timestamp 1677622389
transform 1 0 2500 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4650
timestamp 1677622389
transform 1 0 2460 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5265
timestamp 1677622389
transform 1 0 2532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4675
timestamp 1677622389
transform 1 0 2532 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1677622389
transform 1 0 2468 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1677622389
transform 1 0 2532 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5111
timestamp 1677622389
transform 1 0 2556 0 1 2245
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1677622389
transform 1 0 2548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1677622389
transform 1 0 2588 0 1 2245
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1677622389
transform 1 0 2588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1677622389
transform 1 0 2612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1677622389
transform 1 0 2636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1677622389
transform 1 0 2604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1677622389
transform 1 0 2620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1677622389
transform 1 0 2628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1677622389
transform 1 0 2660 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4651
timestamp 1677622389
transform 1 0 2652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1677622389
transform 1 0 2668 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5174
timestamp 1677622389
transform 1 0 2692 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4592
timestamp 1677622389
transform 1 0 2828 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1677622389
transform 1 0 2820 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5175
timestamp 1677622389
transform 1 0 2756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1677622389
transform 1 0 2812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1677622389
transform 1 0 2732 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4652
timestamp 1677622389
transform 1 0 2780 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1677622389
transform 1 0 2812 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1677622389
transform 1 0 2732 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5318
timestamp 1677622389
transform 1 0 2820 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4705
timestamp 1677622389
transform 1 0 2828 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5177
timestamp 1677622389
transform 1 0 2844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1677622389
transform 1 0 2844 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4706
timestamp 1677622389
transform 1 0 2844 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5272
timestamp 1677622389
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1677622389
transform 1 0 2892 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1677622389
transform 1 0 2908 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1677622389
transform 1 0 2932 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4557
timestamp 1677622389
transform 1 0 2988 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1677622389
transform 1 0 2980 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5273
timestamp 1677622389
transform 1 0 2988 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4678
timestamp 1677622389
transform 1 0 2988 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1677622389
transform 1 0 3004 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5179
timestamp 1677622389
transform 1 0 3052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1677622389
transform 1 0 3084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1677622389
transform 1 0 3004 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4679
timestamp 1677622389
transform 1 0 3020 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1677622389
transform 1 0 3044 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1677622389
transform 1 0 3108 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1677622389
transform 1 0 3100 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1677622389
transform 1 0 3124 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1677622389
transform 1 0 3188 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5275
timestamp 1677622389
transform 1 0 3188 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4550
timestamp 1677622389
transform 1 0 3228 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1677622389
transform 1 0 3220 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5181
timestamp 1677622389
transform 1 0 3220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1677622389
transform 1 0 3228 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4615
timestamp 1677622389
transform 1 0 3268 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5183
timestamp 1677622389
transform 1 0 3252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1677622389
transform 1 0 3244 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4681
timestamp 1677622389
transform 1 0 3244 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5277
timestamp 1677622389
transform 1 0 3268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1677622389
transform 1 0 3284 0 1 2245
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1677622389
transform 1 0 3284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1677622389
transform 1 0 3324 0 1 2245
box -2 -2 2 2
use M3_M2  M3_M2_4616
timestamp 1677622389
transform 1 0 3316 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5278
timestamp 1677622389
transform 1 0 3316 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4594
timestamp 1677622389
transform 1 0 3364 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5185
timestamp 1677622389
transform 1 0 3348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1677622389
transform 1 0 3364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1677622389
transform 1 0 3356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1677622389
transform 1 0 3372 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4682
timestamp 1677622389
transform 1 0 3380 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1677622389
transform 1 0 3436 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5187
timestamp 1677622389
transform 1 0 3420 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4655
timestamp 1677622389
transform 1 0 3420 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1677622389
transform 1 0 3444 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5281
timestamp 1677622389
transform 1 0 3460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1677622389
transform 1 0 3476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1677622389
transform 1 0 3484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1677622389
transform 1 0 3500 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4656
timestamp 1677622389
transform 1 0 3476 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5282
timestamp 1677622389
transform 1 0 3492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1677622389
transform 1 0 3508 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4683
timestamp 1677622389
transform 1 0 3492 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5115
timestamp 1677622389
transform 1 0 3524 0 1 2245
box -2 -2 2 2
use M3_M2  M3_M2_4560
timestamp 1677622389
transform 1 0 3540 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1677622389
transform 1 0 3532 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5191
timestamp 1677622389
transform 1 0 3532 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4657
timestamp 1677622389
transform 1 0 3524 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5116
timestamp 1677622389
transform 1 0 3580 0 1 2245
box -2 -2 2 2
use M3_M2  M3_M2_4684
timestamp 1677622389
transform 1 0 3580 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5192
timestamp 1677622389
transform 1 0 3596 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4685
timestamp 1677622389
transform 1 0 3596 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5193
timestamp 1677622389
transform 1 0 3628 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4574
timestamp 1677622389
transform 1 0 3644 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5284
timestamp 1677622389
transform 1 0 3636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1677622389
transform 1 0 3644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1677622389
transform 1 0 3660 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4658
timestamp 1677622389
transform 1 0 3660 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1677622389
transform 1 0 3700 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5195
timestamp 1677622389
transform 1 0 3700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1677622389
transform 1 0 3716 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4618
timestamp 1677622389
transform 1 0 3716 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5196
timestamp 1677622389
transform 1 0 3716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1677622389
transform 1 0 3676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1677622389
transform 1 0 3692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1677622389
transform 1 0 3708 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4686
timestamp 1677622389
transform 1 0 3708 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1677622389
transform 1 0 3748 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5118
timestamp 1677622389
transform 1 0 3740 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4619
timestamp 1677622389
transform 1 0 3740 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1677622389
transform 1 0 3740 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1677622389
transform 1 0 3764 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1677622389
transform 1 0 3828 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1677622389
transform 1 0 3788 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5197
timestamp 1677622389
transform 1 0 3836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1677622389
transform 1 0 3772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1677622389
transform 1 0 3788 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4687
timestamp 1677622389
transform 1 0 3788 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1677622389
transform 1 0 3812 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1677622389
transform 1 0 3836 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1677622389
transform 1 0 3884 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5198
timestamp 1677622389
transform 1 0 3884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1677622389
transform 1 0 3908 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4551
timestamp 1677622389
transform 1 0 3924 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1677622389
transform 1 0 3956 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5199
timestamp 1677622389
transform 1 0 3940 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1677622389
transform 1 0 3956 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4659
timestamp 1677622389
transform 1 0 3940 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5292
timestamp 1677622389
transform 1 0 3948 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4690
timestamp 1677622389
transform 1 0 3948 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1677622389
transform 1 0 3972 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5201
timestamp 1677622389
transform 1 0 3972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1677622389
transform 1 0 4012 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4552
timestamp 1677622389
transform 1 0 4076 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1677622389
transform 1 0 4052 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5202
timestamp 1677622389
transform 1 0 4060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1677622389
transform 1 0 4076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1677622389
transform 1 0 4084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1677622389
transform 1 0 4052 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4660
timestamp 1677622389
transform 1 0 4084 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1677622389
transform 1 0 4124 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1677622389
transform 1 0 4164 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1677622389
transform 1 0 4156 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5205
timestamp 1677622389
transform 1 0 4156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1677622389
transform 1 0 4124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1677622389
transform 1 0 4132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1677622389
transform 1 0 4148 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1677622389
transform 1 0 4164 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4691
timestamp 1677622389
transform 1 0 4148 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5206
timestamp 1677622389
transform 1 0 4196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1677622389
transform 1 0 4228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1677622389
transform 1 0 4276 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4692
timestamp 1677622389
transform 1 0 4228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1677622389
transform 1 0 4276 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1677622389
transform 1 0 4292 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5208
timestamp 1677622389
transform 1 0 4292 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4577
timestamp 1677622389
transform 1 0 4332 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5209
timestamp 1677622389
transform 1 0 4340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1677622389
transform 1 0 4388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1677622389
transform 1 0 4404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1677622389
transform 1 0 4420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1677622389
transform 1 0 4372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1677622389
transform 1 0 4380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1677622389
transform 1 0 4396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1677622389
transform 1 0 4412 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4710
timestamp 1677622389
transform 1 0 4380 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1677622389
transform 1 0 4452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1677622389
transform 1 0 4476 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5119
timestamp 1677622389
transform 1 0 4460 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1677622389
transform 1 0 4452 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4636
timestamp 1677622389
transform 1 0 4460 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5213
timestamp 1677622389
transform 1 0 4468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1677622389
transform 1 0 4444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1677622389
transform 1 0 4484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1677622389
transform 1 0 4500 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4553
timestamp 1677622389
transform 1 0 4548 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1677622389
transform 1 0 4540 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5215
timestamp 1677622389
transform 1 0 4532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1677622389
transform 1 0 4548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1677622389
transform 1 0 4556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1677622389
transform 1 0 4580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1677622389
transform 1 0 4524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1677622389
transform 1 0 4540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1677622389
transform 1 0 4548 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4661
timestamp 1677622389
transform 1 0 4556 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5308
timestamp 1677622389
transform 1 0 4572 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4693
timestamp 1677622389
transform 1 0 4524 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1677622389
transform 1 0 4580 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1677622389
transform 1 0 4548 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5309
timestamp 1677622389
transform 1 0 4596 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4637
timestamp 1677622389
transform 1 0 4604 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5310
timestamp 1677622389
transform 1 0 4620 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4712
timestamp 1677622389
transform 1 0 4620 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1677622389
transform 1 0 4652 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5219
timestamp 1677622389
transform 1 0 4636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1677622389
transform 1 0 4652 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4627
timestamp 1677622389
transform 1 0 4764 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1677622389
transform 1 0 4676 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5221
timestamp 1677622389
transform 1 0 4700 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4639
timestamp 1677622389
transform 1 0 4740 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5222
timestamp 1677622389
transform 1 0 4756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1677622389
transform 1 0 4764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1677622389
transform 1 0 4644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1677622389
transform 1 0 4660 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1677622389
transform 1 0 4676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4695
timestamp 1677622389
transform 1 0 4676 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5314
timestamp 1677622389
transform 1 0 4780 0 1 2205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_50
timestamp 1677622389
transform 1 0 48 0 1 2170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_339
timestamp 1677622389
transform 1 0 72 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_390
timestamp 1677622389
transform -1 0 184 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_4713
timestamp 1677622389
transform 1 0 220 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_238
timestamp 1677622389
transform -1 0 224 0 1 2170
box -8 -3 46 105
use M3_M2  M3_M2_4714
timestamp 1677622389
transform 1 0 244 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_340
timestamp 1677622389
transform 1 0 224 0 1 2170
box -8 -3 104 105
use FILL  FILL_5955
timestamp 1677622389
transform 1 0 320 0 1 2170
box -8 -3 16 105
use FILL  FILL_5956
timestamp 1677622389
transform 1 0 328 0 1 2170
box -8 -3 16 105
use FILL  FILL_5957
timestamp 1677622389
transform 1 0 336 0 1 2170
box -8 -3 16 105
use FILL  FILL_5958
timestamp 1677622389
transform 1 0 344 0 1 2170
box -8 -3 16 105
use FILL  FILL_5959
timestamp 1677622389
transform 1 0 352 0 1 2170
box -8 -3 16 105
use FILL  FILL_5970
timestamp 1677622389
transform 1 0 360 0 1 2170
box -8 -3 16 105
use FILL  FILL_5972
timestamp 1677622389
transform 1 0 368 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_61
timestamp 1677622389
transform -1 0 400 0 1 2170
box -5 -3 28 105
use FILL  FILL_5973
timestamp 1677622389
transform 1 0 400 0 1 2170
box -8 -3 16 105
use FILL  FILL_5974
timestamp 1677622389
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_5975
timestamp 1677622389
transform 1 0 416 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4715
timestamp 1677622389
transform 1 0 436 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_393
timestamp 1677622389
transform 1 0 424 0 1 2170
box -9 -3 26 105
use FILL  FILL_5976
timestamp 1677622389
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_5977
timestamp 1677622389
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_5978
timestamp 1677622389
transform 1 0 456 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_227
timestamp 1677622389
transform 1 0 464 0 1 2170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_342
timestamp 1677622389
transform -1 0 600 0 1 2170
box -8 -3 104 105
use FILL  FILL_5979
timestamp 1677622389
transform 1 0 600 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_62
timestamp 1677622389
transform 1 0 608 0 1 2170
box -5 -3 28 105
use FILL  FILL_5980
timestamp 1677622389
transform 1 0 632 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_63
timestamp 1677622389
transform -1 0 664 0 1 2170
box -5 -3 28 105
use FILL  FILL_5981
timestamp 1677622389
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_5997
timestamp 1677622389
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_5999
timestamp 1677622389
transform 1 0 680 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_56
timestamp 1677622389
transform 1 0 688 0 1 2170
box -8 -3 32 105
use FILL  FILL_6001
timestamp 1677622389
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6002
timestamp 1677622389
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6003
timestamp 1677622389
transform 1 0 728 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_243
timestamp 1677622389
transform 1 0 736 0 1 2170
box -8 -3 46 105
use FILL  FILL_6004
timestamp 1677622389
transform 1 0 776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6005
timestamp 1677622389
transform 1 0 784 0 1 2170
box -8 -3 16 105
use FILL  FILL_6007
timestamp 1677622389
transform 1 0 792 0 1 2170
box -8 -3 16 105
use FILL  FILL_6009
timestamp 1677622389
transform 1 0 800 0 1 2170
box -8 -3 16 105
use FILL  FILL_6011
timestamp 1677622389
transform 1 0 808 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4716
timestamp 1677622389
transform 1 0 884 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_344
timestamp 1677622389
transform 1 0 816 0 1 2170
box -8 -3 104 105
use FILL  FILL_6013
timestamp 1677622389
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_6025
timestamp 1677622389
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_6027
timestamp 1677622389
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_6029
timestamp 1677622389
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_6031
timestamp 1677622389
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_6033
timestamp 1677622389
transform 1 0 952 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_244
timestamp 1677622389
transform 1 0 960 0 1 2170
box -8 -3 46 105
use FILL  FILL_6035
timestamp 1677622389
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6037
timestamp 1677622389
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6039
timestamp 1677622389
transform 1 0 1016 0 1 2170
box -8 -3 16 105
use FILL  FILL_6041
timestamp 1677622389
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6043
timestamp 1677622389
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_57
timestamp 1677622389
transform 1 0 1040 0 1 2170
box -8 -3 32 105
use FILL  FILL_6045
timestamp 1677622389
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_6050
timestamp 1677622389
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_6052
timestamp 1677622389
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_6054
timestamp 1677622389
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6056
timestamp 1677622389
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6058
timestamp 1677622389
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6060
timestamp 1677622389
transform 1 0 1112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6061
timestamp 1677622389
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6062
timestamp 1677622389
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6063
timestamp 1677622389
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_115
timestamp 1677622389
transform 1 0 1144 0 1 2170
box -8 -3 34 105
use FILL  FILL_6064
timestamp 1677622389
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6070
timestamp 1677622389
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_6072
timestamp 1677622389
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6074
timestamp 1677622389
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6076
timestamp 1677622389
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6078
timestamp 1677622389
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6080
timestamp 1677622389
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6082
timestamp 1677622389
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6084
timestamp 1677622389
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_6086
timestamp 1677622389
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_117
timestamp 1677622389
transform -1 0 1288 0 1 2170
box -8 -3 34 105
use FILL  FILL_6087
timestamp 1677622389
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6094
timestamp 1677622389
transform 1 0 1296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6096
timestamp 1677622389
transform 1 0 1304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6098
timestamp 1677622389
transform 1 0 1312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6100
timestamp 1677622389
transform 1 0 1320 0 1 2170
box -8 -3 16 105
use FILL  FILL_6102
timestamp 1677622389
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_6104
timestamp 1677622389
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_345
timestamp 1677622389
transform -1 0 1440 0 1 2170
box -8 -3 104 105
use FILL  FILL_6105
timestamp 1677622389
transform 1 0 1440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6116
timestamp 1677622389
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6118
timestamp 1677622389
transform 1 0 1456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6120
timestamp 1677622389
transform 1 0 1464 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_229
timestamp 1677622389
transform -1 0 1512 0 1 2170
box -8 -3 46 105
use FILL  FILL_6121
timestamp 1677622389
transform 1 0 1512 0 1 2170
box -8 -3 16 105
use FILL  FILL_6124
timestamp 1677622389
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6126
timestamp 1677622389
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6128
timestamp 1677622389
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6129
timestamp 1677622389
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_346
timestamp 1677622389
transform -1 0 1648 0 1 2170
box -8 -3 104 105
use FILL  FILL_6130
timestamp 1677622389
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_6131
timestamp 1677622389
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_6132
timestamp 1677622389
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_6133
timestamp 1677622389
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_6144
timestamp 1677622389
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_6146
timestamp 1677622389
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_231
timestamp 1677622389
transform -1 0 1736 0 1 2170
box -8 -3 46 105
use FILL  FILL_6147
timestamp 1677622389
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use FILL  FILL_6152
timestamp 1677622389
transform 1 0 1744 0 1 2170
box -8 -3 16 105
use FILL  FILL_6153
timestamp 1677622389
transform 1 0 1752 0 1 2170
box -8 -3 16 105
use FILL  FILL_6154
timestamp 1677622389
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_6155
timestamp 1677622389
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_6156
timestamp 1677622389
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6157
timestamp 1677622389
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use FILL  FILL_6158
timestamp 1677622389
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_6159
timestamp 1677622389
transform 1 0 1800 0 1 2170
box -8 -3 16 105
use FILL  FILL_6160
timestamp 1677622389
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_6161
timestamp 1677622389
transform 1 0 1816 0 1 2170
box -8 -3 16 105
use FILL  FILL_6162
timestamp 1677622389
transform 1 0 1824 0 1 2170
box -8 -3 16 105
use FILL  FILL_6163
timestamp 1677622389
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_6164
timestamp 1677622389
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_6165
timestamp 1677622389
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6166
timestamp 1677622389
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6167
timestamp 1677622389
transform 1 0 1864 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4717
timestamp 1677622389
transform 1 0 1884 0 1 2175
box -3 -3 3 3
use FILL  FILL_6168
timestamp 1677622389
transform 1 0 1872 0 1 2170
box -8 -3 16 105
use FILL  FILL_6171
timestamp 1677622389
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_6173
timestamp 1677622389
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6175
timestamp 1677622389
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_6177
timestamp 1677622389
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6179
timestamp 1677622389
transform 1 0 1912 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_232
timestamp 1677622389
transform -1 0 1960 0 1 2170
box -8 -3 46 105
use FILL  FILL_6180
timestamp 1677622389
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_6188
timestamp 1677622389
transform 1 0 1968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6190
timestamp 1677622389
transform 1 0 1976 0 1 2170
box -8 -3 16 105
use FILL  FILL_6192
timestamp 1677622389
transform 1 0 1984 0 1 2170
box -8 -3 16 105
use FILL  FILL_6194
timestamp 1677622389
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_6196
timestamp 1677622389
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6198
timestamp 1677622389
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6200
timestamp 1677622389
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_398
timestamp 1677622389
transform -1 0 2040 0 1 2170
box -9 -3 26 105
use FILL  FILL_6201
timestamp 1677622389
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_6202
timestamp 1677622389
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_6203
timestamp 1677622389
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_6204
timestamp 1677622389
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_6205
timestamp 1677622389
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4718
timestamp 1677622389
transform 1 0 2092 0 1 2175
box -3 -3 3 3
use FILL  FILL_6209
timestamp 1677622389
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_348
timestamp 1677622389
transform -1 0 2184 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_349
timestamp 1677622389
transform -1 0 2280 0 1 2170
box -8 -3 104 105
use FILL  FILL_6210
timestamp 1677622389
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_6211
timestamp 1677622389
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6229
timestamp 1677622389
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6231
timestamp 1677622389
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6233
timestamp 1677622389
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6235
timestamp 1677622389
transform 1 0 2320 0 1 2170
box -8 -3 16 105
use FILL  FILL_6237
timestamp 1677622389
transform 1 0 2328 0 1 2170
box -8 -3 16 105
use FILL  FILL_6239
timestamp 1677622389
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_6240
timestamp 1677622389
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_6241
timestamp 1677622389
transform 1 0 2352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6242
timestamp 1677622389
transform 1 0 2360 0 1 2170
box -8 -3 16 105
use FILL  FILL_6243
timestamp 1677622389
transform 1 0 2368 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_247
timestamp 1677622389
transform -1 0 2416 0 1 2170
box -8 -3 46 105
use FILL  FILL_6244
timestamp 1677622389
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use FILL  FILL_6252
timestamp 1677622389
transform 1 0 2424 0 1 2170
box -8 -3 16 105
use FILL  FILL_6253
timestamp 1677622389
transform 1 0 2432 0 1 2170
box -8 -3 16 105
use FILL  FILL_6254
timestamp 1677622389
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_350
timestamp 1677622389
transform -1 0 2544 0 1 2170
box -8 -3 104 105
use FILL  FILL_6255
timestamp 1677622389
transform 1 0 2544 0 1 2170
box -8 -3 16 105
use FILL  FILL_6256
timestamp 1677622389
transform 1 0 2552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6265
timestamp 1677622389
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use FILL  FILL_6267
timestamp 1677622389
transform 1 0 2568 0 1 2170
box -8 -3 16 105
use FILL  FILL_6269
timestamp 1677622389
transform 1 0 2576 0 1 2170
box -8 -3 16 105
use FILL  FILL_6271
timestamp 1677622389
transform 1 0 2584 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_248
timestamp 1677622389
transform 1 0 2592 0 1 2170
box -8 -3 46 105
use FILL  FILL_6273
timestamp 1677622389
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use FILL  FILL_6274
timestamp 1677622389
transform 1 0 2640 0 1 2170
box -8 -3 16 105
use FILL  FILL_6275
timestamp 1677622389
transform 1 0 2648 0 1 2170
box -8 -3 16 105
use FILL  FILL_6279
timestamp 1677622389
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use FILL  FILL_6281
timestamp 1677622389
transform 1 0 2664 0 1 2170
box -8 -3 16 105
use FILL  FILL_6283
timestamp 1677622389
transform 1 0 2672 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_399
timestamp 1677622389
transform 1 0 2680 0 1 2170
box -9 -3 26 105
use FILL  FILL_6285
timestamp 1677622389
transform 1 0 2696 0 1 2170
box -8 -3 16 105
use FILL  FILL_6286
timestamp 1677622389
transform 1 0 2704 0 1 2170
box -8 -3 16 105
use FILL  FILL_6289
timestamp 1677622389
transform 1 0 2712 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_351
timestamp 1677622389
transform 1 0 2720 0 1 2170
box -8 -3 104 105
use FILL  FILL_6291
timestamp 1677622389
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_58
timestamp 1677622389
transform 1 0 2824 0 1 2170
box -8 -3 32 105
use FILL  FILL_6292
timestamp 1677622389
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6303
timestamp 1677622389
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6305
timestamp 1677622389
transform 1 0 2864 0 1 2170
box -8 -3 16 105
use FILL  FILL_6307
timestamp 1677622389
transform 1 0 2872 0 1 2170
box -8 -3 16 105
use FILL  FILL_6309
timestamp 1677622389
transform 1 0 2880 0 1 2170
box -8 -3 16 105
use FILL  FILL_6310
timestamp 1677622389
transform 1 0 2888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6311
timestamp 1677622389
transform 1 0 2896 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_120
timestamp 1677622389
transform -1 0 2936 0 1 2170
box -8 -3 34 105
use FILL  FILL_6312
timestamp 1677622389
transform 1 0 2936 0 1 2170
box -8 -3 16 105
use FILL  FILL_6317
timestamp 1677622389
transform 1 0 2944 0 1 2170
box -8 -3 16 105
use FILL  FILL_6319
timestamp 1677622389
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use FILL  FILL_6321
timestamp 1677622389
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_6322
timestamp 1677622389
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6323
timestamp 1677622389
transform 1 0 2976 0 1 2170
box -8 -3 16 105
use FILL  FILL_6324
timestamp 1677622389
transform 1 0 2984 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_352
timestamp 1677622389
transform 1 0 2992 0 1 2170
box -8 -3 104 105
use FILL  FILL_6325
timestamp 1677622389
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6334
timestamp 1677622389
transform 1 0 3096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6336
timestamp 1677622389
transform 1 0 3104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6338
timestamp 1677622389
transform 1 0 3112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6339
timestamp 1677622389
transform 1 0 3120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6340
timestamp 1677622389
transform 1 0 3128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6341
timestamp 1677622389
transform 1 0 3136 0 1 2170
box -8 -3 16 105
use FILL  FILL_6342
timestamp 1677622389
transform 1 0 3144 0 1 2170
box -8 -3 16 105
use FILL  FILL_6343
timestamp 1677622389
transform 1 0 3152 0 1 2170
box -8 -3 16 105
use FILL  FILL_6344
timestamp 1677622389
transform 1 0 3160 0 1 2170
box -8 -3 16 105
use FILL  FILL_6347
timestamp 1677622389
transform 1 0 3168 0 1 2170
box -8 -3 16 105
use FILL  FILL_6349
timestamp 1677622389
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_68
timestamp 1677622389
transform -1 0 3208 0 1 2170
box -5 -3 28 105
use FILL  FILL_6350
timestamp 1677622389
transform 1 0 3208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6351
timestamp 1677622389
transform 1 0 3216 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_69
timestamp 1677622389
transform 1 0 3224 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_70
timestamp 1677622389
transform 1 0 3248 0 1 2170
box -5 -3 28 105
use FILL  FILL_6352
timestamp 1677622389
transform 1 0 3272 0 1 2170
box -8 -3 16 105
use FILL  FILL_6353
timestamp 1677622389
transform 1 0 3280 0 1 2170
box -8 -3 16 105
use FILL  FILL_6354
timestamp 1677622389
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6358
timestamp 1677622389
transform 1 0 3296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6359
timestamp 1677622389
transform 1 0 3304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6360
timestamp 1677622389
transform 1 0 3312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6362
timestamp 1677622389
transform 1 0 3320 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_250
timestamp 1677622389
transform 1 0 3328 0 1 2170
box -8 -3 46 105
use FILL  FILL_6364
timestamp 1677622389
transform 1 0 3368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6365
timestamp 1677622389
transform 1 0 3376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6366
timestamp 1677622389
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6367
timestamp 1677622389
transform 1 0 3392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6368
timestamp 1677622389
transform 1 0 3400 0 1 2170
box -8 -3 16 105
use AND2X2  AND2X2_19
timestamp 1677622389
transform 1 0 3408 0 1 2170
box -8 -3 40 105
use FILL  FILL_6375
timestamp 1677622389
transform 1 0 3440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6381
timestamp 1677622389
transform 1 0 3448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6383
timestamp 1677622389
transform 1 0 3456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6385
timestamp 1677622389
transform 1 0 3464 0 1 2170
box -8 -3 16 105
use FILL  FILL_6387
timestamp 1677622389
transform 1 0 3472 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_251
timestamp 1677622389
transform 1 0 3480 0 1 2170
box -8 -3 46 105
use FILL  FILL_6389
timestamp 1677622389
transform 1 0 3520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6392
timestamp 1677622389
transform 1 0 3528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6394
timestamp 1677622389
transform 1 0 3536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6396
timestamp 1677622389
transform 1 0 3544 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4719
timestamp 1677622389
transform 1 0 3564 0 1 2175
box -3 -3 3 3
use FILL  FILL_6398
timestamp 1677622389
transform 1 0 3552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6400
timestamp 1677622389
transform 1 0 3560 0 1 2170
box -8 -3 16 105
use FILL  FILL_6401
timestamp 1677622389
transform 1 0 3568 0 1 2170
box -8 -3 16 105
use FILL  FILL_6402
timestamp 1677622389
transform 1 0 3576 0 1 2170
box -8 -3 16 105
use FILL  FILL_6403
timestamp 1677622389
transform 1 0 3584 0 1 2170
box -8 -3 16 105
use FILL  FILL_6404
timestamp 1677622389
transform 1 0 3592 0 1 2170
box -8 -3 16 105
use FILL  FILL_6405
timestamp 1677622389
transform 1 0 3600 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_403
timestamp 1677622389
transform -1 0 3624 0 1 2170
box -9 -3 26 105
use FILL  FILL_6406
timestamp 1677622389
transform 1 0 3624 0 1 2170
box -8 -3 16 105
use FILL  FILL_6411
timestamp 1677622389
transform 1 0 3632 0 1 2170
box -8 -3 16 105
use FILL  FILL_6413
timestamp 1677622389
transform 1 0 3640 0 1 2170
box -8 -3 16 105
use FILL  FILL_6415
timestamp 1677622389
transform 1 0 3648 0 1 2170
box -8 -3 16 105
use FILL  FILL_6416
timestamp 1677622389
transform 1 0 3656 0 1 2170
box -8 -3 16 105
use FILL  FILL_6417
timestamp 1677622389
transform 1 0 3664 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4720
timestamp 1677622389
transform 1 0 3708 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_238
timestamp 1677622389
transform 1 0 3672 0 1 2170
box -8 -3 46 105
use FILL  FILL_6418
timestamp 1677622389
transform 1 0 3712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6419
timestamp 1677622389
transform 1 0 3720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6420
timestamp 1677622389
transform 1 0 3728 0 1 2170
box -8 -3 16 105
use FILL  FILL_6421
timestamp 1677622389
transform 1 0 3736 0 1 2170
box -8 -3 16 105
use FILL  FILL_6422
timestamp 1677622389
transform 1 0 3744 0 1 2170
box -8 -3 16 105
use FILL  FILL_6423
timestamp 1677622389
transform 1 0 3752 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_404
timestamp 1677622389
transform -1 0 3776 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_354
timestamp 1677622389
transform 1 0 3776 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_405
timestamp 1677622389
transform 1 0 3872 0 1 2170
box -9 -3 26 105
use FILL  FILL_6435
timestamp 1677622389
transform 1 0 3888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6437
timestamp 1677622389
transform 1 0 3896 0 1 2170
box -8 -3 16 105
use FILL  FILL_6439
timestamp 1677622389
transform 1 0 3904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6441
timestamp 1677622389
transform 1 0 3912 0 1 2170
box -8 -3 16 105
use FILL  FILL_6443
timestamp 1677622389
transform 1 0 3920 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_240
timestamp 1677622389
transform 1 0 3928 0 1 2170
box -8 -3 46 105
use FILL  FILL_6444
timestamp 1677622389
transform 1 0 3968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6447
timestamp 1677622389
transform 1 0 3976 0 1 2170
box -8 -3 16 105
use FILL  FILL_6449
timestamp 1677622389
transform 1 0 3984 0 1 2170
box -8 -3 16 105
use FILL  FILL_6450
timestamp 1677622389
transform 1 0 3992 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4721
timestamp 1677622389
transform 1 0 4012 0 1 2175
box -3 -3 3 3
use FILL  FILL_6451
timestamp 1677622389
transform 1 0 4000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6452
timestamp 1677622389
transform 1 0 4008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6453
timestamp 1677622389
transform 1 0 4016 0 1 2170
box -8 -3 16 105
use FILL  FILL_6454
timestamp 1677622389
transform 1 0 4024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6455
timestamp 1677622389
transform 1 0 4032 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_252
timestamp 1677622389
transform 1 0 4040 0 1 2170
box -8 -3 46 105
use FILL  FILL_6456
timestamp 1677622389
transform 1 0 4080 0 1 2170
box -8 -3 16 105
use FILL  FILL_6457
timestamp 1677622389
transform 1 0 4088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6458
timestamp 1677622389
transform 1 0 4096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6460
timestamp 1677622389
transform 1 0 4104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6462
timestamp 1677622389
transform 1 0 4112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6463
timestamp 1677622389
transform 1 0 4120 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4722
timestamp 1677622389
transform 1 0 4164 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_242
timestamp 1677622389
transform 1 0 4128 0 1 2170
box -8 -3 46 105
use FILL  FILL_6464
timestamp 1677622389
transform 1 0 4168 0 1 2170
box -8 -3 16 105
use FILL  FILL_6465
timestamp 1677622389
transform 1 0 4176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6466
timestamp 1677622389
transform 1 0 4184 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4723
timestamp 1677622389
transform 1 0 4236 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_357
timestamp 1677622389
transform -1 0 4288 0 1 2170
box -8 -3 104 105
use FILL  FILL_6467
timestamp 1677622389
transform 1 0 4288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6477
timestamp 1677622389
transform 1 0 4296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6478
timestamp 1677622389
transform 1 0 4304 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_410
timestamp 1677622389
transform -1 0 4328 0 1 2170
box -9 -3 26 105
use FILL  FILL_6479
timestamp 1677622389
transform 1 0 4328 0 1 2170
box -8 -3 16 105
use FILL  FILL_6480
timestamp 1677622389
transform 1 0 4336 0 1 2170
box -8 -3 16 105
use FILL  FILL_6481
timestamp 1677622389
transform 1 0 4344 0 1 2170
box -8 -3 16 105
use FILL  FILL_6482
timestamp 1677622389
transform 1 0 4352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6483
timestamp 1677622389
transform 1 0 4360 0 1 2170
box -8 -3 16 105
use FILL  FILL_6484
timestamp 1677622389
transform 1 0 4368 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4724
timestamp 1677622389
transform 1 0 4388 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_245
timestamp 1677622389
transform 1 0 4376 0 1 2170
box -8 -3 46 105
use FILL  FILL_6485
timestamp 1677622389
transform 1 0 4416 0 1 2170
box -8 -3 16 105
use FILL  FILL_6490
timestamp 1677622389
transform 1 0 4424 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_411
timestamp 1677622389
transform -1 0 4448 0 1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_40
timestamp 1677622389
transform -1 0 4480 0 1 2170
box -8 -3 40 105
use FILL  FILL_6491
timestamp 1677622389
transform 1 0 4480 0 1 2170
box -8 -3 16 105
use FILL  FILL_6492
timestamp 1677622389
transform 1 0 4488 0 1 2170
box -8 -3 16 105
use FILL  FILL_6493
timestamp 1677622389
transform 1 0 4496 0 1 2170
box -8 -3 16 105
use FILL  FILL_6494
timestamp 1677622389
transform 1 0 4504 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_253
timestamp 1677622389
transform 1 0 4512 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_246
timestamp 1677622389
transform 1 0 4552 0 1 2170
box -8 -3 46 105
use FILL  FILL_6495
timestamp 1677622389
transform 1 0 4592 0 1 2170
box -8 -3 16 105
use FILL  FILL_6496
timestamp 1677622389
transform 1 0 4600 0 1 2170
box -8 -3 16 105
use FILL  FILL_6497
timestamp 1677622389
transform 1 0 4608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6498
timestamp 1677622389
transform 1 0 4616 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_247
timestamp 1677622389
transform 1 0 4624 0 1 2170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_359
timestamp 1677622389
transform 1 0 4664 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_412
timestamp 1677622389
transform -1 0 4776 0 1 2170
box -9 -3 26 105
use FILL  FILL_6499
timestamp 1677622389
transform 1 0 4776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6500
timestamp 1677622389
transform 1 0 4784 0 1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_51
timestamp 1677622389
transform 1 0 4819 0 1 2170
box -10 -3 10 3
use M2_M1  M2_M1_5322
timestamp 1677622389
transform 1 0 92 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4787
timestamp 1677622389
transform 1 0 172 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5407
timestamp 1677622389
transform 1 0 140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1677622389
transform 1 0 172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1677622389
transform 1 0 180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4833
timestamp 1677622389
transform 1 0 140 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1677622389
transform 1 0 180 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5323
timestamp 1677622389
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4758
timestamp 1677622389
transform 1 0 212 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5324
timestamp 1677622389
transform 1 0 212 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4788
timestamp 1677622389
transform 1 0 220 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5325
timestamp 1677622389
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1677622389
transform 1 0 204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1677622389
transform 1 0 220 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4835
timestamp 1677622389
transform 1 0 196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1677622389
transform 1 0 228 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5412
timestamp 1677622389
transform 1 0 236 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4836
timestamp 1677622389
transform 1 0 220 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1677622389
transform 1 0 236 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1677622389
transform 1 0 204 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5413
timestamp 1677622389
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1677622389
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4838
timestamp 1677622389
transform 1 0 284 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1677622389
transform 1 0 340 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5326
timestamp 1677622389
transform 1 0 316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1677622389
transform 1 0 324 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4789
timestamp 1677622389
transform 1 0 332 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5328
timestamp 1677622389
transform 1 0 340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1677622389
transform 1 0 332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1677622389
transform 1 0 380 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4854
timestamp 1677622389
transform 1 0 380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1677622389
transform 1 0 396 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5329
timestamp 1677622389
transform 1 0 396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1677622389
transform 1 0 404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1677622389
transform 1 0 428 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4743
timestamp 1677622389
transform 1 0 444 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1677622389
transform 1 0 460 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1677622389
transform 1 0 436 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5330
timestamp 1677622389
transform 1 0 436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1677622389
transform 1 0 444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1677622389
transform 1 0 460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1677622389
transform 1 0 452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1677622389
transform 1 0 460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1677622389
transform 1 0 476 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4839
timestamp 1677622389
transform 1 0 444 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1677622389
transform 1 0 476 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1677622389
transform 1 0 460 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1677622389
transform 1 0 508 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1677622389
transform 1 0 524 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1677622389
transform 1 0 540 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1677622389
transform 1 0 556 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1677622389
transform 1 0 564 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5333
timestamp 1677622389
transform 1 0 532 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1677622389
transform 1 0 516 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4791
timestamp 1677622389
transform 1 0 540 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1677622389
transform 1 0 580 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5334
timestamp 1677622389
transform 1 0 548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1677622389
transform 1 0 564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1677622389
transform 1 0 524 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4819
timestamp 1677622389
transform 1 0 532 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5424
timestamp 1677622389
transform 1 0 540 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4820
timestamp 1677622389
transform 1 0 548 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5425
timestamp 1677622389
transform 1 0 556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4792
timestamp 1677622389
transform 1 0 572 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5426
timestamp 1677622389
transform 1 0 572 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4793
timestamp 1677622389
transform 1 0 612 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5427
timestamp 1677622389
transform 1 0 628 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4855
timestamp 1677622389
transform 1 0 612 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1677622389
transform 1 0 628 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1677622389
transform 1 0 620 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1677622389
transform 1 0 660 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5336
timestamp 1677622389
transform 1 0 644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1677622389
transform 1 0 652 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4725
timestamp 1677622389
transform 1 0 676 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5428
timestamp 1677622389
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4841
timestamp 1677622389
transform 1 0 668 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1677622389
transform 1 0 716 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1677622389
transform 1 0 748 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1677622389
transform 1 0 740 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1677622389
transform 1 0 700 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1677622389
transform 1 0 740 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5338
timestamp 1677622389
transform 1 0 700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1677622389
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1677622389
transform 1 0 780 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4842
timestamp 1677622389
transform 1 0 724 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1677622389
transform 1 0 756 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1677622389
transform 1 0 828 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5431
timestamp 1677622389
transform 1 0 852 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4821
timestamp 1677622389
transform 1 0 860 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5432
timestamp 1677622389
transform 1 0 900 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4843
timestamp 1677622389
transform 1 0 900 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1677622389
transform 1 0 972 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1677622389
transform 1 0 964 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1677622389
transform 1 0 964 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1677622389
transform 1 0 980 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5339
timestamp 1677622389
transform 1 0 964 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1677622389
transform 1 0 972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1677622389
transform 1 0 980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1677622389
transform 1 0 996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1677622389
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1677622389
transform 1 0 1060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1677622389
transform 1 0 1084 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4822
timestamp 1677622389
transform 1 0 1084 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1677622389
transform 1 0 1124 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5436
timestamp 1677622389
transform 1 0 1124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1677622389
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4769
timestamp 1677622389
transform 1 0 1156 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1677622389
transform 1 0 1156 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1677622389
transform 1 0 1220 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5438
timestamp 1677622389
transform 1 0 1252 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4845
timestamp 1677622389
transform 1 0 1252 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1677622389
transform 1 0 1308 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5510
timestamp 1677622389
transform 1 0 1308 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1677622389
transform 1 0 1348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1677622389
transform 1 0 1340 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4795
timestamp 1677622389
transform 1 0 1388 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5439
timestamp 1677622389
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4729
timestamp 1677622389
transform 1 0 1460 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5319
timestamp 1677622389
transform 1 0 1444 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_4770
timestamp 1677622389
transform 1 0 1452 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5344
timestamp 1677622389
transform 1 0 1452 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4751
timestamp 1677622389
transform 1 0 1468 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5440
timestamp 1677622389
transform 1 0 1460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1677622389
transform 1 0 1484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1677622389
transform 1 0 1492 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4846
timestamp 1677622389
transform 1 0 1492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1677622389
transform 1 0 1516 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1677622389
transform 1 0 1516 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1677622389
transform 1 0 1508 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5346
timestamp 1677622389
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1677622389
transform 1 0 1508 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4847
timestamp 1677622389
transform 1 0 1508 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1677622389
transform 1 0 1508 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5347
timestamp 1677622389
transform 1 0 1556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1677622389
transform 1 0 1612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1677622389
transform 1 0 1644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1677622389
transform 1 0 1652 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4883
timestamp 1677622389
transform 1 0 1652 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5349
timestamp 1677622389
transform 1 0 1668 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4753
timestamp 1677622389
transform 1 0 1692 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5445
timestamp 1677622389
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4884
timestamp 1677622389
transform 1 0 1684 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1677622389
transform 1 0 1708 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1677622389
transform 1 0 1716 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5350
timestamp 1677622389
transform 1 0 1740 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4731
timestamp 1677622389
transform 1 0 1764 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1677622389
transform 1 0 1780 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1677622389
transform 1 0 1788 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5351
timestamp 1677622389
transform 1 0 1836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1677622389
transform 1 0 1756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1677622389
transform 1 0 1788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1677622389
transform 1 0 1852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1677622389
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4799
timestamp 1677622389
transform 1 0 1876 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1677622389
transform 1 0 1868 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1677622389
transform 1 0 1892 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1677622389
transform 1 0 1916 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5353
timestamp 1677622389
transform 1 0 1964 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1677622389
transform 1 0 1972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1677622389
transform 1 0 2060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1677622389
transform 1 0 2052 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1677622389
transform 1 0 2068 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4772
timestamp 1677622389
transform 1 0 2084 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1677622389
transform 1 0 2076 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1677622389
transform 1 0 2172 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5355
timestamp 1677622389
transform 1 0 2156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1677622389
transform 1 0 2172 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1677622389
transform 1 0 2148 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4859
timestamp 1677622389
transform 1 0 2148 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1677622389
transform 1 0 2180 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5357
timestamp 1677622389
transform 1 0 2188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1677622389
transform 1 0 2180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1677622389
transform 1 0 2228 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4801
timestamp 1677622389
transform 1 0 2236 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1677622389
transform 1 0 2260 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5359
timestamp 1677622389
transform 1 0 2268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1677622389
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1677622389
transform 1 0 2276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1677622389
transform 1 0 2284 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4860
timestamp 1677622389
transform 1 0 2276 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1677622389
transform 1 0 2276 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5457
timestamp 1677622389
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1677622389
transform 1 0 2372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1677622389
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1677622389
transform 1 0 2364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1677622389
transform 1 0 2404 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4733
timestamp 1677622389
transform 1 0 2436 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5361
timestamp 1677622389
transform 1 0 2444 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4803
timestamp 1677622389
transform 1 0 2452 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5362
timestamp 1677622389
transform 1 0 2460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1677622389
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1677622389
transform 1 0 2452 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4886
timestamp 1677622389
transform 1 0 2436 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1677622389
transform 1 0 2508 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5363
timestamp 1677622389
transform 1 0 2524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1677622389
transform 1 0 2532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1677622389
transform 1 0 2548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1677622389
transform 1 0 2556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4849
timestamp 1677622389
transform 1 0 2556 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5364
timestamp 1677622389
transform 1 0 2572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1677622389
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1677622389
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1677622389
transform 1 0 2644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1677622389
transform 1 0 2628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1677622389
transform 1 0 2660 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4734
timestamp 1677622389
transform 1 0 2708 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5320
timestamp 1677622389
transform 1 0 2708 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_4735
timestamp 1677622389
transform 1 0 2724 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1677622389
transform 1 0 2724 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5468
timestamp 1677622389
transform 1 0 2748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1677622389
transform 1 0 2780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1677622389
transform 1 0 2788 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4773
timestamp 1677622389
transform 1 0 2804 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5469
timestamp 1677622389
transform 1 0 2796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1677622389
transform 1 0 2804 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1677622389
transform 1 0 2884 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4850
timestamp 1677622389
transform 1 0 2884 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1677622389
transform 1 0 2908 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1677622389
transform 1 0 2924 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5321
timestamp 1677622389
transform 1 0 2924 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1677622389
transform 1 0 2916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1677622389
transform 1 0 2908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1677622389
transform 1 0 2892 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1677622389
transform 1 0 2932 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4774
timestamp 1677622389
transform 1 0 2996 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5372
timestamp 1677622389
transform 1 0 2972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1677622389
transform 1 0 2980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1677622389
transform 1 0 2980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1677622389
transform 1 0 2996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1677622389
transform 1 0 3012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1677622389
transform 1 0 3020 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4851
timestamp 1677622389
transform 1 0 2980 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1677622389
transform 1 0 2972 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1677622389
transform 1 0 3076 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5374
timestamp 1677622389
transform 1 0 3084 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4775
timestamp 1677622389
transform 1 0 3100 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5375
timestamp 1677622389
transform 1 0 3116 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4776
timestamp 1677622389
transform 1 0 3140 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1677622389
transform 1 0 3132 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5376
timestamp 1677622389
transform 1 0 3140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1677622389
transform 1 0 3156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1677622389
transform 1 0 3132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1677622389
transform 1 0 3148 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4824
timestamp 1677622389
transform 1 0 3156 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1677622389
transform 1 0 3228 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5378
timestamp 1677622389
transform 1 0 3204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1677622389
transform 1 0 3228 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4808
timestamp 1677622389
transform 1 0 3308 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5480
timestamp 1677622389
transform 1 0 3308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1677622389
transform 1 0 3332 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1677622389
transform 1 0 3356 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4736
timestamp 1677622389
transform 1 0 3380 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1677622389
transform 1 0 3388 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5380
timestamp 1677622389
transform 1 0 3372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1677622389
transform 1 0 3364 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4861
timestamp 1677622389
transform 1 0 3364 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5481
timestamp 1677622389
transform 1 0 3380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1677622389
transform 1 0 3404 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4862
timestamp 1677622389
transform 1 0 3404 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1677622389
transform 1 0 3436 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1677622389
transform 1 0 3452 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5482
timestamp 1677622389
transform 1 0 3484 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4863
timestamp 1677622389
transform 1 0 3484 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1677622389
transform 1 0 3508 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1677622389
transform 1 0 3500 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5483
timestamp 1677622389
transform 1 0 3508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1677622389
transform 1 0 3500 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4888
timestamp 1677622389
transform 1 0 3500 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5381
timestamp 1677622389
transform 1 0 3524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1677622389
transform 1 0 3564 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4880
timestamp 1677622389
transform 1 0 3564 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1677622389
transform 1 0 3588 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5382
timestamp 1677622389
transform 1 0 3588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1677622389
transform 1 0 3604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1677622389
transform 1 0 3580 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4827
timestamp 1677622389
transform 1 0 3604 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1677622389
transform 1 0 3604 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5384
timestamp 1677622389
transform 1 0 3644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1677622389
transform 1 0 3628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1677622389
transform 1 0 3636 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4779
timestamp 1677622389
transform 1 0 3692 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5385
timestamp 1677622389
transform 1 0 3740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1677622389
transform 1 0 3692 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4865
timestamp 1677622389
transform 1 0 3700 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5386
timestamp 1677622389
transform 1 0 3764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1677622389
transform 1 0 3764 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4866
timestamp 1677622389
transform 1 0 3764 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5387
timestamp 1677622389
transform 1 0 3812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1677622389
transform 1 0 3820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1677622389
transform 1 0 3836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1677622389
transform 1 0 3844 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4828
timestamp 1677622389
transform 1 0 3844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1677622389
transform 1 0 3860 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5389
timestamp 1677622389
transform 1 0 3860 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4809
timestamp 1677622389
transform 1 0 3892 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5491
timestamp 1677622389
transform 1 0 3892 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4867
timestamp 1677622389
transform 1 0 3892 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5390
timestamp 1677622389
transform 1 0 3908 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4780
timestamp 1677622389
transform 1 0 3940 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5391
timestamp 1677622389
transform 1 0 3940 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4810
timestamp 1677622389
transform 1 0 3948 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5392
timestamp 1677622389
transform 1 0 3956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1677622389
transform 1 0 3932 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4829
timestamp 1677622389
transform 1 0 3940 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5493
timestamp 1677622389
transform 1 0 3948 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4868
timestamp 1677622389
transform 1 0 3948 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1677622389
transform 1 0 4060 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1677622389
transform 1 0 4020 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5393
timestamp 1677622389
transform 1 0 3996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1677622389
transform 1 0 4020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1677622389
transform 1 0 4092 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4869
timestamp 1677622389
transform 1 0 4092 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1677622389
transform 1 0 4084 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5394
timestamp 1677622389
transform 1 0 4108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1677622389
transform 1 0 4116 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4870
timestamp 1677622389
transform 1 0 4116 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1677622389
transform 1 0 4132 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5396
timestamp 1677622389
transform 1 0 4140 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4811
timestamp 1677622389
transform 1 0 4148 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5496
timestamp 1677622389
transform 1 0 4132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1677622389
transform 1 0 4148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1677622389
transform 1 0 4164 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4740
timestamp 1677622389
transform 1 0 4172 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5397
timestamp 1677622389
transform 1 0 4172 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4812
timestamp 1677622389
transform 1 0 4180 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1677622389
transform 1 0 4172 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5398
timestamp 1677622389
transform 1 0 4196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1677622389
transform 1 0 4188 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4871
timestamp 1677622389
transform 1 0 4188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1677622389
transform 1 0 4228 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5399
timestamp 1677622389
transform 1 0 4244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1677622389
transform 1 0 4252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1677622389
transform 1 0 4268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1677622389
transform 1 0 4236 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4813
timestamp 1677622389
transform 1 0 4276 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5501
timestamp 1677622389
transform 1 0 4276 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4853
timestamp 1677622389
transform 1 0 4252 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1677622389
transform 1 0 4276 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1677622389
transform 1 0 4292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1677622389
transform 1 0 4324 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5402
timestamp 1677622389
transform 1 0 4292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1677622389
transform 1 0 4308 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4814
timestamp 1677622389
transform 1 0 4396 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5502
timestamp 1677622389
transform 1 0 4332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1677622389
transform 1 0 4388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4784
timestamp 1677622389
transform 1 0 4412 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1677622389
transform 1 0 4468 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5404
timestamp 1677622389
transform 1 0 4516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1677622389
transform 1 0 4436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1677622389
transform 1 0 4468 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4741
timestamp 1677622389
transform 1 0 4596 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1677622389
transform 1 0 4572 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1677622389
transform 1 0 4596 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5405
timestamp 1677622389
transform 1 0 4572 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4816
timestamp 1677622389
transform 1 0 4644 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1677622389
transform 1 0 4572 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5506
timestamp 1677622389
transform 1 0 4596 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4832
timestamp 1677622389
transform 1 0 4604 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5507
timestamp 1677622389
transform 1 0 4676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1677622389
transform 1 0 4700 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4817
timestamp 1677622389
transform 1 0 4724 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5508
timestamp 1677622389
transform 1 0 4724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1677622389
transform 1 0 4780 0 1 2125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_52
timestamp 1677622389
transform 1 0 24 0 1 2070
box -10 -3 10 3
use FILL  FILL_5960
timestamp 1677622389
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_341
timestamp 1677622389
transform 1 0 80 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_391
timestamp 1677622389
transform -1 0 192 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5961
timestamp 1677622389
transform 1 0 192 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_239
timestamp 1677622389
transform 1 0 200 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5962
timestamp 1677622389
transform 1 0 240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5963
timestamp 1677622389
transform 1 0 248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5964
timestamp 1677622389
transform 1 0 256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5965
timestamp 1677622389
transform 1 0 264 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_392
timestamp 1677622389
transform -1 0 288 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5966
timestamp 1677622389
transform 1 0 288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5967
timestamp 1677622389
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5968
timestamp 1677622389
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_240
timestamp 1677622389
transform -1 0 352 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5969
timestamp 1677622389
transform 1 0 352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5971
timestamp 1677622389
transform 1 0 360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5982
timestamp 1677622389
transform 1 0 368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5983
timestamp 1677622389
transform 1 0 376 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_241
timestamp 1677622389
transform 1 0 384 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5984
timestamp 1677622389
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5985
timestamp 1677622389
transform 1 0 432 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_394
timestamp 1677622389
transform 1 0 440 0 -1 2170
box -9 -3 26 105
use AOI22X1  AOI22X1_242
timestamp 1677622389
transform 1 0 456 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5986
timestamp 1677622389
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5987
timestamp 1677622389
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5988
timestamp 1677622389
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5989
timestamp 1677622389
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_228
timestamp 1677622389
transform -1 0 568 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5990
timestamp 1677622389
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5991
timestamp 1677622389
transform 1 0 576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5992
timestamp 1677622389
transform 1 0 584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5993
timestamp 1677622389
transform 1 0 592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5994
timestamp 1677622389
transform 1 0 600 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1677622389
transform -1 0 640 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5995
timestamp 1677622389
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_395
timestamp 1677622389
transform 1 0 648 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5996
timestamp 1677622389
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5998
timestamp 1677622389
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6000
timestamp 1677622389
transform 1 0 680 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_343
timestamp 1677622389
transform 1 0 688 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6006
timestamp 1677622389
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6008
timestamp 1677622389
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6010
timestamp 1677622389
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6012
timestamp 1677622389
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6014
timestamp 1677622389
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6015
timestamp 1677622389
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6016
timestamp 1677622389
transform 1 0 832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6017
timestamp 1677622389
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6018
timestamp 1677622389
transform 1 0 848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6019
timestamp 1677622389
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6020
timestamp 1677622389
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6021
timestamp 1677622389
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_396
timestamp 1677622389
transform -1 0 896 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6022
timestamp 1677622389
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6023
timestamp 1677622389
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6024
timestamp 1677622389
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6026
timestamp 1677622389
transform 1 0 920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6028
timestamp 1677622389
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6030
timestamp 1677622389
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6032
timestamp 1677622389
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6034
timestamp 1677622389
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_245
timestamp 1677622389
transform 1 0 960 0 -1 2170
box -8 -3 46 105
use M3_M2  M3_M2_4889
timestamp 1677622389
transform 1 0 1012 0 1 2075
box -3 -3 3 3
use FILL  FILL_6036
timestamp 1677622389
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6038
timestamp 1677622389
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6040
timestamp 1677622389
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4890
timestamp 1677622389
transform 1 0 1036 0 1 2075
box -3 -3 3 3
use FILL  FILL_6042
timestamp 1677622389
transform 1 0 1024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6044
timestamp 1677622389
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6046
timestamp 1677622389
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6047
timestamp 1677622389
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6048
timestamp 1677622389
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6049
timestamp 1677622389
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4891
timestamp 1677622389
transform 1 0 1084 0 1 2075
box -3 -3 3 3
use FILL  FILL_6051
timestamp 1677622389
transform 1 0 1072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6053
timestamp 1677622389
transform 1 0 1080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6055
timestamp 1677622389
transform 1 0 1088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6057
timestamp 1677622389
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6059
timestamp 1677622389
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_116
timestamp 1677622389
transform 1 0 1112 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6065
timestamp 1677622389
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6066
timestamp 1677622389
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6067
timestamp 1677622389
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6068
timestamp 1677622389
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6069
timestamp 1677622389
transform 1 0 1176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6071
timestamp 1677622389
transform 1 0 1184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6073
timestamp 1677622389
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6075
timestamp 1677622389
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6077
timestamp 1677622389
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6079
timestamp 1677622389
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6081
timestamp 1677622389
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6083
timestamp 1677622389
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6085
timestamp 1677622389
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6088
timestamp 1677622389
transform 1 0 1248 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4892
timestamp 1677622389
transform 1 0 1268 0 1 2075
box -3 -3 3 3
use FILL  FILL_6089
timestamp 1677622389
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6090
timestamp 1677622389
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6091
timestamp 1677622389
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6092
timestamp 1677622389
transform 1 0 1280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6093
timestamp 1677622389
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6095
timestamp 1677622389
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6097
timestamp 1677622389
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6099
timestamp 1677622389
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6101
timestamp 1677622389
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6103
timestamp 1677622389
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6106
timestamp 1677622389
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6107
timestamp 1677622389
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6108
timestamp 1677622389
transform 1 0 1352 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_118
timestamp 1677622389
transform -1 0 1392 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6109
timestamp 1677622389
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6110
timestamp 1677622389
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6111
timestamp 1677622389
transform 1 0 1408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6112
timestamp 1677622389
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6113
timestamp 1677622389
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6114
timestamp 1677622389
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6115
timestamp 1677622389
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6117
timestamp 1677622389
transform 1 0 1448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6119
timestamp 1677622389
transform 1 0 1456 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_230
timestamp 1677622389
transform 1 0 1464 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6122
timestamp 1677622389
transform 1 0 1504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6123
timestamp 1677622389
transform 1 0 1512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6125
timestamp 1677622389
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6127
timestamp 1677622389
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6134
timestamp 1677622389
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_397
timestamp 1677622389
transform -1 0 1560 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6135
timestamp 1677622389
transform 1 0 1560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6136
timestamp 1677622389
transform 1 0 1568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6137
timestamp 1677622389
transform 1 0 1576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6138
timestamp 1677622389
transform 1 0 1584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6139
timestamp 1677622389
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6140
timestamp 1677622389
transform 1 0 1600 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_64
timestamp 1677622389
transform -1 0 1632 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6141
timestamp 1677622389
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6142
timestamp 1677622389
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_65
timestamp 1677622389
transform 1 0 1648 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6143
timestamp 1677622389
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6145
timestamp 1677622389
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_66
timestamp 1677622389
transform 1 0 1688 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6148
timestamp 1677622389
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6149
timestamp 1677622389
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6150
timestamp 1677622389
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6151
timestamp 1677622389
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6169
timestamp 1677622389
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_347
timestamp 1677622389
transform -1 0 1848 0 -1 2170
box -8 -3 104 105
use BUFX2  BUFX2_67
timestamp 1677622389
transform 1 0 1848 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6170
timestamp 1677622389
transform 1 0 1872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6172
timestamp 1677622389
transform 1 0 1880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6174
timestamp 1677622389
transform 1 0 1888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6176
timestamp 1677622389
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6178
timestamp 1677622389
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6181
timestamp 1677622389
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6182
timestamp 1677622389
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6183
timestamp 1677622389
transform 1 0 1928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6184
timestamp 1677622389
transform 1 0 1936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6185
timestamp 1677622389
transform 1 0 1944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6186
timestamp 1677622389
transform 1 0 1952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6187
timestamp 1677622389
transform 1 0 1960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6189
timestamp 1677622389
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6191
timestamp 1677622389
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6193
timestamp 1677622389
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6195
timestamp 1677622389
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6197
timestamp 1677622389
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6199
timestamp 1677622389
transform 1 0 2008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6206
timestamp 1677622389
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6207
timestamp 1677622389
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_246
timestamp 1677622389
transform -1 0 2072 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6208
timestamp 1677622389
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6212
timestamp 1677622389
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6213
timestamp 1677622389
transform 1 0 2088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6214
timestamp 1677622389
transform 1 0 2096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6215
timestamp 1677622389
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6216
timestamp 1677622389
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6217
timestamp 1677622389
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6218
timestamp 1677622389
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6219
timestamp 1677622389
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6220
timestamp 1677622389
transform 1 0 2144 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_233
timestamp 1677622389
transform 1 0 2152 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6221
timestamp 1677622389
transform 1 0 2192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6222
timestamp 1677622389
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4893
timestamp 1677622389
transform 1 0 2220 0 1 2075
box -3 -3 3 3
use FILL  FILL_6223
timestamp 1677622389
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6224
timestamp 1677622389
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6225
timestamp 1677622389
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6226
timestamp 1677622389
transform 1 0 2232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6227
timestamp 1677622389
transform 1 0 2240 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4894
timestamp 1677622389
transform 1 0 2292 0 1 2075
box -3 -3 3 3
use OAI22X1  OAI22X1_234
timestamp 1677622389
transform -1 0 2288 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6228
timestamp 1677622389
transform 1 0 2288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6230
timestamp 1677622389
transform 1 0 2296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6232
timestamp 1677622389
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6234
timestamp 1677622389
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6236
timestamp 1677622389
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6238
timestamp 1677622389
transform 1 0 2328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6245
timestamp 1677622389
transform 1 0 2336 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4895
timestamp 1677622389
transform 1 0 2364 0 1 2075
box -3 -3 3 3
use AND2X2  AND2X2_15
timestamp 1677622389
transform -1 0 2376 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6246
timestamp 1677622389
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6247
timestamp 1677622389
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6248
timestamp 1677622389
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6249
timestamp 1677622389
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6250
timestamp 1677622389
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6251
timestamp 1677622389
transform 1 0 2416 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_235
timestamp 1677622389
transform 1 0 2424 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6257
timestamp 1677622389
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6258
timestamp 1677622389
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6259
timestamp 1677622389
transform 1 0 2480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6260
timestamp 1677622389
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6261
timestamp 1677622389
transform 1 0 2496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6262
timestamp 1677622389
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6263
timestamp 1677622389
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_16
timestamp 1677622389
transform 1 0 2520 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6264
timestamp 1677622389
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6266
timestamp 1677622389
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6268
timestamp 1677622389
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6270
timestamp 1677622389
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6272
timestamp 1677622389
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6276
timestamp 1677622389
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6277
timestamp 1677622389
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_249
timestamp 1677622389
transform 1 0 2608 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6278
timestamp 1677622389
transform 1 0 2648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6280
timestamp 1677622389
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6282
timestamp 1677622389
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6284
timestamp 1677622389
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6287
timestamp 1677622389
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_400
timestamp 1677622389
transform 1 0 2688 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6288
timestamp 1677622389
transform 1 0 2704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6290
timestamp 1677622389
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6293
timestamp 1677622389
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6294
timestamp 1677622389
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6295
timestamp 1677622389
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6296
timestamp 1677622389
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_59
timestamp 1677622389
transform 1 0 2752 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6297
timestamp 1677622389
transform 1 0 2776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6298
timestamp 1677622389
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6299
timestamp 1677622389
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6300
timestamp 1677622389
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_119
timestamp 1677622389
transform 1 0 2808 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6301
timestamp 1677622389
transform 1 0 2840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6302
timestamp 1677622389
transform 1 0 2848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6304
timestamp 1677622389
transform 1 0 2856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6306
timestamp 1677622389
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6308
timestamp 1677622389
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6313
timestamp 1677622389
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_121
timestamp 1677622389
transform -1 0 2920 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6314
timestamp 1677622389
transform 1 0 2920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6315
timestamp 1677622389
transform 1 0 2928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6316
timestamp 1677622389
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6318
timestamp 1677622389
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6320
timestamp 1677622389
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1677622389
transform 1 0 2960 0 -1 2170
box -8 -3 32 105
use AND2X2  AND2X2_17
timestamp 1677622389
transform 1 0 2984 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6326
timestamp 1677622389
transform 1 0 3016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6327
timestamp 1677622389
transform 1 0 3024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6328
timestamp 1677622389
transform 1 0 3032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6329
timestamp 1677622389
transform 1 0 3040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6330
timestamp 1677622389
transform 1 0 3048 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_401
timestamp 1677622389
transform -1 0 3072 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6331
timestamp 1677622389
transform 1 0 3072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6332
timestamp 1677622389
transform 1 0 3080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6333
timestamp 1677622389
transform 1 0 3088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6335
timestamp 1677622389
transform 1 0 3096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6337
timestamp 1677622389
transform 1 0 3104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6345
timestamp 1677622389
transform 1 0 3112 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_236
timestamp 1677622389
transform -1 0 3160 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6346
timestamp 1677622389
transform 1 0 3160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6348
timestamp 1677622389
transform 1 0 3168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6355
timestamp 1677622389
transform 1 0 3176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6356
timestamp 1677622389
transform 1 0 3184 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_353
timestamp 1677622389
transform 1 0 3192 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6357
timestamp 1677622389
transform 1 0 3288 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_402
timestamp 1677622389
transform 1 0 3296 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6361
timestamp 1677622389
transform 1 0 3312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6363
timestamp 1677622389
transform 1 0 3320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6369
timestamp 1677622389
transform 1 0 3328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6370
timestamp 1677622389
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6371
timestamp 1677622389
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6372
timestamp 1677622389
transform 1 0 3352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6373
timestamp 1677622389
transform 1 0 3360 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_18
timestamp 1677622389
transform 1 0 3368 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6374
timestamp 1677622389
transform 1 0 3400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6376
timestamp 1677622389
transform 1 0 3408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6377
timestamp 1677622389
transform 1 0 3416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6378
timestamp 1677622389
transform 1 0 3424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6379
timestamp 1677622389
transform 1 0 3432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6380
timestamp 1677622389
transform 1 0 3440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6382
timestamp 1677622389
transform 1 0 3448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6384
timestamp 1677622389
transform 1 0 3456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6386
timestamp 1677622389
transform 1 0 3464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6388
timestamp 1677622389
transform 1 0 3472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6390
timestamp 1677622389
transform 1 0 3480 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_39
timestamp 1677622389
transform -1 0 3520 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6391
timestamp 1677622389
transform 1 0 3520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6393
timestamp 1677622389
transform 1 0 3528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6395
timestamp 1677622389
transform 1 0 3536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6397
timestamp 1677622389
transform 1 0 3544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6399
timestamp 1677622389
transform 1 0 3552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6407
timestamp 1677622389
transform 1 0 3560 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_237
timestamp 1677622389
transform -1 0 3608 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6408
timestamp 1677622389
transform 1 0 3608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6409
timestamp 1677622389
transform 1 0 3616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6410
timestamp 1677622389
transform 1 0 3624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6412
timestamp 1677622389
transform 1 0 3632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6414
timestamp 1677622389
transform 1 0 3640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6424
timestamp 1677622389
transform 1 0 3648 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_355
timestamp 1677622389
transform -1 0 3752 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6425
timestamp 1677622389
transform 1 0 3752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6426
timestamp 1677622389
transform 1 0 3760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6427
timestamp 1677622389
transform 1 0 3768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6428
timestamp 1677622389
transform 1 0 3776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6429
timestamp 1677622389
transform 1 0 3784 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_239
timestamp 1677622389
transform 1 0 3792 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6430
timestamp 1677622389
transform 1 0 3832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6431
timestamp 1677622389
transform 1 0 3840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6432
timestamp 1677622389
transform 1 0 3848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6433
timestamp 1677622389
transform 1 0 3856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6434
timestamp 1677622389
transform 1 0 3864 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_406
timestamp 1677622389
transform 1 0 3872 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6436
timestamp 1677622389
transform 1 0 3888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6438
timestamp 1677622389
transform 1 0 3896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6440
timestamp 1677622389
transform 1 0 3904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6442
timestamp 1677622389
transform 1 0 3912 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_241
timestamp 1677622389
transform 1 0 3920 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6445
timestamp 1677622389
transform 1 0 3960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6446
timestamp 1677622389
transform 1 0 3968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6448
timestamp 1677622389
transform 1 0 3976 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_356
timestamp 1677622389
transform 1 0 3984 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_407
timestamp 1677622389
transform 1 0 4080 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6459
timestamp 1677622389
transform 1 0 4096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6461
timestamp 1677622389
transform 1 0 4104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6468
timestamp 1677622389
transform 1 0 4112 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_243
timestamp 1677622389
transform -1 0 4160 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6469
timestamp 1677622389
transform 1 0 4160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6470
timestamp 1677622389
transform 1 0 4168 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_408
timestamp 1677622389
transform -1 0 4192 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6471
timestamp 1677622389
transform 1 0 4192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6472
timestamp 1677622389
transform 1 0 4200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6473
timestamp 1677622389
transform 1 0 4208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6474
timestamp 1677622389
transform 1 0 4216 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_409
timestamp 1677622389
transform -1 0 4240 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6475
timestamp 1677622389
transform 1 0 4240 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_244
timestamp 1677622389
transform 1 0 4248 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6476
timestamp 1677622389
transform 1 0 4288 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_358
timestamp 1677622389
transform 1 0 4296 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6486
timestamp 1677622389
transform 1 0 4392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6487
timestamp 1677622389
transform 1 0 4400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6488
timestamp 1677622389
transform 1 0 4408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6489
timestamp 1677622389
transform 1 0 4416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6501
timestamp 1677622389
transform 1 0 4424 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_360
timestamp 1677622389
transform -1 0 4528 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6502
timestamp 1677622389
transform 1 0 4528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6503
timestamp 1677622389
transform 1 0 4536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6504
timestamp 1677622389
transform 1 0 4544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6505
timestamp 1677622389
transform 1 0 4552 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_361
timestamp 1677622389
transform 1 0 4560 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6506
timestamp 1677622389
transform 1 0 4656 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_413
timestamp 1677622389
transform 1 0 4664 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6507
timestamp 1677622389
transform 1 0 4680 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_362
timestamp 1677622389
transform 1 0 4688 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6508
timestamp 1677622389
transform 1 0 4784 0 -1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_53
timestamp 1677622389
transform 1 0 4843 0 1 2070
box -10 -3 10 3
use M3_M2  M3_M2_4927
timestamp 1677622389
transform 1 0 172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1677622389
transform 1 0 140 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1677622389
transform 1 0 180 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5532
timestamp 1677622389
transform 1 0 140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1677622389
transform 1 0 172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1677622389
transform 1 0 180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1677622389
transform 1 0 92 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5008
timestamp 1677622389
transform 1 0 92 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1677622389
transform 1 0 212 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1677622389
transform 1 0 204 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1677622389
transform 1 0 236 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5535
timestamp 1677622389
transform 1 0 204 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1677622389
transform 1 0 220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1677622389
transform 1 0 204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1677622389
transform 1 0 212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1677622389
transform 1 0 228 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4911
timestamp 1677622389
transform 1 0 252 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5537
timestamp 1677622389
transform 1 0 252 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5009
timestamp 1677622389
transform 1 0 252 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5538
timestamp 1677622389
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1677622389
transform 1 0 284 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5010
timestamp 1677622389
transform 1 0 284 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1677622389
transform 1 0 396 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1677622389
transform 1 0 340 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1677622389
transform 1 0 388 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1677622389
transform 1 0 420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1677622389
transform 1 0 516 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1677622389
transform 1 0 548 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1677622389
transform 1 0 556 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1677622389
transform 1 0 524 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1677622389
transform 1 0 564 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5539
timestamp 1677622389
transform 1 0 340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1677622389
transform 1 0 388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1677622389
transform 1 0 396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1677622389
transform 1 0 412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1677622389
transform 1 0 428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1677622389
transform 1 0 468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1677622389
transform 1 0 524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1677622389
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1677622389
transform 1 0 308 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4992
timestamp 1677622389
transform 1 0 372 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1677622389
transform 1 0 308 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5630
timestamp 1677622389
transform 1 0 404 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1677622389
transform 1 0 420 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4993
timestamp 1677622389
transform 1 0 428 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1677622389
transform 1 0 548 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5547
timestamp 1677622389
transform 1 0 556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1677622389
transform 1 0 444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1677622389
transform 1 0 532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1677622389
transform 1 0 548 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1677622389
transform 1 0 564 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1677622389
transform 1 0 572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5011
timestamp 1677622389
transform 1 0 420 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1677622389
transform 1 0 444 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1677622389
transform 1 0 548 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1677622389
transform 1 0 572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1677622389
transform 1 0 604 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1677622389
transform 1 0 636 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1677622389
transform 1 0 628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1677622389
transform 1 0 612 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5548
timestamp 1677622389
transform 1 0 620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1677622389
transform 1 0 612 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4994
timestamp 1677622389
transform 1 0 620 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5549
timestamp 1677622389
transform 1 0 636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1677622389
transform 1 0 628 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4987
timestamp 1677622389
transform 1 0 644 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5550
timestamp 1677622389
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5013
timestamp 1677622389
transform 1 0 668 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1677622389
transform 1 0 684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1677622389
transform 1 0 684 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5639
timestamp 1677622389
transform 1 0 684 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4930
timestamp 1677622389
transform 1 0 748 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1677622389
transform 1 0 748 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5551
timestamp 1677622389
transform 1 0 716 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4989
timestamp 1677622389
transform 1 0 724 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5552
timestamp 1677622389
transform 1 0 732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1677622389
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1677622389
transform 1 0 756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1677622389
transform 1 0 716 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4953
timestamp 1677622389
transform 1 0 772 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5641
timestamp 1677622389
transform 1 0 764 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4923
timestamp 1677622389
transform 1 0 804 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1677622389
transform 1 0 804 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1677622389
transform 1 0 836 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5555
timestamp 1677622389
transform 1 0 820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1677622389
transform 1 0 836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1677622389
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1677622389
transform 1 0 844 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_4924
timestamp 1677622389
transform 1 0 852 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1677622389
transform 1 0 844 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5643
timestamp 1677622389
transform 1 0 860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1677622389
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4995
timestamp 1677622389
transform 1 0 908 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5701
timestamp 1677622389
transform 1 0 908 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_4925
timestamp 1677622389
transform 1 0 972 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1677622389
transform 1 0 972 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1677622389
transform 1 0 996 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5645
timestamp 1677622389
transform 1 0 1020 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4956
timestamp 1677622389
transform 1 0 1036 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5557
timestamp 1677622389
transform 1 0 1036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1677622389
transform 1 0 1060 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4957
timestamp 1677622389
transform 1 0 1140 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1677622389
transform 1 0 1236 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5558
timestamp 1677622389
transform 1 0 1236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1677622389
transform 1 0 1236 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5014
timestamp 1677622389
transform 1 0 1236 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5559
timestamp 1677622389
transform 1 0 1252 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5015
timestamp 1677622389
transform 1 0 1252 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1677622389
transform 1 0 1284 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1677622389
transform 1 0 1276 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5648
timestamp 1677622389
transform 1 0 1276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1677622389
transform 1 0 1308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1677622389
transform 1 0 1348 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1677622389
transform 1 0 1340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1677622389
transform 1 0 1388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1677622389
transform 1 0 1428 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4960
timestamp 1677622389
transform 1 0 1460 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1677622389
transform 1 0 1476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1677622389
transform 1 0 1492 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5563
timestamp 1677622389
transform 1 0 1476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1677622389
transform 1 0 1460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1677622389
transform 1 0 1468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1677622389
transform 1 0 1516 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1677622389
transform 1 0 1548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5016
timestamp 1677622389
transform 1 0 1548 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1677622389
transform 1 0 1564 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1677622389
transform 1 0 1564 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1677622389
transform 1 0 1612 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5653
timestamp 1677622389
transform 1 0 1612 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4900
timestamp 1677622389
transform 1 0 1628 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5565
timestamp 1677622389
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4901
timestamp 1677622389
transform 1 0 1740 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5566
timestamp 1677622389
transform 1 0 1668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1677622389
transform 1 0 1716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1677622389
transform 1 0 1764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1677622389
transform 1 0 1748 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5018
timestamp 1677622389
transform 1 0 1748 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1677622389
transform 1 0 1780 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5655
timestamp 1677622389
transform 1 0 1780 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4902
timestamp 1677622389
transform 1 0 1828 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5569
timestamp 1677622389
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1677622389
transform 1 0 1916 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4934
timestamp 1677622389
transform 1 0 1940 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5571
timestamp 1677622389
transform 1 0 1948 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4962
timestamp 1677622389
transform 1 0 1972 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5572
timestamp 1677622389
transform 1 0 1972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1677622389
transform 1 0 1932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1677622389
transform 1 0 1940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1677622389
transform 1 0 1956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1677622389
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4935
timestamp 1677622389
transform 1 0 2060 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5573
timestamp 1677622389
transform 1 0 2052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1677622389
transform 1 0 2020 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4915
timestamp 1677622389
transform 1 0 2148 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1677622389
transform 1 0 2172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1677622389
transform 1 0 2148 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1677622389
transform 1 0 2188 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5574
timestamp 1677622389
transform 1 0 2148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1677622389
transform 1 0 2164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1677622389
transform 1 0 2180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1677622389
transform 1 0 2188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1677622389
transform 1 0 2156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1677622389
transform 1 0 2172 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5037
timestamp 1677622389
transform 1 0 2212 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1677622389
transform 1 0 2252 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1677622389
transform 1 0 2300 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1677622389
transform 1 0 2276 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5578
timestamp 1677622389
transform 1 0 2276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1677622389
transform 1 0 2292 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4996
timestamp 1677622389
transform 1 0 2268 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5518
timestamp 1677622389
transform 1 0 2316 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_4966
timestamp 1677622389
transform 1 0 2316 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5580
timestamp 1677622389
transform 1 0 2316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1677622389
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1677622389
transform 1 0 2284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1677622389
transform 1 0 2300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1677622389
transform 1 0 2308 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5020
timestamp 1677622389
transform 1 0 2308 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5519
timestamp 1677622389
transform 1 0 2340 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5038
timestamp 1677622389
transform 1 0 2340 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1677622389
transform 1 0 2364 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1677622389
transform 1 0 2388 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1677622389
transform 1 0 2428 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1677622389
transform 1 0 2436 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5581
timestamp 1677622389
transform 1 0 2412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1677622389
transform 1 0 2428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1677622389
transform 1 0 2404 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4998
timestamp 1677622389
transform 1 0 2412 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5668
timestamp 1677622389
transform 1 0 2436 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4917
timestamp 1677622389
transform 1 0 2508 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1677622389
transform 1 0 2508 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5669
timestamp 1677622389
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4918
timestamp 1677622389
transform 1 0 2524 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1677622389
transform 1 0 2556 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5583
timestamp 1677622389
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4904
timestamp 1677622389
transform 1 0 2580 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5584
timestamp 1677622389
transform 1 0 2580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1677622389
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4905
timestamp 1677622389
transform 1 0 2620 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1677622389
transform 1 0 2604 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5585
timestamp 1677622389
transform 1 0 2604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1677622389
transform 1 0 2620 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4969
timestamp 1677622389
transform 1 0 2644 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5671
timestamp 1677622389
transform 1 0 2644 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4906
timestamp 1677622389
transform 1 0 2660 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1677622389
transform 1 0 2684 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1677622389
transform 1 0 2740 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5587
timestamp 1677622389
transform 1 0 2684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1677622389
transform 1 0 2740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1677622389
transform 1 0 2660 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4907
timestamp 1677622389
transform 1 0 2780 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1677622389
transform 1 0 2780 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5589
timestamp 1677622389
transform 1 0 2780 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4972
timestamp 1677622389
transform 1 0 2804 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5673
timestamp 1677622389
transform 1 0 2796 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5021
timestamp 1677622389
transform 1 0 2780 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5525
timestamp 1677622389
transform 1 0 2892 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1677622389
transform 1 0 2908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1677622389
transform 1 0 2956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1677622389
transform 1 0 3012 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5022
timestamp 1677622389
transform 1 0 3012 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5591
timestamp 1677622389
transform 1 0 3028 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4973
timestamp 1677622389
transform 1 0 3068 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5592
timestamp 1677622389
transform 1 0 3044 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4974
timestamp 1677622389
transform 1 0 3084 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5593
timestamp 1677622389
transform 1 0 3084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1677622389
transform 1 0 3052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1677622389
transform 1 0 3068 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1677622389
transform 1 0 3076 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5023
timestamp 1677622389
transform 1 0 3076 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1677622389
transform 1 0 3100 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1677622389
transform 1 0 3140 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5594
timestamp 1677622389
transform 1 0 3124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1677622389
transform 1 0 3140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1677622389
transform 1 0 3116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1677622389
transform 1 0 3132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1677622389
transform 1 0 3156 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5000
timestamp 1677622389
transform 1 0 3156 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5681
timestamp 1677622389
transform 1 0 3188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1677622389
transform 1 0 3204 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1677622389
transform 1 0 3220 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_4908
timestamp 1677622389
transform 1 0 3260 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1677622389
transform 1 0 3252 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5521
timestamp 1677622389
transform 1 0 3260 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_4976
timestamp 1677622389
transform 1 0 3268 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5596
timestamp 1677622389
transform 1 0 3268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1677622389
transform 1 0 3324 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1677622389
transform 1 0 3308 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1677622389
transform 1 0 3316 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_4990
timestamp 1677622389
transform 1 0 3308 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1677622389
transform 1 0 3356 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5530
timestamp 1677622389
transform 1 0 3340 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5001
timestamp 1677622389
transform 1 0 3324 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1677622389
transform 1 0 3348 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1677622389
transform 1 0 3412 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1677622389
transform 1 0 3420 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5523
timestamp 1677622389
transform 1 0 3444 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1677622389
transform 1 0 3452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1677622389
transform 1 0 3484 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1677622389
transform 1 0 3492 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5002
timestamp 1677622389
transform 1 0 3492 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5599
timestamp 1677622389
transform 1 0 3564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1677622389
transform 1 0 3588 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5024
timestamp 1677622389
transform 1 0 3564 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1677622389
transform 1 0 3588 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5683
timestamp 1677622389
transform 1 0 3604 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4942
timestamp 1677622389
transform 1 0 3620 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5600
timestamp 1677622389
transform 1 0 3652 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5003
timestamp 1677622389
transform 1 0 3652 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5684
timestamp 1677622389
transform 1 0 3660 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1677622389
transform 1 0 3676 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5025
timestamp 1677622389
transform 1 0 3660 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1677622389
transform 1 0 3668 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5601
timestamp 1677622389
transform 1 0 3700 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4978
timestamp 1677622389
transform 1 0 3764 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5602
timestamp 1677622389
transform 1 0 3764 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4991
timestamp 1677622389
transform 1 0 3780 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5686
timestamp 1677622389
transform 1 0 3716 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5042
timestamp 1677622389
transform 1 0 3716 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1677622389
transform 1 0 3812 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1677622389
transform 1 0 3836 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5603
timestamp 1677622389
transform 1 0 3860 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5004
timestamp 1677622389
transform 1 0 3924 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1677622389
transform 1 0 3940 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5604
timestamp 1677622389
transform 1 0 3964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1677622389
transform 1 0 4004 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5005
timestamp 1677622389
transform 1 0 4004 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1677622389
transform 1 0 4108 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5606
timestamp 1677622389
transform 1 0 4084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1677622389
transform 1 0 4100 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1677622389
transform 1 0 4108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1677622389
transform 1 0 4052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1677622389
transform 1 0 4068 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1677622389
transform 1 0 4076 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5026
timestamp 1677622389
transform 1 0 4076 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1677622389
transform 1 0 4108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1677622389
transform 1 0 4100 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5609
timestamp 1677622389
transform 1 0 4132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1677622389
transform 1 0 4116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1677622389
transform 1 0 4124 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1677622389
transform 1 0 4244 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4980
timestamp 1677622389
transform 1 0 4332 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1677622389
transform 1 0 4348 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5611
timestamp 1677622389
transform 1 0 4284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1677622389
transform 1 0 4348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1677622389
transform 1 0 4380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1677622389
transform 1 0 4444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1677622389
transform 1 0 4460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1677622389
transform 1 0 4332 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1677622389
transform 1 0 4428 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5028
timestamp 1677622389
transform 1 0 4428 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1677622389
transform 1 0 4460 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1677622389
transform 1 0 4516 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5616
timestamp 1677622389
transform 1 0 4484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1677622389
transform 1 0 4500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1677622389
transform 1 0 4516 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1677622389
transform 1 0 4468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1677622389
transform 1 0 4476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1677622389
transform 1 0 4492 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5007
timestamp 1677622389
transform 1 0 4500 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1677622389
transform 1 0 4572 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1677622389
transform 1 0 4628 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5619
timestamp 1677622389
transform 1 0 4564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1677622389
transform 1 0 4620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1677622389
transform 1 0 4628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1677622389
transform 1 0 4540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1677622389
transform 1 0 4636 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5029
timestamp 1677622389
transform 1 0 4540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1677622389
transform 1 0 4628 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5622
timestamp 1677622389
transform 1 0 4732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1677622389
transform 1 0 4788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1677622389
transform 1 0 4708 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5031
timestamp 1677622389
transform 1 0 4732 0 1 1995
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_54
timestamp 1677622389
transform 1 0 48 0 1 1970
box -10 -3 10 3
use FILL  FILL_6509
timestamp 1677622389
transform 1 0 72 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_363
timestamp 1677622389
transform 1 0 80 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_414
timestamp 1677622389
transform -1 0 192 0 1 1970
box -9 -3 26 105
use FILL  FILL_6511
timestamp 1677622389
transform 1 0 192 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_254
timestamp 1677622389
transform -1 0 240 0 1 1970
box -8 -3 46 105
use FILL  FILL_6512
timestamp 1677622389
transform 1 0 240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6513
timestamp 1677622389
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6517
timestamp 1677622389
transform 1 0 256 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_71
timestamp 1677622389
transform 1 0 264 0 1 1970
box -5 -3 28 105
use FILL  FILL_6519
timestamp 1677622389
transform 1 0 288 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_365
timestamp 1677622389
transform 1 0 296 0 1 1970
box -8 -3 104 105
use AOI22X1  AOI22X1_256
timestamp 1677622389
transform 1 0 392 0 1 1970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_366
timestamp 1677622389
transform 1 0 432 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5045
timestamp 1677622389
transform 1 0 548 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_248
timestamp 1677622389
transform -1 0 568 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5046
timestamp 1677622389
transform 1 0 580 0 1 1975
box -3 -3 3 3
use FILL  FILL_6520
timestamp 1677622389
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6537
timestamp 1677622389
transform 1 0 576 0 1 1970
box -8 -3 16 105
use FILL  FILL_6539
timestamp 1677622389
transform 1 0 584 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_249
timestamp 1677622389
transform 1 0 592 0 1 1970
box -8 -3 46 105
use FILL  FILL_6541
timestamp 1677622389
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6542
timestamp 1677622389
transform 1 0 640 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5047
timestamp 1677622389
transform 1 0 684 0 1 1975
box -3 -3 3 3
use AND2X2  AND2X2_20
timestamp 1677622389
transform -1 0 680 0 1 1970
box -8 -3 40 105
use FILL  FILL_6543
timestamp 1677622389
transform 1 0 680 0 1 1970
box -8 -3 16 105
use FILL  FILL_6544
timestamp 1677622389
transform 1 0 688 0 1 1970
box -8 -3 16 105
use FILL  FILL_6545
timestamp 1677622389
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_6553
timestamp 1677622389
transform 1 0 704 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_257
timestamp 1677622389
transform 1 0 712 0 1 1970
box -8 -3 46 105
use FILL  FILL_6555
timestamp 1677622389
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6556
timestamp 1677622389
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_6557
timestamp 1677622389
transform 1 0 768 0 1 1970
box -8 -3 16 105
use FILL  FILL_6558
timestamp 1677622389
transform 1 0 776 0 1 1970
box -8 -3 16 105
use FILL  FILL_6559
timestamp 1677622389
transform 1 0 784 0 1 1970
box -8 -3 16 105
use FILL  FILL_6560
timestamp 1677622389
transform 1 0 792 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_258
timestamp 1677622389
transform 1 0 800 0 1 1970
box -8 -3 46 105
use FILL  FILL_6561
timestamp 1677622389
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6562
timestamp 1677622389
transform 1 0 848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6563
timestamp 1677622389
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6567
timestamp 1677622389
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6569
timestamp 1677622389
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6571
timestamp 1677622389
transform 1 0 880 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_62
timestamp 1677622389
transform 1 0 888 0 1 1970
box -8 -3 32 105
use FILL  FILL_6573
timestamp 1677622389
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6578
timestamp 1677622389
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6579
timestamp 1677622389
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6580
timestamp 1677622389
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6581
timestamp 1677622389
transform 1 0 944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6582
timestamp 1677622389
transform 1 0 952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6583
timestamp 1677622389
transform 1 0 960 0 1 1970
box -8 -3 16 105
use FILL  FILL_6585
timestamp 1677622389
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_6587
timestamp 1677622389
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_6589
timestamp 1677622389
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_6591
timestamp 1677622389
transform 1 0 992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6593
timestamp 1677622389
transform 1 0 1000 0 1 1970
box -8 -3 16 105
use FILL  FILL_6595
timestamp 1677622389
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_6597
timestamp 1677622389
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_6599
timestamp 1677622389
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_63
timestamp 1677622389
transform 1 0 1032 0 1 1970
box -8 -3 32 105
use FILL  FILL_6601
timestamp 1677622389
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_6606
timestamp 1677622389
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_6608
timestamp 1677622389
transform 1 0 1072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6610
timestamp 1677622389
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_6612
timestamp 1677622389
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use FILL  FILL_6614
timestamp 1677622389
transform 1 0 1096 0 1 1970
box -8 -3 16 105
use FILL  FILL_6616
timestamp 1677622389
transform 1 0 1104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6618
timestamp 1677622389
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_6619
timestamp 1677622389
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_6620
timestamp 1677622389
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6622
timestamp 1677622389
transform 1 0 1136 0 1 1970
box -8 -3 16 105
use FILL  FILL_6624
timestamp 1677622389
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_6626
timestamp 1677622389
transform 1 0 1152 0 1 1970
box -8 -3 16 105
use FILL  FILL_6628
timestamp 1677622389
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6629
timestamp 1677622389
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6630
timestamp 1677622389
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6631
timestamp 1677622389
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6632
timestamp 1677622389
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6633
timestamp 1677622389
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_6634
timestamp 1677622389
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_6635
timestamp 1677622389
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6636
timestamp 1677622389
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6637
timestamp 1677622389
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_122
timestamp 1677622389
transform 1 0 1240 0 1 1970
box -8 -3 34 105
use FILL  FILL_6638
timestamp 1677622389
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use FILL  FILL_6642
timestamp 1677622389
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use FILL  FILL_6644
timestamp 1677622389
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6645
timestamp 1677622389
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6646
timestamp 1677622389
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_6647
timestamp 1677622389
transform 1 0 1312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6648
timestamp 1677622389
transform 1 0 1320 0 1 1970
box -8 -3 16 105
use FILL  FILL_6649
timestamp 1677622389
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_6652
timestamp 1677622389
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_6654
timestamp 1677622389
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_123
timestamp 1677622389
transform -1 0 1384 0 1 1970
box -8 -3 34 105
use FILL  FILL_6655
timestamp 1677622389
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6656
timestamp 1677622389
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6657
timestamp 1677622389
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_6658
timestamp 1677622389
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6659
timestamp 1677622389
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6660
timestamp 1677622389
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_6661
timestamp 1677622389
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6662
timestamp 1677622389
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6663
timestamp 1677622389
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5048
timestamp 1677622389
transform 1 0 1468 0 1 1975
box -3 -3 3 3
use FILL  FILL_6664
timestamp 1677622389
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1677622389
transform 1 0 1464 0 1 1970
box -8 -3 40 105
use FILL  FILL_6665
timestamp 1677622389
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6666
timestamp 1677622389
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_6667
timestamp 1677622389
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6668
timestamp 1677622389
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6677
timestamp 1677622389
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6678
timestamp 1677622389
transform 1 0 1536 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_76
timestamp 1677622389
transform -1 0 1568 0 1 1970
box -5 -3 28 105
use FILL  FILL_6679
timestamp 1677622389
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6683
timestamp 1677622389
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_6685
timestamp 1677622389
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_6687
timestamp 1677622389
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_6689
timestamp 1677622389
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_78
timestamp 1677622389
transform -1 0 1632 0 1 1970
box -5 -3 28 105
use FILL  FILL_6690
timestamp 1677622389
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6693
timestamp 1677622389
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6695
timestamp 1677622389
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_6697
timestamp 1677622389
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_371
timestamp 1677622389
transform -1 0 1760 0 1 1970
box -8 -3 104 105
use BUFX2  BUFX2_80
timestamp 1677622389
transform 1 0 1760 0 1 1970
box -5 -3 28 105
use FILL  FILL_6698
timestamp 1677622389
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_6714
timestamp 1677622389
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_6716
timestamp 1677622389
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_6717
timestamp 1677622389
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_6718
timestamp 1677622389
transform 1 0 1816 0 1 1970
box -8 -3 16 105
use FILL  FILL_6720
timestamp 1677622389
transform 1 0 1824 0 1 1970
box -8 -3 16 105
use FILL  FILL_6722
timestamp 1677622389
transform 1 0 1832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6723
timestamp 1677622389
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6724
timestamp 1677622389
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6725
timestamp 1677622389
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_422
timestamp 1677622389
transform -1 0 1880 0 1 1970
box -9 -3 26 105
use FILL  FILL_6726
timestamp 1677622389
transform 1 0 1880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6727
timestamp 1677622389
transform 1 0 1888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6728
timestamp 1677622389
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6729
timestamp 1677622389
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6730
timestamp 1677622389
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6731
timestamp 1677622389
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5049
timestamp 1677622389
transform 1 0 1972 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_260
timestamp 1677622389
transform 1 0 1928 0 1 1970
box -8 -3 46 105
use FILL  FILL_6732
timestamp 1677622389
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_6736
timestamp 1677622389
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_6738
timestamp 1677622389
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_6740
timestamp 1677622389
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6742
timestamp 1677622389
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5050
timestamp 1677622389
transform 1 0 2028 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_373
timestamp 1677622389
transform 1 0 2008 0 1 1970
box -8 -3 104 105
use FILL  FILL_6744
timestamp 1677622389
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6752
timestamp 1677622389
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_6754
timestamp 1677622389
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_6756
timestamp 1677622389
transform 1 0 2128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6758
timestamp 1677622389
transform 1 0 2136 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_261
timestamp 1677622389
transform -1 0 2184 0 1 1970
box -8 -3 46 105
use FILL  FILL_6759
timestamp 1677622389
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6767
timestamp 1677622389
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6769
timestamp 1677622389
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_6771
timestamp 1677622389
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_6773
timestamp 1677622389
transform 1 0 2216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6775
timestamp 1677622389
transform 1 0 2224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6777
timestamp 1677622389
transform 1 0 2232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6779
timestamp 1677622389
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6780
timestamp 1677622389
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6781
timestamp 1677622389
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6783
timestamp 1677622389
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_262
timestamp 1677622389
transform -1 0 2312 0 1 1970
box -8 -3 46 105
use FILL  FILL_6784
timestamp 1677622389
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6785
timestamp 1677622389
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_6786
timestamp 1677622389
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_6787
timestamp 1677622389
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5051
timestamp 1677622389
transform 1 0 2356 0 1 1975
box -3 -3 3 3
use FILL  FILL_6788
timestamp 1677622389
transform 1 0 2344 0 1 1970
box -8 -3 16 105
use FILL  FILL_6789
timestamp 1677622389
transform 1 0 2352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6790
timestamp 1677622389
transform 1 0 2360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6791
timestamp 1677622389
transform 1 0 2368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6794
timestamp 1677622389
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6796
timestamp 1677622389
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_263
timestamp 1677622389
transform -1 0 2432 0 1 1970
box -8 -3 46 105
use FILL  FILL_6797
timestamp 1677622389
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6798
timestamp 1677622389
transform 1 0 2440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6799
timestamp 1677622389
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6800
timestamp 1677622389
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_6801
timestamp 1677622389
transform 1 0 2464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6802
timestamp 1677622389
transform 1 0 2472 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5052
timestamp 1677622389
transform 1 0 2492 0 1 1975
box -3 -3 3 3
use FILL  FILL_6803
timestamp 1677622389
transform 1 0 2480 0 1 1970
box -8 -3 16 105
use FILL  FILL_6804
timestamp 1677622389
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5053
timestamp 1677622389
transform 1 0 2508 0 1 1975
box -3 -3 3 3
use FILL  FILL_6805
timestamp 1677622389
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_425
timestamp 1677622389
transform 1 0 2504 0 1 1970
box -9 -3 26 105
use FILL  FILL_6806
timestamp 1677622389
transform 1 0 2520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6811
timestamp 1677622389
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6813
timestamp 1677622389
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6815
timestamp 1677622389
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use FILL  FILL_6817
timestamp 1677622389
transform 1 0 2552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6819
timestamp 1677622389
transform 1 0 2560 0 1 1970
box -8 -3 16 105
use FILL  FILL_6820
timestamp 1677622389
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6821
timestamp 1677622389
transform 1 0 2576 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_264
timestamp 1677622389
transform 1 0 2584 0 1 1970
box -8 -3 46 105
use FILL  FILL_6822
timestamp 1677622389
transform 1 0 2624 0 1 1970
box -8 -3 16 105
use FILL  FILL_6827
timestamp 1677622389
transform 1 0 2632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6829
timestamp 1677622389
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5054
timestamp 1677622389
transform 1 0 2660 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1677622389
transform 1 0 2692 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_376
timestamp 1677622389
transform 1 0 2648 0 1 1970
box -8 -3 104 105
use FILL  FILL_6831
timestamp 1677622389
transform 1 0 2744 0 1 1970
box -8 -3 16 105
use FILL  FILL_6832
timestamp 1677622389
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6833
timestamp 1677622389
transform 1 0 2760 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_124
timestamp 1677622389
transform 1 0 2768 0 1 1970
box -8 -3 34 105
use FILL  FILL_6834
timestamp 1677622389
transform 1 0 2800 0 1 1970
box -8 -3 16 105
use FILL  FILL_6841
timestamp 1677622389
transform 1 0 2808 0 1 1970
box -8 -3 16 105
use FILL  FILL_6843
timestamp 1677622389
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use FILL  FILL_6845
timestamp 1677622389
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_6847
timestamp 1677622389
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6848
timestamp 1677622389
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6849
timestamp 1677622389
transform 1 0 2848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6850
timestamp 1677622389
transform 1 0 2856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6852
timestamp 1677622389
transform 1 0 2864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6854
timestamp 1677622389
transform 1 0 2872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6856
timestamp 1677622389
transform 1 0 2880 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_125
timestamp 1677622389
transform -1 0 2920 0 1 1970
box -8 -3 34 105
use FILL  FILL_6857
timestamp 1677622389
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6858
timestamp 1677622389
transform 1 0 2928 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5056
timestamp 1677622389
transform 1 0 2948 0 1 1975
box -3 -3 3 3
use FILL  FILL_6862
timestamp 1677622389
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6864
timestamp 1677622389
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6865
timestamp 1677622389
transform 1 0 2952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6866
timestamp 1677622389
transform 1 0 2960 0 1 1970
box -8 -3 16 105
use FILL  FILL_6867
timestamp 1677622389
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_428
timestamp 1677622389
transform 1 0 2976 0 1 1970
box -9 -3 26 105
use FILL  FILL_6868
timestamp 1677622389
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6869
timestamp 1677622389
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_6870
timestamp 1677622389
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_6871
timestamp 1677622389
transform 1 0 3016 0 1 1970
box -8 -3 16 105
use FILL  FILL_6872
timestamp 1677622389
transform 1 0 3024 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_250
timestamp 1677622389
transform -1 0 3072 0 1 1970
box -8 -3 46 105
use FILL  FILL_6873
timestamp 1677622389
transform 1 0 3072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6874
timestamp 1677622389
transform 1 0 3080 0 1 1970
box -8 -3 16 105
use FILL  FILL_6875
timestamp 1677622389
transform 1 0 3088 0 1 1970
box -8 -3 16 105
use FILL  FILL_6876
timestamp 1677622389
transform 1 0 3096 0 1 1970
box -8 -3 16 105
use FILL  FILL_6877
timestamp 1677622389
transform 1 0 3104 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5057
timestamp 1677622389
transform 1 0 3124 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1677622389
transform 1 0 3140 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_251
timestamp 1677622389
transform -1 0 3152 0 1 1970
box -8 -3 46 105
use FILL  FILL_6878
timestamp 1677622389
transform 1 0 3152 0 1 1970
box -8 -3 16 105
use FILL  FILL_6879
timestamp 1677622389
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6884
timestamp 1677622389
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6886
timestamp 1677622389
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6888
timestamp 1677622389
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_41
timestamp 1677622389
transform -1 0 3224 0 1 1970
box -8 -3 40 105
use FILL  FILL_6889
timestamp 1677622389
transform 1 0 3224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6890
timestamp 1677622389
transform 1 0 3232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6891
timestamp 1677622389
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_42
timestamp 1677622389
transform -1 0 3280 0 1 1970
box -8 -3 40 105
use FILL  FILL_6892
timestamp 1677622389
transform 1 0 3280 0 1 1970
box -8 -3 16 105
use FILL  FILL_6893
timestamp 1677622389
transform 1 0 3288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6894
timestamp 1677622389
transform 1 0 3296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6895
timestamp 1677622389
transform 1 0 3304 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1677622389
transform -1 0 3344 0 1 1970
box -8 -3 40 105
use FILL  FILL_6896
timestamp 1677622389
transform 1 0 3344 0 1 1970
box -8 -3 16 105
use FILL  FILL_6907
timestamp 1677622389
transform 1 0 3352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6908
timestamp 1677622389
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6909
timestamp 1677622389
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6910
timestamp 1677622389
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6911
timestamp 1677622389
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6912
timestamp 1677622389
transform 1 0 3392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6915
timestamp 1677622389
transform 1 0 3400 0 1 1970
box -8 -3 16 105
use FILL  FILL_6917
timestamp 1677622389
transform 1 0 3408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6919
timestamp 1677622389
transform 1 0 3416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6920
timestamp 1677622389
transform 1 0 3424 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_46
timestamp 1677622389
transform -1 0 3464 0 1 1970
box -8 -3 40 105
use FILL  FILL_6921
timestamp 1677622389
transform 1 0 3464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6925
timestamp 1677622389
transform 1 0 3472 0 1 1970
box -8 -3 16 105
use FILL  FILL_6927
timestamp 1677622389
transform 1 0 3480 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_431
timestamp 1677622389
transform -1 0 3504 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_380
timestamp 1677622389
transform -1 0 3600 0 1 1970
box -8 -3 104 105
use FILL  FILL_6928
timestamp 1677622389
transform 1 0 3600 0 1 1970
box -8 -3 16 105
use FILL  FILL_6929
timestamp 1677622389
transform 1 0 3608 0 1 1970
box -8 -3 16 105
use FILL  FILL_6930
timestamp 1677622389
transform 1 0 3616 0 1 1970
box -8 -3 16 105
use FILL  FILL_6931
timestamp 1677622389
transform 1 0 3624 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5059
timestamp 1677622389
transform 1 0 3644 0 1 1975
box -3 -3 3 3
use FILL  FILL_6932
timestamp 1677622389
transform 1 0 3632 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5060
timestamp 1677622389
transform 1 0 3676 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_252
timestamp 1677622389
transform -1 0 3680 0 1 1970
box -8 -3 46 105
use FILL  FILL_6933
timestamp 1677622389
transform 1 0 3680 0 1 1970
box -8 -3 16 105
use FILL  FILL_6934
timestamp 1677622389
transform 1 0 3688 0 1 1970
box -8 -3 16 105
use FILL  FILL_6935
timestamp 1677622389
transform 1 0 3696 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5061
timestamp 1677622389
transform 1 0 3716 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_381
timestamp 1677622389
transform 1 0 3704 0 1 1970
box -8 -3 104 105
use FILL  FILL_6936
timestamp 1677622389
transform 1 0 3800 0 1 1970
box -8 -3 16 105
use FILL  FILL_6956
timestamp 1677622389
transform 1 0 3808 0 1 1970
box -8 -3 16 105
use FILL  FILL_6958
timestamp 1677622389
transform 1 0 3816 0 1 1970
box -8 -3 16 105
use FILL  FILL_6960
timestamp 1677622389
transform 1 0 3824 0 1 1970
box -8 -3 16 105
use FILL  FILL_6962
timestamp 1677622389
transform 1 0 3832 0 1 1970
box -8 -3 16 105
use FILL  FILL_6963
timestamp 1677622389
transform 1 0 3840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6964
timestamp 1677622389
transform 1 0 3848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6965
timestamp 1677622389
transform 1 0 3856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6966
timestamp 1677622389
transform 1 0 3864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6967
timestamp 1677622389
transform 1 0 3872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6969
timestamp 1677622389
transform 1 0 3880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6971
timestamp 1677622389
transform 1 0 3888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6973
timestamp 1677622389
transform 1 0 3896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6975
timestamp 1677622389
transform 1 0 3904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6976
timestamp 1677622389
transform 1 0 3912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6977
timestamp 1677622389
transform 1 0 3920 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5062
timestamp 1677622389
transform 1 0 3940 0 1 1975
box -3 -3 3 3
use FILL  FILL_6978
timestamp 1677622389
transform 1 0 3928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6979
timestamp 1677622389
transform 1 0 3936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6980
timestamp 1677622389
transform 1 0 3944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6981
timestamp 1677622389
transform 1 0 3952 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5063
timestamp 1677622389
transform 1 0 3972 0 1 1975
box -3 -3 3 3
use FILL  FILL_6982
timestamp 1677622389
transform 1 0 3960 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_382
timestamp 1677622389
transform -1 0 4064 0 1 1970
box -8 -3 104 105
use AOI22X1  AOI22X1_269
timestamp 1677622389
transform -1 0 4104 0 1 1970
box -8 -3 46 105
use FILL  FILL_6983
timestamp 1677622389
transform 1 0 4104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6984
timestamp 1677622389
transform 1 0 4112 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_433
timestamp 1677622389
transform 1 0 4120 0 1 1970
box -9 -3 26 105
use FILL  FILL_6985
timestamp 1677622389
transform 1 0 4136 0 1 1970
box -8 -3 16 105
use FILL  FILL_6986
timestamp 1677622389
transform 1 0 4144 0 1 1970
box -8 -3 16 105
use FILL  FILL_6987
timestamp 1677622389
transform 1 0 4152 0 1 1970
box -8 -3 16 105
use FILL  FILL_6988
timestamp 1677622389
transform 1 0 4160 0 1 1970
box -8 -3 16 105
use FILL  FILL_6989
timestamp 1677622389
transform 1 0 4168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6990
timestamp 1677622389
transform 1 0 4176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6991
timestamp 1677622389
transform 1 0 4184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6992
timestamp 1677622389
transform 1 0 4192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6993
timestamp 1677622389
transform 1 0 4200 0 1 1970
box -8 -3 16 105
use FILL  FILL_6994
timestamp 1677622389
transform 1 0 4208 0 1 1970
box -8 -3 16 105
use FILL  FILL_6995
timestamp 1677622389
transform 1 0 4216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6996
timestamp 1677622389
transform 1 0 4224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6997
timestamp 1677622389
transform 1 0 4232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6998
timestamp 1677622389
transform 1 0 4240 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_383
timestamp 1677622389
transform -1 0 4344 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5064
timestamp 1677622389
transform 1 0 4428 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_384
timestamp 1677622389
transform -1 0 4440 0 1 1970
box -8 -3 104 105
use AND2X2  AND2X2_26
timestamp 1677622389
transform -1 0 4472 0 1 1970
box -8 -3 40 105
use INVX2  INVX2_434
timestamp 1677622389
transform 1 0 4472 0 1 1970
box -9 -3 26 105
use AND2X2  AND2X2_27
timestamp 1677622389
transform 1 0 4488 0 1 1970
box -8 -3 40 105
use FILL  FILL_6999
timestamp 1677622389
transform 1 0 4520 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_388
timestamp 1677622389
transform 1 0 4528 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_439
timestamp 1677622389
transform -1 0 4640 0 1 1970
box -9 -3 26 105
use FILL  FILL_7016
timestamp 1677622389
transform 1 0 4640 0 1 1970
box -8 -3 16 105
use FILL  FILL_7017
timestamp 1677622389
transform 1 0 4648 0 1 1970
box -8 -3 16 105
use FILL  FILL_7022
timestamp 1677622389
transform 1 0 4656 0 1 1970
box -8 -3 16 105
use FILL  FILL_7024
timestamp 1677622389
transform 1 0 4664 0 1 1970
box -8 -3 16 105
use FILL  FILL_7025
timestamp 1677622389
transform 1 0 4672 0 1 1970
box -8 -3 16 105
use FILL  FILL_7026
timestamp 1677622389
transform 1 0 4680 0 1 1970
box -8 -3 16 105
use FILL  FILL_7027
timestamp 1677622389
transform 1 0 4688 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_389
timestamp 1677622389
transform 1 0 4696 0 1 1970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_55
timestamp 1677622389
transform 1 0 4819 0 1 1970
box -10 -3 10 3
use M2_M1  M2_M1_5705
timestamp 1677622389
transform 1 0 92 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1677622389
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1677622389
transform 1 0 172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1677622389
transform 1 0 180 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5151
timestamp 1677622389
transform 1 0 140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1677622389
transform 1 0 180 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1677622389
transform 1 0 172 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5706
timestamp 1677622389
transform 1 0 212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1677622389
transform 1 0 220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1677622389
transform 1 0 236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1677622389
transform 1 0 244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1677622389
transform 1 0 204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1677622389
transform 1 0 228 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5184
timestamp 1677622389
transform 1 0 220 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1677622389
transform 1 0 268 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5793
timestamp 1677622389
transform 1 0 260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1677622389
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5087
timestamp 1677622389
transform 1 0 300 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5710
timestamp 1677622389
transform 1 0 292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1677622389
transform 1 0 300 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5088
timestamp 1677622389
transform 1 0 332 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5795
timestamp 1677622389
transform 1 0 332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1677622389
transform 1 0 340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1677622389
transform 1 0 412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1677622389
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1677622389
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1677622389
transform 1 0 508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5185
timestamp 1677622389
transform 1 0 500 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1677622389
transform 1 0 484 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1677622389
transform 1 0 556 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5799
timestamp 1677622389
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1677622389
transform 1 0 580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1677622389
transform 1 0 572 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5212
timestamp 1677622389
transform 1 0 572 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1677622389
transform 1 0 604 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5801
timestamp 1677622389
transform 1 0 628 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5186
timestamp 1677622389
transform 1 0 628 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5702
timestamp 1677622389
transform 1 0 644 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5123
timestamp 1677622389
transform 1 0 644 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1677622389
transform 1 0 668 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5715
timestamp 1677622389
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5091
timestamp 1677622389
transform 1 0 684 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5716
timestamp 1677622389
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1677622389
transform 1 0 724 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5070
timestamp 1677622389
transform 1 0 740 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5717
timestamp 1677622389
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1677622389
transform 1 0 828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1677622389
transform 1 0 780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1677622389
transform 1 0 828 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5153
timestamp 1677622389
transform 1 0 780 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5805
timestamp 1677622389
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1677622389
transform 1 0 844 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5154
timestamp 1677622389
transform 1 0 836 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1677622389
transform 1 0 828 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1677622389
transform 1 0 836 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1677622389
transform 1 0 860 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5719
timestamp 1677622389
transform 1 0 884 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5092
timestamp 1677622389
transform 1 0 908 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5807
timestamp 1677622389
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5214
timestamp 1677622389
transform 1 0 892 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1677622389
transform 1 0 940 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1677622389
transform 1 0 932 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5720
timestamp 1677622389
transform 1 0 932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1677622389
transform 1 0 964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1677622389
transform 1 0 940 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1677622389
transform 1 0 956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1677622389
transform 1 0 980 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5124
timestamp 1677622389
transform 1 0 980 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1677622389
transform 1 0 1004 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1677622389
transform 1 0 1060 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1677622389
transform 1 0 1132 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1677622389
transform 1 0 1164 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5810
timestamp 1677622389
transform 1 0 1156 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5155
timestamp 1677622389
transform 1 0 1156 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1677622389
transform 1 0 1172 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5722
timestamp 1677622389
transform 1 0 1172 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5073
timestamp 1677622389
transform 1 0 1260 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5811
timestamp 1677622389
transform 1 0 1196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1677622389
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5156
timestamp 1677622389
transform 1 0 1196 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1677622389
transform 1 0 1172 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5813
timestamp 1677622389
transform 1 0 1284 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5187
timestamp 1677622389
transform 1 0 1292 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1677622389
transform 1 0 1316 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5814
timestamp 1677622389
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5157
timestamp 1677622389
transform 1 0 1308 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5893
timestamp 1677622389
transform 1 0 1324 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5188
timestamp 1677622389
transform 1 0 1308 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1677622389
transform 1 0 1340 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5723
timestamp 1677622389
transform 1 0 1372 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5136
timestamp 1677622389
transform 1 0 1372 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1677622389
transform 1 0 1420 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1677622389
transform 1 0 1460 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5724
timestamp 1677622389
transform 1 0 1460 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5137
timestamp 1677622389
transform 1 0 1388 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5815
timestamp 1677622389
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1677622389
transform 1 0 1492 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5189
timestamp 1677622389
transform 1 0 1492 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1677622389
transform 1 0 1516 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5725
timestamp 1677622389
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5205
timestamp 1677622389
transform 1 0 1508 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1677622389
transform 1 0 1532 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5817
timestamp 1677622389
transform 1 0 1532 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5215
timestamp 1677622389
transform 1 0 1524 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1677622389
transform 1 0 1548 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1677622389
transform 1 0 1588 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5818
timestamp 1677622389
transform 1 0 1612 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1677622389
transform 1 0 1644 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5138
timestamp 1677622389
transform 1 0 1644 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5727
timestamp 1677622389
transform 1 0 1700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1677622389
transform 1 0 1716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1677622389
transform 1 0 1804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1677622389
transform 1 0 1820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1677622389
transform 1 0 1828 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5139
timestamp 1677622389
transform 1 0 1844 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5729
timestamp 1677622389
transform 1 0 1868 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5140
timestamp 1677622389
transform 1 0 1868 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1677622389
transform 1 0 1884 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5730
timestamp 1677622389
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1677622389
transform 1 0 1908 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5141
timestamp 1677622389
transform 1 0 1956 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5823
timestamp 1677622389
transform 1 0 1964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1677622389
transform 1 0 1972 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5216
timestamp 1677622389
transform 1 0 1964 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1677622389
transform 1 0 2020 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5825
timestamp 1677622389
transform 1 0 2036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1677622389
transform 1 0 2060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1677622389
transform 1 0 2052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1677622389
transform 1 0 2052 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5074
timestamp 1677622389
transform 1 0 2076 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5895
timestamp 1677622389
transform 1 0 2068 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5192
timestamp 1677622389
transform 1 0 2084 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1677622389
transform 1 0 2124 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5732
timestamp 1677622389
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5100
timestamp 1677622389
transform 1 0 2244 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5733
timestamp 1677622389
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5101
timestamp 1677622389
transform 1 0 2292 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5734
timestamp 1677622389
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1677622389
transform 1 0 2268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1677622389
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1677622389
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5159
timestamp 1677622389
transform 1 0 2268 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1677622389
transform 1 0 2308 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1677622389
transform 1 0 2332 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1677622389
transform 1 0 2372 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5735
timestamp 1677622389
transform 1 0 2388 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5162
timestamp 1677622389
transform 1 0 2380 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5736
timestamp 1677622389
transform 1 0 2404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1677622389
transform 1 0 2412 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5163
timestamp 1677622389
transform 1 0 2412 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1677622389
transform 1 0 2436 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5737
timestamp 1677622389
transform 1 0 2508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1677622389
transform 1 0 2460 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5164
timestamp 1677622389
transform 1 0 2460 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1677622389
transform 1 0 2468 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1677622389
transform 1 0 2580 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5738
timestamp 1677622389
transform 1 0 2572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1677622389
transform 1 0 2588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1677622389
transform 1 0 2564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1677622389
transform 1 0 2580 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5206
timestamp 1677622389
transform 1 0 2556 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1677622389
transform 1 0 2588 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1677622389
transform 1 0 2564 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1677622389
transform 1 0 2604 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5740
timestamp 1677622389
transform 1 0 2604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1677622389
transform 1 0 2620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1677622389
transform 1 0 2636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1677622389
transform 1 0 2676 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5165
timestamp 1677622389
transform 1 0 2676 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5741
timestamp 1677622389
transform 1 0 2692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1677622389
transform 1 0 2716 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5143
timestamp 1677622389
transform 1 0 2764 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5704
timestamp 1677622389
transform 1 0 2780 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1677622389
transform 1 0 2772 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5166
timestamp 1677622389
transform 1 0 2716 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5839
timestamp 1677622389
transform 1 0 2796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1677622389
transform 1 0 2836 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5144
timestamp 1677622389
transform 1 0 2844 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1677622389
transform 1 0 2836 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5743
timestamp 1677622389
transform 1 0 2868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1677622389
transform 1 0 2860 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5145
timestamp 1677622389
transform 1 0 2868 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5896
timestamp 1677622389
transform 1 0 2868 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1677622389
transform 1 0 2892 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1677622389
transform 1 0 2916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1677622389
transform 1 0 2948 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5075
timestamp 1677622389
transform 1 0 3004 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1677622389
transform 1 0 3036 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1677622389
transform 1 0 3012 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5745
timestamp 1677622389
transform 1 0 3036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1677622389
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1677622389
transform 1 0 3012 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5107
timestamp 1677622389
transform 1 0 3052 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1677622389
transform 1 0 3076 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5746
timestamp 1677622389
transform 1 0 3076 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1677622389
transform 1 0 3124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1677622389
transform 1 0 3156 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5219
timestamp 1677622389
transform 1 0 3108 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5898
timestamp 1677622389
transform 1 0 3164 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5078
timestamp 1677622389
transform 1 0 3188 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1677622389
transform 1 0 3188 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1677622389
transform 1 0 3204 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5846
timestamp 1677622389
transform 1 0 3228 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5167
timestamp 1677622389
transform 1 0 3228 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5902
timestamp 1677622389
transform 1 0 3220 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1677622389
transform 1 0 3244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1677622389
transform 1 0 3252 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1677622389
transform 1 0 3284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1677622389
transform 1 0 3292 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5220
timestamp 1677622389
transform 1 0 3276 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5749
timestamp 1677622389
transform 1 0 3308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1677622389
transform 1 0 3316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1677622389
transform 1 0 3332 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5168
timestamp 1677622389
transform 1 0 3332 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5900
timestamp 1677622389
transform 1 0 3340 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5108
timestamp 1677622389
transform 1 0 3388 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5850
timestamp 1677622389
transform 1 0 3380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1677622389
transform 1 0 3372 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5208
timestamp 1677622389
transform 1 0 3372 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5750
timestamp 1677622389
transform 1 0 3412 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5109
timestamp 1677622389
transform 1 0 3428 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5851
timestamp 1677622389
transform 1 0 3428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1677622389
transform 1 0 3420 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5209
timestamp 1677622389
transform 1 0 3420 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1677622389
transform 1 0 3476 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1677622389
transform 1 0 3484 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5751
timestamp 1677622389
transform 1 0 3492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1677622389
transform 1 0 3476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1677622389
transform 1 0 3484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1677622389
transform 1 0 3500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1677622389
transform 1 0 3516 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5193
timestamp 1677622389
transform 1 0 3484 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1677622389
transform 1 0 3516 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1677622389
transform 1 0 3556 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5752
timestamp 1677622389
transform 1 0 3564 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5111
timestamp 1677622389
transform 1 0 3580 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5753
timestamp 1677622389
transform 1 0 3580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1677622389
transform 1 0 3604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1677622389
transform 1 0 3628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1677622389
transform 1 0 3644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1677622389
transform 1 0 3620 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5146
timestamp 1677622389
transform 1 0 3644 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1677622389
transform 1 0 3716 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5756
timestamp 1677622389
transform 1 0 3684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1677622389
transform 1 0 3700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1677622389
transform 1 0 3716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1677622389
transform 1 0 3724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1677622389
transform 1 0 3692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1677622389
transform 1 0 3708 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5169
timestamp 1677622389
transform 1 0 3692 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5760
timestamp 1677622389
transform 1 0 3740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1677622389
transform 1 0 3732 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5195
timestamp 1677622389
transform 1 0 3732 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5861
timestamp 1677622389
transform 1 0 3780 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5147
timestamp 1677622389
transform 1 0 3788 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5862
timestamp 1677622389
transform 1 0 3796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1677622389
transform 1 0 3820 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5113
timestamp 1677622389
transform 1 0 3844 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5762
timestamp 1677622389
transform 1 0 3844 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5132
timestamp 1677622389
transform 1 0 3868 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5863
timestamp 1677622389
transform 1 0 3836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1677622389
transform 1 0 3852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1677622389
transform 1 0 3868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1677622389
transform 1 0 3876 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5170
timestamp 1677622389
transform 1 0 3876 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1677622389
transform 1 0 3868 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1677622389
transform 1 0 3852 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1677622389
transform 1 0 3900 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1677622389
transform 1 0 3916 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1677622389
transform 1 0 3948 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5763
timestamp 1677622389
transform 1 0 3900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1677622389
transform 1 0 3908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1677622389
transform 1 0 3924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1677622389
transform 1 0 3940 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5171
timestamp 1677622389
transform 1 0 3900 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5867
timestamp 1677622389
transform 1 0 3916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1677622389
transform 1 0 3932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1677622389
transform 1 0 3948 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5172
timestamp 1677622389
transform 1 0 3932 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1677622389
transform 1 0 3948 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5767
timestamp 1677622389
transform 1 0 3964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1677622389
transform 1 0 4044 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5133
timestamp 1677622389
transform 1 0 4068 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1677622389
transform 1 0 4092 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1677622389
transform 1 0 4044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1677622389
transform 1 0 4148 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1677622389
transform 1 0 4212 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1677622389
transform 1 0 4140 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5769
timestamp 1677622389
transform 1 0 4212 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5116
timestamp 1677622389
transform 1 0 4284 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1677622389
transform 1 0 4308 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5770
timestamp 1677622389
transform 1 0 4308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1677622389
transform 1 0 4092 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1677622389
transform 1 0 4124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1677622389
transform 1 0 4132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1677622389
transform 1 0 4172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1677622389
transform 1 0 4228 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5197
timestamp 1677622389
transform 1 0 4044 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1677622389
transform 1 0 4164 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1677622389
transform 1 0 4172 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1677622389
transform 1 0 4244 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5875
timestamp 1677622389
transform 1 0 4260 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5175
timestamp 1677622389
transform 1 0 4260 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5876
timestamp 1677622389
transform 1 0 4340 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5176
timestamp 1677622389
transform 1 0 4340 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5771
timestamp 1677622389
transform 1 0 4348 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5082
timestamp 1677622389
transform 1 0 4364 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1677622389
transform 1 0 4396 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5772
timestamp 1677622389
transform 1 0 4364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1677622389
transform 1 0 4380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1677622389
transform 1 0 4396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1677622389
transform 1 0 4372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1677622389
transform 1 0 4388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1677622389
transform 1 0 4396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1677622389
transform 1 0 4420 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5177
timestamp 1677622389
transform 1 0 4364 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1677622389
transform 1 0 4388 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1677622389
transform 1 0 4436 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5775
timestamp 1677622389
transform 1 0 4436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1677622389
transform 1 0 4436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5179
timestamp 1677622389
transform 1 0 4436 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5776
timestamp 1677622389
transform 1 0 4460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1677622389
transform 1 0 4460 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5119
timestamp 1677622389
transform 1 0 4476 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5777
timestamp 1677622389
transform 1 0 4492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1677622389
transform 1 0 4484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1677622389
transform 1 0 4500 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5180
timestamp 1677622389
transform 1 0 4484 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5778
timestamp 1677622389
transform 1 0 4516 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5083
timestamp 1677622389
transform 1 0 4524 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5779
timestamp 1677622389
transform 1 0 4524 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5068
timestamp 1677622389
transform 1 0 4580 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1677622389
transform 1 0 4588 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5780
timestamp 1677622389
transform 1 0 4564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1677622389
transform 1 0 4580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1677622389
transform 1 0 4556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1677622389
transform 1 0 4572 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1677622389
transform 1 0 4588 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5069
timestamp 1677622389
transform 1 0 4604 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1677622389
transform 1 0 4644 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5782
timestamp 1677622389
transform 1 0 4604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1677622389
transform 1 0 4628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1677622389
transform 1 0 4644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1677622389
transform 1 0 4620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1677622389
transform 1 0 4636 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5181
timestamp 1677622389
transform 1 0 4644 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1677622389
transform 1 0 4620 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5785
timestamp 1677622389
transform 1 0 4660 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5120
timestamp 1677622389
transform 1 0 4676 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1677622389
transform 1 0 4708 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5786
timestamp 1677622389
transform 1 0 4676 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5150
timestamp 1677622389
transform 1 0 4676 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5890
timestamp 1677622389
transform 1 0 4700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1677622389
transform 1 0 4756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1677622389
transform 1 0 4764 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5182
timestamp 1677622389
transform 1 0 4700 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1677622389
transform 1 0 4764 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5787
timestamp 1677622389
transform 1 0 4788 0 1 1935
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_56
timestamp 1677622389
transform 1 0 24 0 1 1870
box -10 -3 10 3
use FILL  FILL_6510
timestamp 1677622389
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_364
timestamp 1677622389
transform 1 0 80 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6514
timestamp 1677622389
transform 1 0 176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6515
timestamp 1677622389
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_415
timestamp 1677622389
transform -1 0 208 0 -1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_255
timestamp 1677622389
transform -1 0 248 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6516
timestamp 1677622389
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6518
timestamp 1677622389
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6521
timestamp 1677622389
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_72
timestamp 1677622389
transform 1 0 272 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6522
timestamp 1677622389
transform 1 0 296 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_73
timestamp 1677622389
transform -1 0 328 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6523
timestamp 1677622389
transform 1 0 328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6524
timestamp 1677622389
transform 1 0 336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6525
timestamp 1677622389
transform 1 0 344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6526
timestamp 1677622389
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_416
timestamp 1677622389
transform -1 0 376 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6527
timestamp 1677622389
transform 1 0 376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6528
timestamp 1677622389
transform 1 0 384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6529
timestamp 1677622389
transform 1 0 392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6530
timestamp 1677622389
transform 1 0 400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6531
timestamp 1677622389
transform 1 0 408 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_367
timestamp 1677622389
transform 1 0 416 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6532
timestamp 1677622389
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6533
timestamp 1677622389
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6534
timestamp 1677622389
transform 1 0 528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6535
timestamp 1677622389
transform 1 0 536 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_74
timestamp 1677622389
transform 1 0 544 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6536
timestamp 1677622389
transform 1 0 568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6538
timestamp 1677622389
transform 1 0 576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6540
timestamp 1677622389
transform 1 0 584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6546
timestamp 1677622389
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6547
timestamp 1677622389
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_21
timestamp 1677622389
transform -1 0 640 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6548
timestamp 1677622389
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6549
timestamp 1677622389
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6550
timestamp 1677622389
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6551
timestamp 1677622389
transform 1 0 664 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_61
timestamp 1677622389
transform 1 0 672 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6552
timestamp 1677622389
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6554
timestamp 1677622389
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6564
timestamp 1677622389
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5221
timestamp 1677622389
transform 1 0 732 0 1 1875
box -3 -3 3 3
use FILL  FILL_6565
timestamp 1677622389
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_368
timestamp 1677622389
transform 1 0 728 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5222
timestamp 1677622389
transform 1 0 844 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_417
timestamp 1677622389
transform 1 0 824 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_418
timestamp 1677622389
transform -1 0 856 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6566
timestamp 1677622389
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6568
timestamp 1677622389
transform 1 0 864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6570
timestamp 1677622389
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6572
timestamp 1677622389
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6574
timestamp 1677622389
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6575
timestamp 1677622389
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6576
timestamp 1677622389
transform 1 0 904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6577
timestamp 1677622389
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_259
timestamp 1677622389
transform 1 0 920 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6584
timestamp 1677622389
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6586
timestamp 1677622389
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6588
timestamp 1677622389
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5223
timestamp 1677622389
transform 1 0 996 0 1 1875
box -3 -3 3 3
use FILL  FILL_6590
timestamp 1677622389
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6592
timestamp 1677622389
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6594
timestamp 1677622389
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6596
timestamp 1677622389
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6598
timestamp 1677622389
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6600
timestamp 1677622389
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6602
timestamp 1677622389
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6603
timestamp 1677622389
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6604
timestamp 1677622389
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6605
timestamp 1677622389
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6607
timestamp 1677622389
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6609
timestamp 1677622389
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6611
timestamp 1677622389
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6613
timestamp 1677622389
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6615
timestamp 1677622389
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6617
timestamp 1677622389
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_419
timestamp 1677622389
transform 1 0 1112 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6621
timestamp 1677622389
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6623
timestamp 1677622389
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6625
timestamp 1677622389
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6627
timestamp 1677622389
transform 1 0 1152 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_369
timestamp 1677622389
transform 1 0 1160 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6639
timestamp 1677622389
transform 1 0 1256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6640
timestamp 1677622389
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6641
timestamp 1677622389
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6643
timestamp 1677622389
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6650
timestamp 1677622389
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_22
timestamp 1677622389
transform -1 0 1328 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6651
timestamp 1677622389
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6653
timestamp 1677622389
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6669
timestamp 1677622389
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6670
timestamp 1677622389
transform 1 0 1352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6671
timestamp 1677622389
transform 1 0 1360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6672
timestamp 1677622389
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_370
timestamp 1677622389
transform -1 0 1472 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6673
timestamp 1677622389
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6674
timestamp 1677622389
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6675
timestamp 1677622389
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_75
timestamp 1677622389
transform 1 0 1496 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6676
timestamp 1677622389
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6680
timestamp 1677622389
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_77
timestamp 1677622389
transform -1 0 1560 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6681
timestamp 1677622389
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6682
timestamp 1677622389
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6684
timestamp 1677622389
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6686
timestamp 1677622389
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6688
timestamp 1677622389
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6691
timestamp 1677622389
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_79
timestamp 1677622389
transform 1 0 1608 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6692
timestamp 1677622389
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6694
timestamp 1677622389
transform 1 0 1640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6696
timestamp 1677622389
transform 1 0 1648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6699
timestamp 1677622389
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6700
timestamp 1677622389
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6701
timestamp 1677622389
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6702
timestamp 1677622389
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6703
timestamp 1677622389
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6704
timestamp 1677622389
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6705
timestamp 1677622389
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6706
timestamp 1677622389
transform 1 0 1712 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_420
timestamp 1677622389
transform 1 0 1720 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6707
timestamp 1677622389
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6708
timestamp 1677622389
transform 1 0 1744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6709
timestamp 1677622389
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6710
timestamp 1677622389
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6711
timestamp 1677622389
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6712
timestamp 1677622389
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6713
timestamp 1677622389
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6715
timestamp 1677622389
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_421
timestamp 1677622389
transform 1 0 1800 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6719
timestamp 1677622389
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6721
timestamp 1677622389
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_81
timestamp 1677622389
transform 1 0 1832 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6733
timestamp 1677622389
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6734
timestamp 1677622389
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_372
timestamp 1677622389
transform 1 0 1872 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6735
timestamp 1677622389
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6737
timestamp 1677622389
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6739
timestamp 1677622389
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6741
timestamp 1677622389
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6743
timestamp 1677622389
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6745
timestamp 1677622389
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_24
timestamp 1677622389
transform -1 0 2048 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6746
timestamp 1677622389
transform 1 0 2048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6747
timestamp 1677622389
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6748
timestamp 1677622389
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_423
timestamp 1677622389
transform -1 0 2088 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6749
timestamp 1677622389
transform 1 0 2088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6750
timestamp 1677622389
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6751
timestamp 1677622389
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6753
timestamp 1677622389
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6755
timestamp 1677622389
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6757
timestamp 1677622389
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6760
timestamp 1677622389
transform 1 0 2136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6761
timestamp 1677622389
transform 1 0 2144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6762
timestamp 1677622389
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6763
timestamp 1677622389
transform 1 0 2160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6764
timestamp 1677622389
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6765
timestamp 1677622389
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6766
timestamp 1677622389
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6768
timestamp 1677622389
transform 1 0 2192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6770
timestamp 1677622389
transform 1 0 2200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6772
timestamp 1677622389
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6774
timestamp 1677622389
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6776
timestamp 1677622389
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6778
timestamp 1677622389
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_424
timestamp 1677622389
transform 1 0 2240 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6782
timestamp 1677622389
transform 1 0 2256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6792
timestamp 1677622389
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_374
timestamp 1677622389
transform -1 0 2368 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6793
timestamp 1677622389
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6795
timestamp 1677622389
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_426
timestamp 1677622389
transform 1 0 2384 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6807
timestamp 1677622389
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6808
timestamp 1677622389
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6809
timestamp 1677622389
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_375
timestamp 1677622389
transform -1 0 2520 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6810
timestamp 1677622389
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6812
timestamp 1677622389
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6814
timestamp 1677622389
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6816
timestamp 1677622389
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6818
timestamp 1677622389
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_265
timestamp 1677622389
transform 1 0 2560 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6823
timestamp 1677622389
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6824
timestamp 1677622389
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6825
timestamp 1677622389
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6826
timestamp 1677622389
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6828
timestamp 1677622389
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6830
timestamp 1677622389
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_427
timestamp 1677622389
transform 1 0 2648 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6835
timestamp 1677622389
transform 1 0 2664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6836
timestamp 1677622389
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_377
timestamp 1677622389
transform 1 0 2680 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6837
timestamp 1677622389
transform 1 0 2776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6838
timestamp 1677622389
transform 1 0 2784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6839
timestamp 1677622389
transform 1 0 2792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6840
timestamp 1677622389
transform 1 0 2800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6842
timestamp 1677622389
transform 1 0 2808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6844
timestamp 1677622389
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6846
timestamp 1677622389
transform 1 0 2824 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_64
timestamp 1677622389
transform 1 0 2832 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6851
timestamp 1677622389
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6853
timestamp 1677622389
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6855
timestamp 1677622389
transform 1 0 2872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6859
timestamp 1677622389
transform 1 0 2880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6860
timestamp 1677622389
transform 1 0 2888 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_126
timestamp 1677622389
transform -1 0 2928 0 -1 1970
box -8 -3 34 105
use FILL  FILL_6861
timestamp 1677622389
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6863
timestamp 1677622389
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6880
timestamp 1677622389
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_378
timestamp 1677622389
transform -1 0 3048 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6881
timestamp 1677622389
transform 1 0 3048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6882
timestamp 1677622389
transform 1 0 3056 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_379
timestamp 1677622389
transform 1 0 3064 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6883
timestamp 1677622389
transform 1 0 3160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6885
timestamp 1677622389
transform 1 0 3168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6887
timestamp 1677622389
transform 1 0 3176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6897
timestamp 1677622389
transform 1 0 3184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6898
timestamp 1677622389
transform 1 0 3192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6899
timestamp 1677622389
transform 1 0 3200 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5224
timestamp 1677622389
transform 1 0 3220 0 1 1875
box -3 -3 3 3
use NAND3X1  NAND3X1_44
timestamp 1677622389
transform -1 0 3240 0 -1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5225
timestamp 1677622389
transform 1 0 3252 0 1 1875
box -3 -3 3 3
use FILL  FILL_6900
timestamp 1677622389
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6901
timestamp 1677622389
transform 1 0 3248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6902
timestamp 1677622389
transform 1 0 3256 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5226
timestamp 1677622389
transform 1 0 3292 0 1 1875
box -3 -3 3 3
use BUFX2  BUFX2_82
timestamp 1677622389
transform 1 0 3264 0 -1 1970
box -5 -3 28 105
use INVX2  INVX2_429
timestamp 1677622389
transform 1 0 3288 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6903
timestamp 1677622389
transform 1 0 3304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6904
timestamp 1677622389
transform 1 0 3312 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_430
timestamp 1677622389
transform 1 0 3320 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6905
timestamp 1677622389
transform 1 0 3336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6906
timestamp 1677622389
transform 1 0 3344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6913
timestamp 1677622389
transform 1 0 3352 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_45
timestamp 1677622389
transform -1 0 3392 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6914
timestamp 1677622389
transform 1 0 3392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6916
timestamp 1677622389
transform 1 0 3400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6918
timestamp 1677622389
transform 1 0 3408 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1677622389
transform 1 0 3416 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6922
timestamp 1677622389
transform 1 0 3448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6923
timestamp 1677622389
transform 1 0 3456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6924
timestamp 1677622389
transform 1 0 3464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6926
timestamp 1677622389
transform 1 0 3472 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_266
timestamp 1677622389
transform 1 0 3480 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6937
timestamp 1677622389
transform 1 0 3520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6938
timestamp 1677622389
transform 1 0 3528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6939
timestamp 1677622389
transform 1 0 3536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6940
timestamp 1677622389
transform 1 0 3544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6941
timestamp 1677622389
transform 1 0 3552 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_432
timestamp 1677622389
transform 1 0 3560 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6942
timestamp 1677622389
transform 1 0 3576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6943
timestamp 1677622389
transform 1 0 3584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6944
timestamp 1677622389
transform 1 0 3592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6945
timestamp 1677622389
transform 1 0 3600 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_253
timestamp 1677622389
transform -1 0 3648 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6946
timestamp 1677622389
transform 1 0 3648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6947
timestamp 1677622389
transform 1 0 3656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6948
timestamp 1677622389
transform 1 0 3664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6949
timestamp 1677622389
transform 1 0 3672 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_254
timestamp 1677622389
transform 1 0 3680 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6950
timestamp 1677622389
transform 1 0 3720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6951
timestamp 1677622389
transform 1 0 3728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6952
timestamp 1677622389
transform 1 0 3736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6953
timestamp 1677622389
transform 1 0 3744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6954
timestamp 1677622389
transform 1 0 3752 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_267
timestamp 1677622389
transform -1 0 3800 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6955
timestamp 1677622389
transform 1 0 3800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6957
timestamp 1677622389
transform 1 0 3808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6959
timestamp 1677622389
transform 1 0 3816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6961
timestamp 1677622389
transform 1 0 3824 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_268
timestamp 1677622389
transform 1 0 3832 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6968
timestamp 1677622389
transform 1 0 3872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6970
timestamp 1677622389
transform 1 0 3880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6972
timestamp 1677622389
transform 1 0 3888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6974
timestamp 1677622389
transform 1 0 3896 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_255
timestamp 1677622389
transform 1 0 3904 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_435
timestamp 1677622389
transform -1 0 3960 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7000
timestamp 1677622389
transform 1 0 3960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7001
timestamp 1677622389
transform 1 0 3968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7002
timestamp 1677622389
transform 1 0 3976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7003
timestamp 1677622389
transform 1 0 3984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7004
timestamp 1677622389
transform 1 0 3992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7005
timestamp 1677622389
transform 1 0 4000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7006
timestamp 1677622389
transform 1 0 4008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7007
timestamp 1677622389
transform 1 0 4016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7008
timestamp 1677622389
transform 1 0 4024 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_385
timestamp 1677622389
transform 1 0 4032 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_386
timestamp 1677622389
transform -1 0 4224 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_387
timestamp 1677622389
transform -1 0 4320 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_436
timestamp 1677622389
transform -1 0 4336 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7009
timestamp 1677622389
transform 1 0 4336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7010
timestamp 1677622389
transform 1 0 4344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7011
timestamp 1677622389
transform 1 0 4352 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_256
timestamp 1677622389
transform -1 0 4400 0 -1 1970
box -8 -3 46 105
use AND2X2  AND2X2_28
timestamp 1677622389
transform -1 0 4432 0 -1 1970
box -8 -3 40 105
use FILL  FILL_7012
timestamp 1677622389
transform 1 0 4432 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_437
timestamp 1677622389
transform -1 0 4456 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7013
timestamp 1677622389
transform 1 0 4456 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1677622389
transform -1 0 4496 0 -1 1970
box -8 -3 40 105
use INVX2  INVX2_438
timestamp 1677622389
transform -1 0 4512 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7014
timestamp 1677622389
transform 1 0 4512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7015
timestamp 1677622389
transform 1 0 4520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7018
timestamp 1677622389
transform 1 0 4528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7019
timestamp 1677622389
transform 1 0 4536 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_257
timestamp 1677622389
transform -1 0 4584 0 -1 1970
box -8 -3 46 105
use FILL  FILL_7020
timestamp 1677622389
transform 1 0 4584 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_440
timestamp 1677622389
transform -1 0 4608 0 -1 1970
box -9 -3 26 105
use OAI22X1  OAI22X1_258
timestamp 1677622389
transform 1 0 4608 0 -1 1970
box -8 -3 46 105
use FILL  FILL_7021
timestamp 1677622389
transform 1 0 4648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7023
timestamp 1677622389
transform 1 0 4656 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_390
timestamp 1677622389
transform 1 0 4664 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_441
timestamp 1677622389
transform -1 0 4776 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7028
timestamp 1677622389
transform 1 0 4776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7029
timestamp 1677622389
transform 1 0 4784 0 -1 1970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_57
timestamp 1677622389
transform 1 0 4843 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_5331
timestamp 1677622389
transform 1 0 84 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1677622389
transform 1 0 164 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1677622389
transform 1 0 148 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1677622389
transform 1 0 188 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5918
timestamp 1677622389
transform 1 0 148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1677622389
transform 1 0 180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1677622389
transform 1 0 188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1677622389
transform 1 0 100 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5332
timestamp 1677622389
transform 1 0 220 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6031
timestamp 1677622389
transform 1 0 228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1677622389
transform 1 0 220 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5333
timestamp 1677622389
transform 1 0 236 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1677622389
transform 1 0 260 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1677622389
transform 1 0 292 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1677622389
transform 1 0 332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1677622389
transform 1 0 372 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5921
timestamp 1677622389
transform 1 0 268 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5310
timestamp 1677622389
transform 1 0 284 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5922
timestamp 1677622389
transform 1 0 332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1677622389
transform 1 0 364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1677622389
transform 1 0 372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1677622389
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1677622389
transform 1 0 372 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5354
timestamp 1677622389
transform 1 0 356 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1677622389
transform 1 0 420 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1677622389
transform 1 0 428 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6034
timestamp 1677622389
transform 1 0 420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1677622389
transform 1 0 452 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5257
timestamp 1677622389
transform 1 0 492 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1677622389
transform 1 0 476 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5926
timestamp 1677622389
transform 1 0 476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1677622389
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1677622389
transform 1 0 460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1677622389
transform 1 0 468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1677622389
transform 1 0 484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1677622389
transform 1 0 492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1677622389
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5355
timestamp 1677622389
transform 1 0 460 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1677622389
transform 1 0 468 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1677622389
transform 1 0 508 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1677622389
transform 1 0 548 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5928
timestamp 1677622389
transform 1 0 548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1677622389
transform 1 0 556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1677622389
transform 1 0 572 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5387
timestamp 1677622389
transform 1 0 572 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1677622389
transform 1 0 588 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5929
timestamp 1677622389
transform 1 0 588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1677622389
transform 1 0 604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1677622389
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5259
timestamp 1677622389
transform 1 0 644 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5932
timestamp 1677622389
transform 1 0 644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1677622389
transform 1 0 644 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1677622389
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5356
timestamp 1677622389
transform 1 0 644 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1677622389
transform 1 0 692 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5933
timestamp 1677622389
transform 1 0 676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1677622389
transform 1 0 692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1677622389
transform 1 0 684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1677622389
transform 1 0 708 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5238
timestamp 1677622389
transform 1 0 724 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6045
timestamp 1677622389
transform 1 0 716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5284
timestamp 1677622389
transform 1 0 732 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1677622389
transform 1 0 748 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5935
timestamp 1677622389
transform 1 0 748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1677622389
transform 1 0 756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1677622389
transform 1 0 764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1677622389
transform 1 0 820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1677622389
transform 1 0 836 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5312
timestamp 1677622389
transform 1 0 852 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6048
timestamp 1677622389
transform 1 0 852 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5313
timestamp 1677622389
transform 1 0 884 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6049
timestamp 1677622389
transform 1 0 900 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5388
timestamp 1677622389
transform 1 0 900 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5938
timestamp 1677622389
transform 1 0 980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1677622389
transform 1 0 996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1677622389
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5314
timestamp 1677622389
transform 1 0 1036 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1677622389
transform 1 0 1052 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5940
timestamp 1677622389
transform 1 0 1060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1677622389
transform 1 0 1052 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5227
timestamp 1677622389
transform 1 0 1092 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1677622389
transform 1 0 1132 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1677622389
transform 1 0 1100 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1677622389
transform 1 0 1156 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1677622389
transform 1 0 1076 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5941
timestamp 1677622389
transform 1 0 1116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1677622389
transform 1 0 1164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1677622389
transform 1 0 1084 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5389
timestamp 1677622389
transform 1 0 1084 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1677622389
transform 1 0 1188 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1677622389
transform 1 0 1244 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1677622389
transform 1 0 1252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1677622389
transform 1 0 1276 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5943
timestamp 1677622389
transform 1 0 1244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1677622389
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1677622389
transform 1 0 1268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1677622389
transform 1 0 1252 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5334
timestamp 1677622389
transform 1 0 1268 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1677622389
transform 1 0 1260 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6054
timestamp 1677622389
transform 1 0 1324 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5316
timestamp 1677622389
transform 1 0 1372 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5946
timestamp 1677622389
transform 1 0 1380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1677622389
transform 1 0 1388 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5229
timestamp 1677622389
transform 1 0 1420 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6056
timestamp 1677622389
transform 1 0 1412 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5264
timestamp 1677622389
transform 1 0 1428 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5947
timestamp 1677622389
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1677622389
transform 1 0 1468 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5317
timestamp 1677622389
transform 1 0 1476 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1677622389
transform 1 0 1532 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5949
timestamp 1677622389
transform 1 0 1532 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5357
timestamp 1677622389
transform 1 0 1524 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5950
timestamp 1677622389
transform 1 0 1548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1677622389
transform 1 0 1564 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5231
timestamp 1677622389
transform 1 0 1596 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1677622389
transform 1 0 1620 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5951
timestamp 1677622389
transform 1 0 1620 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5335
timestamp 1677622389
transform 1 0 1628 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5952
timestamp 1677622389
transform 1 0 1644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1677622389
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5391
timestamp 1677622389
transform 1 0 1644 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6059
timestamp 1677622389
transform 1 0 1668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5239
timestamp 1677622389
transform 1 0 1724 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5953
timestamp 1677622389
transform 1 0 1716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1677622389
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1677622389
transform 1 0 1708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1677622389
transform 1 0 1724 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5358
timestamp 1677622389
transform 1 0 1700 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1677622389
transform 1 0 1732 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1677622389
transform 1 0 1724 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1677622389
transform 1 0 1708 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1677622389
transform 1 0 1732 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6062
timestamp 1677622389
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1677622389
transform 1 0 1820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1677622389
transform 1 0 1844 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5360
timestamp 1677622389
transform 1 0 1844 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1677622389
transform 1 0 1844 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5956
timestamp 1677622389
transform 1 0 1860 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5337
timestamp 1677622389
transform 1 0 1860 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1677622389
transform 1 0 1868 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1677622389
transform 1 0 1884 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1677622389
transform 1 0 1916 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5957
timestamp 1677622389
transform 1 0 1924 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5288
timestamp 1677622389
transform 1 0 1940 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6064
timestamp 1677622389
transform 1 0 1932 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1677622389
transform 1 0 1940 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5396
timestamp 1677622389
transform 1 0 1932 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5958
timestamp 1677622389
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1677622389
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1677622389
transform 1 0 2004 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5338
timestamp 1677622389
transform 1 0 2004 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5961
timestamp 1677622389
transform 1 0 2036 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5339
timestamp 1677622389
transform 1 0 2036 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1677622389
transform 1 0 2060 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6066
timestamp 1677622389
transform 1 0 2068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1677622389
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5362
timestamp 1677622389
transform 1 0 2068 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1677622389
transform 1 0 2108 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5962
timestamp 1677622389
transform 1 0 2100 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5249
timestamp 1677622389
transform 1 0 2132 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5963
timestamp 1677622389
transform 1 0 2116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1677622389
transform 1 0 2124 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5341
timestamp 1677622389
transform 1 0 2108 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1677622389
transform 1 0 2124 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6122
timestamp 1677622389
transform 1 0 2124 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5289
timestamp 1677622389
transform 1 0 2140 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5965
timestamp 1677622389
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1677622389
transform 1 0 2148 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5318
timestamp 1677622389
transform 1 0 2156 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6068
timestamp 1677622389
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5343
timestamp 1677622389
transform 1 0 2148 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1677622389
transform 1 0 2180 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1677622389
transform 1 0 2180 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6069
timestamp 1677622389
transform 1 0 2172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1677622389
transform 1 0 2180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1677622389
transform 1 0 2204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1677622389
transform 1 0 2220 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5344
timestamp 1677622389
transform 1 0 2204 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6071
timestamp 1677622389
transform 1 0 2228 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5363
timestamp 1677622389
transform 1 0 2228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1677622389
transform 1 0 2244 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6123
timestamp 1677622389
transform 1 0 2244 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1677622389
transform 1 0 2260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1677622389
transform 1 0 2260 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5250
timestamp 1677622389
transform 1 0 2300 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1677622389
transform 1 0 2292 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1677622389
transform 1 0 2324 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5970
timestamp 1677622389
transform 1 0 2316 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5319
timestamp 1677622389
transform 1 0 2324 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6073
timestamp 1677622389
transform 1 0 2308 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5347
timestamp 1677622389
transform 1 0 2316 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1677622389
transform 1 0 2348 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1677622389
transform 1 0 2340 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5971
timestamp 1677622389
transform 1 0 2348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1677622389
transform 1 0 2340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1677622389
transform 1 0 2364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1677622389
transform 1 0 2380 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5251
timestamp 1677622389
transform 1 0 2428 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1677622389
transform 1 0 2412 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5974
timestamp 1677622389
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1677622389
transform 1 0 2436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1677622389
transform 1 0 2412 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5364
timestamp 1677622389
transform 1 0 2412 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6076
timestamp 1677622389
transform 1 0 2452 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5365
timestamp 1677622389
transform 1 0 2452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1677622389
transform 1 0 2484 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5976
timestamp 1677622389
transform 1 0 2484 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5265
timestamp 1677622389
transform 1 0 2508 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1677622389
transform 1 0 2532 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5977
timestamp 1677622389
transform 1 0 2524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1677622389
transform 1 0 2532 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5235
timestamp 1677622389
transform 1 0 2572 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5978
timestamp 1677622389
transform 1 0 2548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1677622389
transform 1 0 2564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1677622389
transform 1 0 2572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1677622389
transform 1 0 2580 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5266
timestamp 1677622389
transform 1 0 2628 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5981
timestamp 1677622389
transform 1 0 2620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1677622389
transform 1 0 2636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1677622389
transform 1 0 2628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1677622389
transform 1 0 2636 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5294
timestamp 1677622389
transform 1 0 2692 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5983
timestamp 1677622389
transform 1 0 2692 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5267
timestamp 1677622389
transform 1 0 2788 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1677622389
transform 1 0 2740 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5984
timestamp 1677622389
transform 1 0 2740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1677622389
transform 1 0 2788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1677622389
transform 1 0 2708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1677622389
transform 1 0 2804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1677622389
transform 1 0 2796 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5366
timestamp 1677622389
transform 1 0 2796 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1677622389
transform 1 0 2836 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5909
timestamp 1677622389
transform 1 0 2844 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1677622389
transform 1 0 2844 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5367
timestamp 1677622389
transform 1 0 2844 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5987
timestamp 1677622389
transform 1 0 2860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1677622389
transform 1 0 2868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1677622389
transform 1 0 2884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1677622389
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5368
timestamp 1677622389
transform 1 0 2876 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5990
timestamp 1677622389
transform 1 0 2908 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5268
timestamp 1677622389
transform 1 0 2924 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5910
timestamp 1677622389
transform 1 0 2916 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5241
timestamp 1677622389
transform 1 0 2996 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1677622389
transform 1 0 2996 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5911
timestamp 1677622389
transform 1 0 2996 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1677622389
transform 1 0 2980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1677622389
transform 1 0 2972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5369
timestamp 1677622389
transform 1 0 2972 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6086
timestamp 1677622389
transform 1 0 3044 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5270
timestamp 1677622389
transform 1 0 3068 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6087
timestamp 1677622389
transform 1 0 3068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1677622389
transform 1 0 3100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1677622389
transform 1 0 3132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1677622389
transform 1 0 3140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1677622389
transform 1 0 3108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1677622389
transform 1 0 3124 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5370
timestamp 1677622389
transform 1 0 3100 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6124
timestamp 1677622389
transform 1 0 3116 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5371
timestamp 1677622389
transform 1 0 3124 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1677622389
transform 1 0 3164 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6090
timestamp 1677622389
transform 1 0 3156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1677622389
transform 1 0 3156 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1677622389
transform 1 0 3188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1677622389
transform 1 0 3172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1677622389
transform 1 0 3180 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5253
timestamp 1677622389
transform 1 0 3244 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5904
timestamp 1677622389
transform 1 0 3236 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_5372
timestamp 1677622389
transform 1 0 3236 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5912
timestamp 1677622389
transform 1 0 3252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1677622389
transform 1 0 3244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1677622389
transform 1 0 3260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1677622389
transform 1 0 3284 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_5296
timestamp 1677622389
transform 1 0 3284 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5906
timestamp 1677622389
transform 1 0 3300 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1677622389
transform 1 0 3292 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1677622389
transform 1 0 3300 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1677622389
transform 1 0 3276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1677622389
transform 1 0 3324 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1677622389
transform 1 0 3316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1677622389
transform 1 0 3356 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1677622389
transform 1 0 3340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1677622389
transform 1 0 3348 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5322
timestamp 1677622389
transform 1 0 3340 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6000
timestamp 1677622389
transform 1 0 3364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1677622389
transform 1 0 3388 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5323
timestamp 1677622389
transform 1 0 3388 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6093
timestamp 1677622389
transform 1 0 3380 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5297
timestamp 1677622389
transform 1 0 3404 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1677622389
transform 1 0 3436 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1677622389
transform 1 0 3444 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6001
timestamp 1677622389
transform 1 0 3436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1677622389
transform 1 0 3444 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5242
timestamp 1677622389
transform 1 0 3484 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1677622389
transform 1 0 3468 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6003
timestamp 1677622389
transform 1 0 3468 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5324
timestamp 1677622389
transform 1 0 3476 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6094
timestamp 1677622389
transform 1 0 3460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5348
timestamp 1677622389
transform 1 0 3476 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1677622389
transform 1 0 3508 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6095
timestamp 1677622389
transform 1 0 3484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1677622389
transform 1 0 3492 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5397
timestamp 1677622389
transform 1 0 3484 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1677622389
transform 1 0 3500 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6004
timestamp 1677622389
transform 1 0 3516 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5373
timestamp 1677622389
transform 1 0 3508 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1677622389
transform 1 0 3548 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1677622389
transform 1 0 3532 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1677622389
transform 1 0 3564 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1677622389
transform 1 0 3588 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6005
timestamp 1677622389
transform 1 0 3532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1677622389
transform 1 0 3588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1677622389
transform 1 0 3612 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5374
timestamp 1677622389
transform 1 0 3540 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1677622389
transform 1 0 3612 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1677622389
transform 1 0 3628 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6007
timestamp 1677622389
transform 1 0 3692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1677622389
transform 1 0 3644 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5376
timestamp 1677622389
transform 1 0 3644 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6008
timestamp 1677622389
transform 1 0 3740 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5243
timestamp 1677622389
transform 1 0 3756 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6009
timestamp 1677622389
transform 1 0 3764 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5244
timestamp 1677622389
transform 1 0 3796 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6010
timestamp 1677622389
transform 1 0 3804 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5350
timestamp 1677622389
transform 1 0 3812 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6099
timestamp 1677622389
transform 1 0 3852 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5377
timestamp 1677622389
transform 1 0 3852 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6011
timestamp 1677622389
transform 1 0 3916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1677622389
transform 1 0 3884 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5378
timestamp 1677622389
transform 1 0 3884 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1677622389
transform 1 0 3948 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1677622389
transform 1 0 3900 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6012
timestamp 1677622389
transform 1 0 3980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1677622389
transform 1 0 3996 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5325
timestamp 1677622389
transform 1 0 4020 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6014
timestamp 1677622389
transform 1 0 4052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1677622389
transform 1 0 4020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1677622389
transform 1 0 4028 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1677622389
transform 1 0 4044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1677622389
transform 1 0 4060 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5399
timestamp 1677622389
transform 1 0 4028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1677622389
transform 1 0 4132 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6015
timestamp 1677622389
transform 1 0 4156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1677622389
transform 1 0 4164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1677622389
transform 1 0 4180 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5400
timestamp 1677622389
transform 1 0 4180 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6016
timestamp 1677622389
transform 1 0 4212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1677622389
transform 1 0 4236 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5305
timestamp 1677622389
transform 1 0 4356 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6017
timestamp 1677622389
transform 1 0 4324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1677622389
transform 1 0 4284 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5401
timestamp 1677622389
transform 1 0 4284 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1677622389
transform 1 0 4404 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6018
timestamp 1677622389
transform 1 0 4412 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5380
timestamp 1677622389
transform 1 0 4396 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1677622389
transform 1 0 4412 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1677622389
transform 1 0 4428 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6019
timestamp 1677622389
transform 1 0 4428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1677622389
transform 1 0 4444 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5274
timestamp 1677622389
transform 1 0 4500 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1677622389
transform 1 0 4460 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1677622389
transform 1 0 4548 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6020
timestamp 1677622389
transform 1 0 4484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1677622389
transform 1 0 4540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1677622389
transform 1 0 4548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1677622389
transform 1 0 4460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5402
timestamp 1677622389
transform 1 0 4460 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1677622389
transform 1 0 4580 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1677622389
transform 1 0 4604 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1677622389
transform 1 0 4596 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1677622389
transform 1 0 4604 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6023
timestamp 1677622389
transform 1 0 4596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1677622389
transform 1 0 4612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1677622389
transform 1 0 4572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1677622389
transform 1 0 4588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1677622389
transform 1 0 4604 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5382
timestamp 1677622389
transform 1 0 4572 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1677622389
transform 1 0 4612 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1677622389
transform 1 0 4652 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1677622389
transform 1 0 4628 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_6025
timestamp 1677622389
transform 1 0 4652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1677622389
transform 1 0 4668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1677622389
transform 1 0 4628 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5351
timestamp 1677622389
transform 1 0 4636 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6115
timestamp 1677622389
transform 1 0 4644 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5352
timestamp 1677622389
transform 1 0 4652 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6116
timestamp 1677622389
transform 1 0 4660 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5309
timestamp 1677622389
transform 1 0 4780 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1677622389
transform 1 0 4676 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6027
timestamp 1677622389
transform 1 0 4716 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5330
timestamp 1677622389
transform 1 0 4756 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6028
timestamp 1677622389
transform 1 0 4772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1677622389
transform 1 0 4780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1677622389
transform 1 0 4676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1677622389
transform 1 0 4692 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5384
timestamp 1677622389
transform 1 0 4668 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1677622389
transform 1 0 4716 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1677622389
transform 1 0 4692 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6119
timestamp 1677622389
transform 1 0 4788 0 1 1805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_58
timestamp 1677622389
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_7030
timestamp 1677622389
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_7032
timestamp 1677622389
transform 1 0 80 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_391
timestamp 1677622389
transform 1 0 88 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_442
timestamp 1677622389
transform -1 0 200 0 1 1770
box -9 -3 26 105
use FILL  FILL_7033
timestamp 1677622389
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7034
timestamp 1677622389
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7035
timestamp 1677622389
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7036
timestamp 1677622389
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7037
timestamp 1677622389
transform 1 0 232 0 1 1770
box -8 -3 16 105
use FILL  FILL_7038
timestamp 1677622389
transform 1 0 240 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_83
timestamp 1677622389
transform -1 0 272 0 1 1770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_392
timestamp 1677622389
transform 1 0 272 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_5404
timestamp 1677622389
transform 1 0 380 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_443
timestamp 1677622389
transform 1 0 368 0 1 1770
box -9 -3 26 105
use FILL  FILL_7039
timestamp 1677622389
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7040
timestamp 1677622389
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_7052
timestamp 1677622389
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_7054
timestamp 1677622389
transform 1 0 408 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_445
timestamp 1677622389
transform 1 0 416 0 1 1770
box -9 -3 26 105
use FILL  FILL_7055
timestamp 1677622389
transform 1 0 432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7056
timestamp 1677622389
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_7057
timestamp 1677622389
transform 1 0 448 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5405
timestamp 1677622389
transform 1 0 484 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_272
timestamp 1677622389
transform -1 0 496 0 1 1770
box -8 -3 46 105
use FILL  FILL_7058
timestamp 1677622389
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7059
timestamp 1677622389
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7060
timestamp 1677622389
transform 1 0 512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7061
timestamp 1677622389
transform 1 0 520 0 1 1770
box -8 -3 16 105
use FILL  FILL_7062
timestamp 1677622389
transform 1 0 528 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_260
timestamp 1677622389
transform -1 0 576 0 1 1770
box -8 -3 46 105
use FILL  FILL_7063
timestamp 1677622389
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_7064
timestamp 1677622389
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7065
timestamp 1677622389
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7066
timestamp 1677622389
transform 1 0 600 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_30
timestamp 1677622389
transform -1 0 640 0 1 1770
box -8 -3 40 105
use FILL  FILL_7067
timestamp 1677622389
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_7068
timestamp 1677622389
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_7069
timestamp 1677622389
transform 1 0 656 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5406
timestamp 1677622389
transform 1 0 692 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_262
timestamp 1677622389
transform 1 0 664 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_5407
timestamp 1677622389
transform 1 0 716 0 1 1775
box -3 -3 3 3
use FILL  FILL_7078
timestamp 1677622389
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_7079
timestamp 1677622389
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_7080
timestamp 1677622389
transform 1 0 720 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_65
timestamp 1677622389
transform 1 0 728 0 1 1770
box -8 -3 32 105
use FILL  FILL_7081
timestamp 1677622389
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_7082
timestamp 1677622389
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_7083
timestamp 1677622389
transform 1 0 768 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_447
timestamp 1677622389
transform -1 0 792 0 1 1770
box -9 -3 26 105
use FILL  FILL_7084
timestamp 1677622389
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_7090
timestamp 1677622389
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_7092
timestamp 1677622389
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_7094
timestamp 1677622389
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_7096
timestamp 1677622389
transform 1 0 824 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_84
timestamp 1677622389
transform 1 0 832 0 1 1770
box -5 -3 28 105
use FILL  FILL_7097
timestamp 1677622389
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_7100
timestamp 1677622389
transform 1 0 864 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_86
timestamp 1677622389
transform 1 0 872 0 1 1770
box -5 -3 28 105
use FILL  FILL_7102
timestamp 1677622389
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_7103
timestamp 1677622389
transform 1 0 904 0 1 1770
box -8 -3 16 105
use FILL  FILL_7104
timestamp 1677622389
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7108
timestamp 1677622389
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_7110
timestamp 1677622389
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_7112
timestamp 1677622389
transform 1 0 936 0 1 1770
box -8 -3 16 105
use FILL  FILL_7114
timestamp 1677622389
transform 1 0 944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7116
timestamp 1677622389
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_7118
timestamp 1677622389
transform 1 0 960 0 1 1770
box -8 -3 16 105
use FILL  FILL_7119
timestamp 1677622389
transform 1 0 968 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_274
timestamp 1677622389
transform 1 0 976 0 1 1770
box -8 -3 46 105
use FILL  FILL_7120
timestamp 1677622389
transform 1 0 1016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7124
timestamp 1677622389
transform 1 0 1024 0 1 1770
box -8 -3 16 105
use FILL  FILL_7126
timestamp 1677622389
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_7128
timestamp 1677622389
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7130
timestamp 1677622389
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_7132
timestamp 1677622389
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_7134
timestamp 1677622389
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_396
timestamp 1677622389
transform 1 0 1072 0 1 1770
box -8 -3 104 105
use FILL  FILL_7136
timestamp 1677622389
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_7145
timestamp 1677622389
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_7147
timestamp 1677622389
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_7149
timestamp 1677622389
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7150
timestamp 1677622389
transform 1 0 1200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7151
timestamp 1677622389
transform 1 0 1208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7152
timestamp 1677622389
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7153
timestamp 1677622389
transform 1 0 1224 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_263
timestamp 1677622389
transform -1 0 1272 0 1 1770
box -8 -3 46 105
use FILL  FILL_7154
timestamp 1677622389
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_7162
timestamp 1677622389
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_7163
timestamp 1677622389
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use FILL  FILL_7164
timestamp 1677622389
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use FILL  FILL_7165
timestamp 1677622389
transform 1 0 1304 0 1 1770
box -8 -3 16 105
use FILL  FILL_7166
timestamp 1677622389
transform 1 0 1312 0 1 1770
box -8 -3 16 105
use FILL  FILL_7167
timestamp 1677622389
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_7170
timestamp 1677622389
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_7172
timestamp 1677622389
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_7174
timestamp 1677622389
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_7176
timestamp 1677622389
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5408
timestamp 1677622389
transform 1 0 1388 0 1 1775
box -3 -3 3 3
use AND2X2  AND2X2_33
timestamp 1677622389
transform -1 0 1392 0 1 1770
box -8 -3 40 105
use FILL  FILL_7177
timestamp 1677622389
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_7178
timestamp 1677622389
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_7179
timestamp 1677622389
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use FILL  FILL_7180
timestamp 1677622389
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_7181
timestamp 1677622389
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7182
timestamp 1677622389
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7189
timestamp 1677622389
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_449
timestamp 1677622389
transform 1 0 1448 0 1 1770
box -9 -3 26 105
use FILL  FILL_7191
timestamp 1677622389
transform 1 0 1464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7195
timestamp 1677622389
transform 1 0 1472 0 1 1770
box -8 -3 16 105
use FILL  FILL_7197
timestamp 1677622389
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_7199
timestamp 1677622389
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_7201
timestamp 1677622389
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7203
timestamp 1677622389
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_34
timestamp 1677622389
transform -1 0 1544 0 1 1770
box -8 -3 40 105
use FILL  FILL_7204
timestamp 1677622389
transform 1 0 1544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7211
timestamp 1677622389
transform 1 0 1552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7213
timestamp 1677622389
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_7215
timestamp 1677622389
transform 1 0 1568 0 1 1770
box -8 -3 16 105
use FILL  FILL_7217
timestamp 1677622389
transform 1 0 1576 0 1 1770
box -8 -3 16 105
use FILL  FILL_7219
timestamp 1677622389
transform 1 0 1584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7221
timestamp 1677622389
transform 1 0 1592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7223
timestamp 1677622389
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_7224
timestamp 1677622389
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_87
timestamp 1677622389
transform 1 0 1616 0 1 1770
box -5 -3 28 105
use FILL  FILL_7225
timestamp 1677622389
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use FILL  FILL_7227
timestamp 1677622389
transform 1 0 1648 0 1 1770
box -8 -3 16 105
use FILL  FILL_7229
timestamp 1677622389
transform 1 0 1656 0 1 1770
box -8 -3 16 105
use FILL  FILL_7231
timestamp 1677622389
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7233
timestamp 1677622389
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7235
timestamp 1677622389
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7237
timestamp 1677622389
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_7239
timestamp 1677622389
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_265
timestamp 1677622389
transform 1 0 1704 0 1 1770
box -8 -3 46 105
use FILL  FILL_7241
timestamp 1677622389
transform 1 0 1744 0 1 1770
box -8 -3 16 105
use FILL  FILL_7243
timestamp 1677622389
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_397
timestamp 1677622389
transform -1 0 1856 0 1 1770
box -8 -3 104 105
use FILL  FILL_7244
timestamp 1677622389
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_7254
timestamp 1677622389
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_7256
timestamp 1677622389
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7258
timestamp 1677622389
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_7259
timestamp 1677622389
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5409
timestamp 1677622389
transform 1 0 1916 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_450
timestamp 1677622389
transform -1 0 1912 0 1 1770
box -9 -3 26 105
use FILL  FILL_7260
timestamp 1677622389
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7261
timestamp 1677622389
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use FILL  FILL_7264
timestamp 1677622389
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_88
timestamp 1677622389
transform -1 0 1960 0 1 1770
box -5 -3 28 105
use FILL  FILL_7265
timestamp 1677622389
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_7266
timestamp 1677622389
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_7267
timestamp 1677622389
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_36
timestamp 1677622389
transform -1 0 2016 0 1 1770
box -8 -3 40 105
use FILL  FILL_7268
timestamp 1677622389
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5410
timestamp 1677622389
transform 1 0 2044 0 1 1775
box -3 -3 3 3
use FILL  FILL_7269
timestamp 1677622389
transform 1 0 2024 0 1 1770
box -8 -3 16 105
use FILL  FILL_7270
timestamp 1677622389
transform 1 0 2032 0 1 1770
box -8 -3 16 105
use FILL  FILL_7271
timestamp 1677622389
transform 1 0 2040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7279
timestamp 1677622389
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_7281
timestamp 1677622389
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_7283
timestamp 1677622389
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_89
timestamp 1677622389
transform -1 0 2096 0 1 1770
box -5 -3 28 105
use FILL  FILL_7284
timestamp 1677622389
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7285
timestamp 1677622389
transform 1 0 2104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7286
timestamp 1677622389
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5411
timestamp 1677622389
transform 1 0 2140 0 1 1775
box -3 -3 3 3
use NOR2X1  NOR2X1_68
timestamp 1677622389
transform 1 0 2120 0 1 1770
box -8 -3 32 105
use FILL  FILL_7290
timestamp 1677622389
transform 1 0 2144 0 1 1770
box -8 -3 16 105
use FILL  FILL_7291
timestamp 1677622389
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_451
timestamp 1677622389
transform -1 0 2176 0 1 1770
box -9 -3 26 105
use FILL  FILL_7292
timestamp 1677622389
transform 1 0 2176 0 1 1770
box -8 -3 16 105
use FILL  FILL_7293
timestamp 1677622389
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_41
timestamp 1677622389
transform 1 0 2192 0 1 1770
box -8 -3 40 105
use FILL  FILL_7299
timestamp 1677622389
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7302
timestamp 1677622389
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_70
timestamp 1677622389
transform 1 0 2240 0 1 1770
box -8 -3 32 105
use FILL  FILL_7304
timestamp 1677622389
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_7306
timestamp 1677622389
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_7308
timestamp 1677622389
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_7309
timestamp 1677622389
transform 1 0 2288 0 1 1770
box -8 -3 16 105
use FILL  FILL_7310
timestamp 1677622389
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_42
timestamp 1677622389
transform 1 0 2304 0 1 1770
box -8 -3 40 105
use FILL  FILL_7312
timestamp 1677622389
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_7313
timestamp 1677622389
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_44
timestamp 1677622389
transform 1 0 2352 0 1 1770
box -8 -3 40 105
use FILL  FILL_7316
timestamp 1677622389
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7322
timestamp 1677622389
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_7324
timestamp 1677622389
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_45
timestamp 1677622389
transform 1 0 2408 0 1 1770
box -8 -3 40 105
use FILL  FILL_7325
timestamp 1677622389
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_7326
timestamp 1677622389
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use FILL  FILL_7327
timestamp 1677622389
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_7330
timestamp 1677622389
transform 1 0 2464 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_47
timestamp 1677622389
transform 1 0 2472 0 1 1770
box -8 -3 40 105
use FILL  FILL_7332
timestamp 1677622389
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7335
timestamp 1677622389
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7336
timestamp 1677622389
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5412
timestamp 1677622389
transform 1 0 2540 0 1 1775
box -3 -3 3 3
use FILL  FILL_7337
timestamp 1677622389
transform 1 0 2528 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_48
timestamp 1677622389
transform 1 0 2536 0 1 1770
box -8 -3 40 105
use FILL  FILL_7338
timestamp 1677622389
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use FILL  FILL_7339
timestamp 1677622389
transform 1 0 2576 0 1 1770
box -8 -3 16 105
use FILL  FILL_7340
timestamp 1677622389
transform 1 0 2584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7341
timestamp 1677622389
transform 1 0 2592 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_279
timestamp 1677622389
transform 1 0 2600 0 1 1770
box -8 -3 46 105
use FILL  FILL_7342
timestamp 1677622389
transform 1 0 2640 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_455
timestamp 1677622389
transform 1 0 2648 0 1 1770
box -9 -3 26 105
use FILL  FILL_7350
timestamp 1677622389
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7354
timestamp 1677622389
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7356
timestamp 1677622389
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7357
timestamp 1677622389
transform 1 0 2688 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5413
timestamp 1677622389
transform 1 0 2708 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_398
timestamp 1677622389
transform 1 0 2696 0 1 1770
box -8 -3 104 105
use FILL  FILL_7358
timestamp 1677622389
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use FILL  FILL_7359
timestamp 1677622389
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_127
timestamp 1677622389
transform 1 0 2808 0 1 1770
box -8 -3 34 105
use M3_M2  M3_M2_5414
timestamp 1677622389
transform 1 0 2852 0 1 1775
box -3 -3 3 3
use FILL  FILL_7360
timestamp 1677622389
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_7369
timestamp 1677622389
transform 1 0 2848 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1677622389
transform 1 0 2856 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_457
timestamp 1677622389
transform 1 0 2880 0 1 1770
box -9 -3 26 105
use FILL  FILL_7370
timestamp 1677622389
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_7374
timestamp 1677622389
transform 1 0 2904 0 1 1770
box -8 -3 16 105
use FILL  FILL_7375
timestamp 1677622389
transform 1 0 2912 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_458
timestamp 1677622389
transform -1 0 2936 0 1 1770
box -9 -3 26 105
use FILL  FILL_7376
timestamp 1677622389
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_7377
timestamp 1677622389
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7378
timestamp 1677622389
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_7379
timestamp 1677622389
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_128
timestamp 1677622389
transform 1 0 2968 0 1 1770
box -8 -3 34 105
use FILL  FILL_7380
timestamp 1677622389
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_7381
timestamp 1677622389
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7384
timestamp 1677622389
transform 1 0 3016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7385
timestamp 1677622389
transform 1 0 3024 0 1 1770
box -8 -3 16 105
use FILL  FILL_7386
timestamp 1677622389
transform 1 0 3032 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_129
timestamp 1677622389
transform -1 0 3072 0 1 1770
box -8 -3 34 105
use FILL  FILL_7387
timestamp 1677622389
transform 1 0 3072 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5415
timestamp 1677622389
transform 1 0 3092 0 1 1775
box -3 -3 3 3
use AND2X2  AND2X2_49
timestamp 1677622389
transform -1 0 3112 0 1 1770
box -8 -3 40 105
use NOR2X1  NOR2X1_74
timestamp 1677622389
transform 1 0 3112 0 1 1770
box -8 -3 32 105
use M3_M2  M3_M2_5416
timestamp 1677622389
transform 1 0 3156 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_460
timestamp 1677622389
transform -1 0 3152 0 1 1770
box -9 -3 26 105
use FILL  FILL_7388
timestamp 1677622389
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_75
timestamp 1677622389
transform 1 0 3160 0 1 1770
box -8 -3 32 105
use FILL  FILL_7389
timestamp 1677622389
transform 1 0 3184 0 1 1770
box -8 -3 16 105
use FILL  FILL_7390
timestamp 1677622389
transform 1 0 3192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7402
timestamp 1677622389
transform 1 0 3200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7404
timestamp 1677622389
transform 1 0 3208 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_462
timestamp 1677622389
transform 1 0 3216 0 1 1770
box -9 -3 26 105
use FILL  FILL_7406
timestamp 1677622389
transform 1 0 3232 0 1 1770
box -8 -3 16 105
use FILL  FILL_7407
timestamp 1677622389
transform 1 0 3240 0 1 1770
box -8 -3 16 105
use FILL  FILL_7408
timestamp 1677622389
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_7409
timestamp 1677622389
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_54
timestamp 1677622389
transform 1 0 3264 0 1 1770
box -8 -3 40 105
use FILL  FILL_7412
timestamp 1677622389
transform 1 0 3296 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_55
timestamp 1677622389
transform 1 0 3304 0 1 1770
box -8 -3 40 105
use FILL  FILL_7418
timestamp 1677622389
transform 1 0 3336 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_56
timestamp 1677622389
transform -1 0 3376 0 1 1770
box -8 -3 40 105
use FILL  FILL_7419
timestamp 1677622389
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_7420
timestamp 1677622389
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_90
timestamp 1677622389
transform -1 0 3416 0 1 1770
box -5 -3 28 105
use FILL  FILL_7421
timestamp 1677622389
transform 1 0 3416 0 1 1770
box -8 -3 16 105
use FILL  FILL_7422
timestamp 1677622389
transform 1 0 3424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7423
timestamp 1677622389
transform 1 0 3432 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_91
timestamp 1677622389
transform 1 0 3440 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_92
timestamp 1677622389
transform 1 0 3464 0 1 1770
box -5 -3 28 105
use FILL  FILL_7430
timestamp 1677622389
transform 1 0 3488 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_466
timestamp 1677622389
transform 1 0 3496 0 1 1770
box -9 -3 26 105
use FILL  FILL_7434
timestamp 1677622389
transform 1 0 3512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7435
timestamp 1677622389
transform 1 0 3520 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_399
timestamp 1677622389
transform -1 0 3624 0 1 1770
box -8 -3 104 105
use FILL  FILL_7436
timestamp 1677622389
transform 1 0 3624 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_400
timestamp 1677622389
transform 1 0 3632 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_467
timestamp 1677622389
transform 1 0 3728 0 1 1770
box -9 -3 26 105
use FILL  FILL_7437
timestamp 1677622389
transform 1 0 3744 0 1 1770
box -8 -3 16 105
use FILL  FILL_7438
timestamp 1677622389
transform 1 0 3752 0 1 1770
box -8 -3 16 105
use FILL  FILL_7439
timestamp 1677622389
transform 1 0 3760 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_401
timestamp 1677622389
transform -1 0 3864 0 1 1770
box -8 -3 104 105
use FILL  FILL_7440
timestamp 1677622389
transform 1 0 3864 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_402
timestamp 1677622389
transform 1 0 3872 0 1 1770
box -8 -3 104 105
use FILL  FILL_7441
timestamp 1677622389
transform 1 0 3968 0 1 1770
box -8 -3 16 105
use FILL  FILL_7442
timestamp 1677622389
transform 1 0 3976 0 1 1770
box -8 -3 16 105
use FILL  FILL_7443
timestamp 1677622389
transform 1 0 3984 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_468
timestamp 1677622389
transform -1 0 4008 0 1 1770
box -9 -3 26 105
use FILL  FILL_7444
timestamp 1677622389
transform 1 0 4008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7445
timestamp 1677622389
transform 1 0 4016 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_267
timestamp 1677622389
transform 1 0 4024 0 1 1770
box -8 -3 46 105
use FILL  FILL_7446
timestamp 1677622389
transform 1 0 4064 0 1 1770
box -8 -3 16 105
use FILL  FILL_7447
timestamp 1677622389
transform 1 0 4072 0 1 1770
box -8 -3 16 105
use FILL  FILL_7448
timestamp 1677622389
transform 1 0 4080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7449
timestamp 1677622389
transform 1 0 4088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7450
timestamp 1677622389
transform 1 0 4096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7451
timestamp 1677622389
transform 1 0 4104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7452
timestamp 1677622389
transform 1 0 4112 0 1 1770
box -8 -3 16 105
use FILL  FILL_7453
timestamp 1677622389
transform 1 0 4120 0 1 1770
box -8 -3 16 105
use FILL  FILL_7475
timestamp 1677622389
transform 1 0 4128 0 1 1770
box -8 -3 16 105
use FILL  FILL_7477
timestamp 1677622389
transform 1 0 4136 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_272
timestamp 1677622389
transform -1 0 4184 0 1 1770
box -8 -3 46 105
use FILL  FILL_7478
timestamp 1677622389
transform 1 0 4184 0 1 1770
box -8 -3 16 105
use FILL  FILL_7479
timestamp 1677622389
transform 1 0 4192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7480
timestamp 1677622389
transform 1 0 4200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7481
timestamp 1677622389
transform 1 0 4208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7482
timestamp 1677622389
transform 1 0 4216 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_474
timestamp 1677622389
transform -1 0 4240 0 1 1770
box -9 -3 26 105
use FILL  FILL_7483
timestamp 1677622389
transform 1 0 4240 0 1 1770
box -8 -3 16 105
use FILL  FILL_7484
timestamp 1677622389
transform 1 0 4248 0 1 1770
box -8 -3 16 105
use FILL  FILL_7485
timestamp 1677622389
transform 1 0 4256 0 1 1770
box -8 -3 16 105
use FILL  FILL_7486
timestamp 1677622389
transform 1 0 4264 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_405
timestamp 1677622389
transform 1 0 4272 0 1 1770
box -8 -3 104 105
use FILL  FILL_7487
timestamp 1677622389
transform 1 0 4368 0 1 1770
box -8 -3 16 105
use FILL  FILL_7499
timestamp 1677622389
transform 1 0 4376 0 1 1770
box -8 -3 16 105
use FILL  FILL_7501
timestamp 1677622389
transform 1 0 4384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7503
timestamp 1677622389
transform 1 0 4392 0 1 1770
box -8 -3 16 105
use FILL  FILL_7505
timestamp 1677622389
transform 1 0 4400 0 1 1770
box -8 -3 16 105
use FILL  FILL_7506
timestamp 1677622389
transform 1 0 4408 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_476
timestamp 1677622389
transform -1 0 4432 0 1 1770
box -9 -3 26 105
use FILL  FILL_7507
timestamp 1677622389
transform 1 0 4432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7511
timestamp 1677622389
transform 1 0 4440 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_407
timestamp 1677622389
transform 1 0 4448 0 1 1770
box -8 -3 104 105
use FILL  FILL_7513
timestamp 1677622389
transform 1 0 4544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7520
timestamp 1677622389
transform 1 0 4552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7522
timestamp 1677622389
transform 1 0 4560 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_275
timestamp 1677622389
transform 1 0 4568 0 1 1770
box -8 -3 46 105
use FILL  FILL_7524
timestamp 1677622389
transform 1 0 4608 0 1 1770
box -8 -3 16 105
use FILL  FILL_7526
timestamp 1677622389
transform 1 0 4616 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5417
timestamp 1677622389
transform 1 0 4644 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_277
timestamp 1677622389
transform 1 0 4624 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_479
timestamp 1677622389
transform -1 0 4680 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5418
timestamp 1677622389
transform 1 0 4740 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_408
timestamp 1677622389
transform 1 0 4680 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_480
timestamp 1677622389
transform -1 0 4792 0 1 1770
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_59
timestamp 1677622389
transform 1 0 4819 0 1 1770
box -10 -3 10 3
use M3_M2  M3_M2_5419
timestamp 1677622389
transform 1 0 100 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1677622389
transform 1 0 156 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6133
timestamp 1677622389
transform 1 0 92 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5436
timestamp 1677622389
transform 1 0 180 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6134
timestamp 1677622389
transform 1 0 180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1677622389
transform 1 0 116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1677622389
transform 1 0 172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1677622389
transform 1 0 180 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5542
timestamp 1677622389
transform 1 0 172 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6135
timestamp 1677622389
transform 1 0 228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1677622389
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1677622389
transform 1 0 220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1677622389
transform 1 0 236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1677622389
transform 1 0 244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5584
timestamp 1677622389
transform 1 0 236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1677622389
transform 1 0 332 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6136
timestamp 1677622389
transform 1 0 308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1677622389
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1677622389
transform 1 0 332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1677622389
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5518
timestamp 1677622389
transform 1 0 332 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1677622389
transform 1 0 388 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1677622389
transform 1 0 364 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6139
timestamp 1677622389
transform 1 0 364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1677622389
transform 1 0 380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1677622389
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1677622389
transform 1 0 340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1677622389
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1677622389
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1677622389
transform 1 0 372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1677622389
transform 1 0 388 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5543
timestamp 1677622389
transform 1 0 316 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1677622389
transform 1 0 340 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1677622389
transform 1 0 388 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1677622389
transform 1 0 404 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1677622389
transform 1 0 428 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1677622389
transform 1 0 452 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6142
timestamp 1677622389
transform 1 0 436 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5500
timestamp 1677622389
transform 1 0 444 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6143
timestamp 1677622389
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5520
timestamp 1677622389
transform 1 0 420 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6242
timestamp 1677622389
transform 1 0 428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1677622389
transform 1 0 444 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5545
timestamp 1677622389
transform 1 0 444 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6144
timestamp 1677622389
transform 1 0 508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1677622389
transform 1 0 516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1677622389
transform 1 0 500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1677622389
transform 1 0 508 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5521
timestamp 1677622389
transform 1 0 516 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6246
timestamp 1677622389
transform 1 0 524 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5546
timestamp 1677622389
transform 1 0 500 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1677622389
transform 1 0 508 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1677622389
transform 1 0 500 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1677622389
transform 1 0 548 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1677622389
transform 1 0 556 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6146
timestamp 1677622389
transform 1 0 556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1677622389
transform 1 0 556 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5467
timestamp 1677622389
transform 1 0 652 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6147
timestamp 1677622389
transform 1 0 572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1677622389
transform 1 0 596 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5522
timestamp 1677622389
transform 1 0 604 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6249
timestamp 1677622389
transform 1 0 652 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5547
timestamp 1677622389
transform 1 0 596 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1677622389
transform 1 0 772 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6148
timestamp 1677622389
transform 1 0 772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1677622389
transform 1 0 692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1677622389
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5469
timestamp 1677622389
transform 1 0 796 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6149
timestamp 1677622389
transform 1 0 796 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5587
timestamp 1677622389
transform 1 0 836 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1677622389
transform 1 0 860 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6126
timestamp 1677622389
transform 1 0 860 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1677622389
transform 1 0 852 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5470
timestamp 1677622389
transform 1 0 868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1677622389
transform 1 0 892 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1677622389
transform 1 0 940 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6150
timestamp 1677622389
transform 1 0 932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1677622389
transform 1 0 956 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5588
timestamp 1677622389
transform 1 0 956 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1677622389
transform 1 0 988 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1677622389
transform 1 0 1012 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1677622389
transform 1 0 980 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1677622389
transform 1 0 1004 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6127
timestamp 1677622389
transform 1 0 1012 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1677622389
transform 1 0 980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1677622389
transform 1 0 996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1677622389
transform 1 0 1004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1677622389
transform 1 0 972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1677622389
transform 1 0 988 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5615
timestamp 1677622389
transform 1 0 988 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1677622389
transform 1 0 1012 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6256
timestamp 1677622389
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5473
timestamp 1677622389
transform 1 0 1100 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6257
timestamp 1677622389
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1677622389
transform 1 0 1124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1677622389
transform 1 0 1116 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5605
timestamp 1677622389
transform 1 0 1132 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6259
timestamp 1677622389
transform 1 0 1180 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5606
timestamp 1677622389
transform 1 0 1180 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1677622389
transform 1 0 1228 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6155
timestamp 1677622389
transform 1 0 1228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1677622389
transform 1 0 1220 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5523
timestamp 1677622389
transform 1 0 1228 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6261
timestamp 1677622389
transform 1 0 1252 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5502
timestamp 1677622389
transform 1 0 1308 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6156
timestamp 1677622389
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1677622389
transform 1 0 1324 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5524
timestamp 1677622389
transform 1 0 1300 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6262
timestamp 1677622389
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1677622389
transform 1 0 1316 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1677622389
transform 1 0 1340 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5503
timestamp 1677622389
transform 1 0 1372 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1677622389
transform 1 0 1396 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6158
timestamp 1677622389
transform 1 0 1420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1677622389
transform 1 0 1396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1677622389
transform 1 0 1412 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5548
timestamp 1677622389
transform 1 0 1396 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6265
timestamp 1677622389
transform 1 0 1436 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5549
timestamp 1677622389
transform 1 0 1444 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6159
timestamp 1677622389
transform 1 0 1468 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5443
timestamp 1677622389
transform 1 0 1532 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1677622389
transform 1 0 1532 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1677622389
transform 1 0 1564 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1677622389
transform 1 0 1620 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6160
timestamp 1677622389
transform 1 0 1604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1677622389
transform 1 0 1620 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5526
timestamp 1677622389
transform 1 0 1604 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6266
timestamp 1677622389
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1677622389
transform 1 0 1628 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5527
timestamp 1677622389
transform 1 0 1636 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1677622389
transform 1 0 1612 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6162
timestamp 1677622389
transform 1 0 1700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1677622389
transform 1 0 1692 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5528
timestamp 1677622389
transform 1 0 1700 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1677622389
transform 1 0 1716 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6163
timestamp 1677622389
transform 1 0 1716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1677622389
transform 1 0 1732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1677622389
transform 1 0 1724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1677622389
transform 1 0 1740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1677622389
transform 1 0 1756 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5529
timestamp 1677622389
transform 1 0 1756 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6271
timestamp 1677622389
transform 1 0 1804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1677622389
transform 1 0 1820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1677622389
transform 1 0 1836 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5425
timestamp 1677622389
transform 1 0 1908 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6166
timestamp 1677622389
transform 1 0 1916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1677622389
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1677622389
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5589
timestamp 1677622389
transform 1 0 1932 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1677622389
transform 1 0 1940 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1677622389
transform 1 0 1956 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1677622389
transform 1 0 1980 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6276
timestamp 1677622389
transform 1 0 1956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1677622389
transform 1 0 1972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1677622389
transform 1 0 1980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5551
timestamp 1677622389
transform 1 0 1956 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1677622389
transform 1 0 2012 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1677622389
transform 1 0 2004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1677622389
transform 1 0 2036 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6167
timestamp 1677622389
transform 1 0 2036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1677622389
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5552
timestamp 1677622389
transform 1 0 2028 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6280
timestamp 1677622389
transform 1 0 2044 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5590
timestamp 1677622389
transform 1 0 2060 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1677622389
transform 1 0 2092 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1677622389
transform 1 0 2108 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6168
timestamp 1677622389
transform 1 0 2108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1677622389
transform 1 0 2100 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5553
timestamp 1677622389
transform 1 0 2100 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1677622389
transform 1 0 2172 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6169
timestamp 1677622389
transform 1 0 2180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1677622389
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1677622389
transform 1 0 2172 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5591
timestamp 1677622389
transform 1 0 2164 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1677622389
transform 1 0 2220 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6128
timestamp 1677622389
transform 1 0 2220 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1677622389
transform 1 0 2212 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5508
timestamp 1677622389
transform 1 0 2220 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6284
timestamp 1677622389
transform 1 0 2204 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5530
timestamp 1677622389
transform 1 0 2212 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1677622389
transform 1 0 2244 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6129
timestamp 1677622389
transform 1 0 2244 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1677622389
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5554
timestamp 1677622389
transform 1 0 2244 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1677622389
transform 1 0 2268 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6172
timestamp 1677622389
transform 1 0 2268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1677622389
transform 1 0 2260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1677622389
transform 1 0 2292 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5448
timestamp 1677622389
transform 1 0 2324 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6173
timestamp 1677622389
transform 1 0 2308 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5509
timestamp 1677622389
transform 1 0 2316 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6287
timestamp 1677622389
transform 1 0 2324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1677622389
transform 1 0 2340 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5427
timestamp 1677622389
transform 1 0 2364 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1677622389
transform 1 0 2412 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6174
timestamp 1677622389
transform 1 0 2436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1677622389
transform 1 0 2444 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1677622389
transform 1 0 2412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1677622389
transform 1 0 2428 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5555
timestamp 1677622389
transform 1 0 2436 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1677622389
transform 1 0 2484 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6176
timestamp 1677622389
transform 1 0 2484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1677622389
transform 1 0 2492 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5556
timestamp 1677622389
transform 1 0 2492 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6347
timestamp 1677622389
transform 1 0 2508 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5429
timestamp 1677622389
transform 1 0 2548 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1677622389
transform 1 0 2532 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6292
timestamp 1677622389
transform 1 0 2540 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5557
timestamp 1677622389
transform 1 0 2540 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6348
timestamp 1677622389
transform 1 0 2548 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1677622389
transform 1 0 2556 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1677622389
transform 1 0 2532 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5609
timestamp 1677622389
transform 1 0 2548 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6293
timestamp 1677622389
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5558
timestamp 1677622389
transform 1 0 2588 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6362
timestamp 1677622389
transform 1 0 2580 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5610
timestamp 1677622389
transform 1 0 2580 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6177
timestamp 1677622389
transform 1 0 2604 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5532
timestamp 1677622389
transform 1 0 2604 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1677622389
transform 1 0 2604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1677622389
transform 1 0 2660 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6363
timestamp 1677622389
transform 1 0 2644 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5593
timestamp 1677622389
transform 1 0 2652 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6294
timestamp 1677622389
transform 1 0 2692 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5559
timestamp 1677622389
transform 1 0 2692 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6350
timestamp 1677622389
transform 1 0 2708 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1677622389
transform 1 0 2716 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1677622389
transform 1 0 2700 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5611
timestamp 1677622389
transform 1 0 2700 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1677622389
transform 1 0 2716 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6365
timestamp 1677622389
transform 1 0 2724 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5612
timestamp 1677622389
transform 1 0 2724 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6295
timestamp 1677622389
transform 1 0 2756 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5560
timestamp 1677622389
transform 1 0 2756 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6178
timestamp 1677622389
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1677622389
transform 1 0 2796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1677622389
transform 1 0 2804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5534
timestamp 1677622389
transform 1 0 2812 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6352
timestamp 1677622389
transform 1 0 2828 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1677622389
transform 1 0 2844 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5430
timestamp 1677622389
transform 1 0 2860 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1677622389
transform 1 0 2852 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1677622389
transform 1 0 2868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1677622389
transform 1 0 2884 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6298
timestamp 1677622389
transform 1 0 2876 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5431
timestamp 1677622389
transform 1 0 2900 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6299
timestamp 1677622389
transform 1 0 2892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1677622389
transform 1 0 2900 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1677622389
transform 1 0 2908 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5449
timestamp 1677622389
transform 1 0 2932 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1677622389
transform 1 0 2924 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6179
timestamp 1677622389
transform 1 0 2924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1677622389
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1677622389
transform 1 0 2924 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5450
timestamp 1677622389
transform 1 0 2988 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1677622389
transform 1 0 2980 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6181
timestamp 1677622389
transform 1 0 2980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1677622389
transform 1 0 2988 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5451
timestamp 1677622389
transform 1 0 3012 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1677622389
transform 1 0 3004 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6131
timestamp 1677622389
transform 1 0 3012 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1677622389
transform 1 0 2980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1677622389
transform 1 0 2996 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5562
timestamp 1677622389
transform 1 0 2980 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6354
timestamp 1677622389
transform 1 0 3004 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5484
timestamp 1677622389
transform 1 0 3036 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6183
timestamp 1677622389
transform 1 0 3028 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5563
timestamp 1677622389
transform 1 0 3020 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6184
timestamp 1677622389
transform 1 0 3044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1677622389
transform 1 0 3036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1677622389
transform 1 0 3044 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5564
timestamp 1677622389
transform 1 0 3044 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6185
timestamp 1677622389
transform 1 0 3076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1677622389
transform 1 0 3092 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1677622389
transform 1 0 3116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1677622389
transform 1 0 3132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1677622389
transform 1 0 3140 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5595
timestamp 1677622389
transform 1 0 3132 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6187
timestamp 1677622389
transform 1 0 3156 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5535
timestamp 1677622389
transform 1 0 3156 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1677622389
transform 1 0 3188 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1677622389
transform 1 0 3180 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6306
timestamp 1677622389
transform 1 0 3180 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5565
timestamp 1677622389
transform 1 0 3180 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6356
timestamp 1677622389
transform 1 0 3188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1677622389
transform 1 0 3172 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5596
timestamp 1677622389
transform 1 0 3188 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6357
timestamp 1677622389
transform 1 0 3212 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5432
timestamp 1677622389
transform 1 0 3228 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1677622389
transform 1 0 3252 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1677622389
transform 1 0 3236 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6307
timestamp 1677622389
transform 1 0 3244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5566
timestamp 1677622389
transform 1 0 3244 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1677622389
transform 1 0 3260 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6358
timestamp 1677622389
transform 1 0 3252 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1677622389
transform 1 0 3236 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1677622389
transform 1 0 3260 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5487
timestamp 1677622389
transform 1 0 3316 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6359
timestamp 1677622389
transform 1 0 3324 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5488
timestamp 1677622389
transform 1 0 3340 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6308
timestamp 1677622389
transform 1 0 3340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1677622389
transform 1 0 3348 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1677622389
transform 1 0 3364 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5616
timestamp 1677622389
transform 1 0 3356 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1677622389
transform 1 0 3380 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1677622389
transform 1 0 3372 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1677622389
transform 1 0 3380 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6188
timestamp 1677622389
transform 1 0 3388 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5512
timestamp 1677622389
transform 1 0 3396 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6189
timestamp 1677622389
transform 1 0 3412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1677622389
transform 1 0 3428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1677622389
transform 1 0 3372 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1677622389
transform 1 0 3396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1677622389
transform 1 0 3404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1677622389
transform 1 0 3420 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5567
timestamp 1677622389
transform 1 0 3420 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1677622389
transform 1 0 3396 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1677622389
transform 1 0 3388 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6313
timestamp 1677622389
transform 1 0 3436 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5618
timestamp 1677622389
transform 1 0 3444 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1677622389
transform 1 0 3460 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6191
timestamp 1677622389
transform 1 0 3460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1677622389
transform 1 0 3460 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5568
timestamp 1677622389
transform 1 0 3460 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6315
timestamp 1677622389
transform 1 0 3476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5598
timestamp 1677622389
transform 1 0 3476 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6192
timestamp 1677622389
transform 1 0 3508 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5491
timestamp 1677622389
transform 1 0 3596 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6193
timestamp 1677622389
transform 1 0 3548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1677622389
transform 1 0 3516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1677622389
transform 1 0 3532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1677622389
transform 1 0 3596 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5569
timestamp 1677622389
transform 1 0 3548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1677622389
transform 1 0 3596 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6194
timestamp 1677622389
transform 1 0 3668 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5492
timestamp 1677622389
transform 1 0 3700 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6195
timestamp 1677622389
transform 1 0 3700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1677622389
transform 1 0 3716 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5537
timestamp 1677622389
transform 1 0 3684 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6319
timestamp 1677622389
transform 1 0 3692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1677622389
transform 1 0 3708 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5538
timestamp 1677622389
transform 1 0 3716 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1677622389
transform 1 0 3692 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1677622389
transform 1 0 3708 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6321
timestamp 1677622389
transform 1 0 3740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1677622389
transform 1 0 3764 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5572
timestamp 1677622389
transform 1 0 3756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1677622389
transform 1 0 3780 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6198
timestamp 1677622389
transform 1 0 3780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1677622389
transform 1 0 3796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1677622389
transform 1 0 3804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5600
timestamp 1677622389
transform 1 0 3788 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1677622389
transform 1 0 3836 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1677622389
transform 1 0 3828 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6200
timestamp 1677622389
transform 1 0 3828 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1677622389
transform 1 0 3836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1677622389
transform 1 0 3852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1677622389
transform 1 0 3844 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5456
timestamp 1677622389
transform 1 0 3900 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1677622389
transform 1 0 3932 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6203
timestamp 1677622389
transform 1 0 3876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1677622389
transform 1 0 3892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1677622389
transform 1 0 3900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1677622389
transform 1 0 3916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1677622389
transform 1 0 3932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1677622389
transform 1 0 3860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1677622389
transform 1 0 3884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1677622389
transform 1 0 3900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1677622389
transform 1 0 3924 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5573
timestamp 1677622389
transform 1 0 3852 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1677622389
transform 1 0 3900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1677622389
transform 1 0 3924 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6328
timestamp 1677622389
transform 1 0 3940 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5575
timestamp 1677622389
transform 1 0 3940 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6208
timestamp 1677622389
transform 1 0 3980 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5457
timestamp 1677622389
transform 1 0 4004 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1677622389
transform 1 0 4004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1677622389
transform 1 0 4020 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1677622389
transform 1 0 4060 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6209
timestamp 1677622389
transform 1 0 4020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1677622389
transform 1 0 4044 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5539
timestamp 1677622389
transform 1 0 4052 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6210
timestamp 1677622389
transform 1 0 4116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1677622389
transform 1 0 4100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1677622389
transform 1 0 4116 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5576
timestamp 1677622389
transform 1 0 4020 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1677622389
transform 1 0 4044 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1677622389
transform 1 0 4108 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1677622389
transform 1 0 4148 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1677622389
transform 1 0 4164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1677622389
transform 1 0 4244 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6211
timestamp 1677622389
transform 1 0 4164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1677622389
transform 1 0 4188 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5579
timestamp 1677622389
transform 1 0 4188 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6212
timestamp 1677622389
transform 1 0 4268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1677622389
transform 1 0 4252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1677622389
transform 1 0 4260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5461
timestamp 1677622389
transform 1 0 4308 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6213
timestamp 1677622389
transform 1 0 4308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1677622389
transform 1 0 4324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1677622389
transform 1 0 4316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1677622389
transform 1 0 4332 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5580
timestamp 1677622389
transform 1 0 4316 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1677622389
transform 1 0 4332 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6337
timestamp 1677622389
transform 1 0 4348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1677622389
transform 1 0 4356 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5581
timestamp 1677622389
transform 1 0 4348 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1677622389
transform 1 0 4372 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1677622389
transform 1 0 4388 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6216
timestamp 1677622389
transform 1 0 4388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1677622389
transform 1 0 4396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1677622389
transform 1 0 4420 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5462
timestamp 1677622389
transform 1 0 4436 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6218
timestamp 1677622389
transform 1 0 4436 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5497
timestamp 1677622389
transform 1 0 4484 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6219
timestamp 1677622389
transform 1 0 4468 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5514
timestamp 1677622389
transform 1 0 4476 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6220
timestamp 1677622389
transform 1 0 4484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1677622389
transform 1 0 4460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1677622389
transform 1 0 4476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5582
timestamp 1677622389
transform 1 0 4460 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1677622389
transform 1 0 4476 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6341
timestamp 1677622389
transform 1 0 4516 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5583
timestamp 1677622389
transform 1 0 4516 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6221
timestamp 1677622389
transform 1 0 4540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1677622389
transform 1 0 4532 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5515
timestamp 1677622389
transform 1 0 4556 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1677622389
transform 1 0 4588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1677622389
transform 1 0 4612 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6222
timestamp 1677622389
transform 1 0 4572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1677622389
transform 1 0 4588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1677622389
transform 1 0 4604 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5540
timestamp 1677622389
transform 1 0 4580 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6343
timestamp 1677622389
transform 1 0 4596 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5434
timestamp 1677622389
transform 1 0 4628 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6225
timestamp 1677622389
transform 1 0 4628 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5463
timestamp 1677622389
transform 1 0 4668 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1677622389
transform 1 0 4644 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6226
timestamp 1677622389
transform 1 0 4652 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5517
timestamp 1677622389
transform 1 0 4660 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6227
timestamp 1677622389
transform 1 0 4668 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5541
timestamp 1677622389
transform 1 0 4652 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6344
timestamp 1677622389
transform 1 0 4660 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5435
timestamp 1677622389
transform 1 0 4716 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6228
timestamp 1677622389
transform 1 0 4764 0 1 1735
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_60
timestamp 1677622389
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_7031
timestamp 1677622389
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_393
timestamp 1677622389
transform 1 0 80 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7041
timestamp 1677622389
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7042
timestamp 1677622389
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7043
timestamp 1677622389
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_270
timestamp 1677622389
transform -1 0 240 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7044
timestamp 1677622389
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7045
timestamp 1677622389
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7046
timestamp 1677622389
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_444
timestamp 1677622389
transform -1 0 280 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7047
timestamp 1677622389
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7048
timestamp 1677622389
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7049
timestamp 1677622389
transform 1 0 296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7050
timestamp 1677622389
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_259
timestamp 1677622389
transform -1 0 352 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_271
timestamp 1677622389
transform -1 0 392 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7051
timestamp 1677622389
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7053
timestamp 1677622389
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7070
timestamp 1677622389
transform 1 0 408 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_261
timestamp 1677622389
transform -1 0 456 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7071
timestamp 1677622389
transform 1 0 456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7072
timestamp 1677622389
transform 1 0 464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7073
timestamp 1677622389
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7074
timestamp 1677622389
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_446
timestamp 1677622389
transform -1 0 504 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_273
timestamp 1677622389
transform 1 0 504 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7075
timestamp 1677622389
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7076
timestamp 1677622389
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_394
timestamp 1677622389
transform 1 0 560 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7077
timestamp 1677622389
transform 1 0 656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7085
timestamp 1677622389
transform 1 0 664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7086
timestamp 1677622389
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7087
timestamp 1677622389
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_395
timestamp 1677622389
transform -1 0 784 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7088
timestamp 1677622389
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7089
timestamp 1677622389
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7091
timestamp 1677622389
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7093
timestamp 1677622389
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7095
timestamp 1677622389
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7098
timestamp 1677622389
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_85
timestamp 1677622389
transform -1 0 856 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7099
timestamp 1677622389
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7101
timestamp 1677622389
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7105
timestamp 1677622389
transform 1 0 872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7106
timestamp 1677622389
transform 1 0 880 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_66
timestamp 1677622389
transform 1 0 888 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7107
timestamp 1677622389
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7109
timestamp 1677622389
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5619
timestamp 1677622389
transform 1 0 940 0 1 1675
box -3 -3 3 3
use FILL  FILL_7111
timestamp 1677622389
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7113
timestamp 1677622389
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7115
timestamp 1677622389
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7117
timestamp 1677622389
transform 1 0 952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7121
timestamp 1677622389
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5620
timestamp 1677622389
transform 1 0 988 0 1 1675
box -3 -3 3 3
use AOI22X1  AOI22X1_275
timestamp 1677622389
transform -1 0 1008 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7122
timestamp 1677622389
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7123
timestamp 1677622389
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7125
timestamp 1677622389
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7127
timestamp 1677622389
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7129
timestamp 1677622389
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7131
timestamp 1677622389
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7133
timestamp 1677622389
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7135
timestamp 1677622389
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_67
timestamp 1677622389
transform 1 0 1072 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7137
timestamp 1677622389
transform 1 0 1096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7138
timestamp 1677622389
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7139
timestamp 1677622389
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7140
timestamp 1677622389
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7141
timestamp 1677622389
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_448
timestamp 1677622389
transform 1 0 1136 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7142
timestamp 1677622389
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7143
timestamp 1677622389
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7144
timestamp 1677622389
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7146
timestamp 1677622389
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7148
timestamp 1677622389
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7155
timestamp 1677622389
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_31
timestamp 1677622389
transform -1 0 1232 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7156
timestamp 1677622389
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7157
timestamp 1677622389
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7158
timestamp 1677622389
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7159
timestamp 1677622389
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7160
timestamp 1677622389
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7161
timestamp 1677622389
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7168
timestamp 1677622389
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_32
timestamp 1677622389
transform -1 0 1320 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7169
timestamp 1677622389
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7171
timestamp 1677622389
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7173
timestamp 1677622389
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7175
timestamp 1677622389
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7183
timestamp 1677622389
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7184
timestamp 1677622389
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7185
timestamp 1677622389
transform 1 0 1368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7186
timestamp 1677622389
transform 1 0 1376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7187
timestamp 1677622389
transform 1 0 1384 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_276
timestamp 1677622389
transform -1 0 1432 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7188
timestamp 1677622389
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7190
timestamp 1677622389
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7192
timestamp 1677622389
transform 1 0 1448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7193
timestamp 1677622389
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7194
timestamp 1677622389
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7196
timestamp 1677622389
transform 1 0 1472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7198
timestamp 1677622389
transform 1 0 1480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7200
timestamp 1677622389
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7202
timestamp 1677622389
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7205
timestamp 1677622389
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7206
timestamp 1677622389
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7207
timestamp 1677622389
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7208
timestamp 1677622389
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7209
timestamp 1677622389
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7210
timestamp 1677622389
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7212
timestamp 1677622389
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7214
timestamp 1677622389
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7216
timestamp 1677622389
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7218
timestamp 1677622389
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7220
timestamp 1677622389
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7222
timestamp 1677622389
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_264
timestamp 1677622389
transform 1 0 1600 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7226
timestamp 1677622389
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7228
timestamp 1677622389
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7230
timestamp 1677622389
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7232
timestamp 1677622389
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7234
timestamp 1677622389
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7236
timestamp 1677622389
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7238
timestamp 1677622389
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7240
timestamp 1677622389
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_277
timestamp 1677622389
transform 1 0 1704 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7242
timestamp 1677622389
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7245
timestamp 1677622389
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7246
timestamp 1677622389
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7247
timestamp 1677622389
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7248
timestamp 1677622389
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7249
timestamp 1677622389
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7250
timestamp 1677622389
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_278
timestamp 1677622389
transform -1 0 1840 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7251
timestamp 1677622389
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7252
timestamp 1677622389
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7253
timestamp 1677622389
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5621
timestamp 1677622389
transform 1 0 1876 0 1 1675
box -3 -3 3 3
use FILL  FILL_7255
timestamp 1677622389
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7257
timestamp 1677622389
transform 1 0 1872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7262
timestamp 1677622389
transform 1 0 1880 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_35
timestamp 1677622389
transform -1 0 1920 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7263
timestamp 1677622389
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7272
timestamp 1677622389
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7273
timestamp 1677622389
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_37
timestamp 1677622389
transform 1 0 1944 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7274
timestamp 1677622389
transform 1 0 1976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7275
timestamp 1677622389
transform 1 0 1984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7276
timestamp 1677622389
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7277
timestamp 1677622389
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5622
timestamp 1677622389
transform 1 0 2044 0 1 1675
box -3 -3 3 3
use AND2X2  AND2X2_38
timestamp 1677622389
transform -1 0 2040 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7278
timestamp 1677622389
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7280
timestamp 1677622389
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7282
timestamp 1677622389
transform 1 0 2056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7287
timestamp 1677622389
transform 1 0 2064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7288
timestamp 1677622389
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_39
timestamp 1677622389
transform -1 0 2112 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7289
timestamp 1677622389
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7294
timestamp 1677622389
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7295
timestamp 1677622389
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7296
timestamp 1677622389
transform 1 0 2136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7297
timestamp 1677622389
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_40
timestamp 1677622389
transform -1 0 2184 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7298
timestamp 1677622389
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7300
timestamp 1677622389
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_69
timestamp 1677622389
transform -1 0 2224 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7301
timestamp 1677622389
transform 1 0 2224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7303
timestamp 1677622389
transform 1 0 2232 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_71
timestamp 1677622389
transform 1 0 2240 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7305
timestamp 1677622389
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7307
timestamp 1677622389
transform 1 0 2272 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_452
timestamp 1677622389
transform 1 0 2280 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7311
timestamp 1677622389
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7314
timestamp 1677622389
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_43
timestamp 1677622389
transform 1 0 2312 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7315
timestamp 1677622389
transform 1 0 2344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7317
timestamp 1677622389
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7318
timestamp 1677622389
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7319
timestamp 1677622389
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7320
timestamp 1677622389
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7321
timestamp 1677622389
transform 1 0 2384 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5623
timestamp 1677622389
transform 1 0 2404 0 1 1675
box -3 -3 3 3
use FILL  FILL_7323
timestamp 1677622389
transform 1 0 2392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7328
timestamp 1677622389
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_46
timestamp 1677622389
transform -1 0 2440 0 -1 1770
box -8 -3 40 105
use INVX2  INVX2_453
timestamp 1677622389
transform 1 0 2440 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7329
timestamp 1677622389
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7331
timestamp 1677622389
transform 1 0 2464 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_72
timestamp 1677622389
transform 1 0 2472 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7333
timestamp 1677622389
transform 1 0 2496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7334
timestamp 1677622389
transform 1 0 2504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7343
timestamp 1677622389
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_47
timestamp 1677622389
transform -1 0 2552 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7344
timestamp 1677622389
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7345
timestamp 1677622389
transform 1 0 2560 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_48
timestamp 1677622389
transform -1 0 2600 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7346
timestamp 1677622389
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7347
timestamp 1677622389
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7348
timestamp 1677622389
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_454
timestamp 1677622389
transform 1 0 2624 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7349
timestamp 1677622389
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7351
timestamp 1677622389
transform 1 0 2648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7352
timestamp 1677622389
transform 1 0 2656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7353
timestamp 1677622389
transform 1 0 2664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7355
timestamp 1677622389
transform 1 0 2672 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_49
timestamp 1677622389
transform 1 0 2680 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7361
timestamp 1677622389
transform 1 0 2712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7362
timestamp 1677622389
transform 1 0 2720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7363
timestamp 1677622389
transform 1 0 2728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7364
timestamp 1677622389
transform 1 0 2736 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_50
timestamp 1677622389
transform 1 0 2744 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7365
timestamp 1677622389
transform 1 0 2776 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_456
timestamp 1677622389
transform 1 0 2784 0 -1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_73
timestamp 1677622389
transform -1 0 2824 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7366
timestamp 1677622389
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7367
timestamp 1677622389
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7368
timestamp 1677622389
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7371
timestamp 1677622389
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1677622389
transform -1 0 2888 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7372
timestamp 1677622389
transform 1 0 2888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7373
timestamp 1677622389
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7382
timestamp 1677622389
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_459
timestamp 1677622389
transform -1 0 2928 0 -1 1770
box -9 -3 26 105
use XNOR2X1  XNOR2X1_0
timestamp 1677622389
transform -1 0 2984 0 -1 1770
box -8 -3 64 105
use NAND2X1  NAND2X1_4
timestamp 1677622389
transform 1 0 2984 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7383
timestamp 1677622389
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_76
timestamp 1677622389
transform 1 0 3016 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7391
timestamp 1677622389
transform 1 0 3040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7392
timestamp 1677622389
transform 1 0 3048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7393
timestamp 1677622389
transform 1 0 3056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7394
timestamp 1677622389
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_461
timestamp 1677622389
transform 1 0 3072 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7395
timestamp 1677622389
transform 1 0 3088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7396
timestamp 1677622389
transform 1 0 3096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7397
timestamp 1677622389
transform 1 0 3104 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_77
timestamp 1677622389
transform 1 0 3112 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7398
timestamp 1677622389
transform 1 0 3136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7399
timestamp 1677622389
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7400
timestamp 1677622389
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_52
timestamp 1677622389
transform -1 0 3192 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7401
timestamp 1677622389
transform 1 0 3192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7403
timestamp 1677622389
transform 1 0 3200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7405
timestamp 1677622389
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7410
timestamp 1677622389
transform 1 0 3216 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_53
timestamp 1677622389
transform -1 0 3256 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7411
timestamp 1677622389
transform 1 0 3256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7413
timestamp 1677622389
transform 1 0 3264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7414
timestamp 1677622389
transform 1 0 3272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7415
timestamp 1677622389
transform 1 0 3280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7416
timestamp 1677622389
transform 1 0 3288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7417
timestamp 1677622389
transform 1 0 3296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7424
timestamp 1677622389
transform 1 0 3304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7425
timestamp 1677622389
transform 1 0 3312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7426
timestamp 1677622389
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_57
timestamp 1677622389
transform 1 0 3328 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7427
timestamp 1677622389
transform 1 0 3360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7428
timestamp 1677622389
transform 1 0 3368 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_463
timestamp 1677622389
transform -1 0 3392 0 -1 1770
box -9 -3 26 105
use OAI22X1  OAI22X1_266
timestamp 1677622389
transform 1 0 3392 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7429
timestamp 1677622389
transform 1 0 3432 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5624
timestamp 1677622389
transform 1 0 3452 0 1 1675
box -3 -3 3 3
use FILL  FILL_7431
timestamp 1677622389
transform 1 0 3440 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_464
timestamp 1677622389
transform -1 0 3464 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_465
timestamp 1677622389
transform -1 0 3480 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7432
timestamp 1677622389
transform 1 0 3480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7433
timestamp 1677622389
transform 1 0 3488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7454
timestamp 1677622389
transform 1 0 3496 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_50
timestamp 1677622389
transform 1 0 3504 0 -1 1770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_403
timestamp 1677622389
transform 1 0 3536 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7455
timestamp 1677622389
transform 1 0 3632 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_469
timestamp 1677622389
transform 1 0 3640 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7456
timestamp 1677622389
transform 1 0 3656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7457
timestamp 1677622389
transform 1 0 3664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7458
timestamp 1677622389
transform 1 0 3672 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_268
timestamp 1677622389
transform 1 0 3680 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7459
timestamp 1677622389
transform 1 0 3720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7460
timestamp 1677622389
transform 1 0 3728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7461
timestamp 1677622389
transform 1 0 3736 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_470
timestamp 1677622389
transform -1 0 3760 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7462
timestamp 1677622389
transform 1 0 3760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7463
timestamp 1677622389
transform 1 0 3768 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_269
timestamp 1677622389
transform 1 0 3776 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7464
timestamp 1677622389
transform 1 0 3816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7465
timestamp 1677622389
transform 1 0 3824 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_471
timestamp 1677622389
transform 1 0 3832 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7466
timestamp 1677622389
transform 1 0 3848 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_270
timestamp 1677622389
transform 1 0 3856 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_271
timestamp 1677622389
transform 1 0 3896 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7467
timestamp 1677622389
transform 1 0 3936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7468
timestamp 1677622389
transform 1 0 3944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7469
timestamp 1677622389
transform 1 0 3952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7470
timestamp 1677622389
transform 1 0 3960 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_472
timestamp 1677622389
transform -1 0 3984 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7471
timestamp 1677622389
transform 1 0 3984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7472
timestamp 1677622389
transform 1 0 3992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7473
timestamp 1677622389
transform 1 0 4000 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_404
timestamp 1677622389
transform 1 0 4008 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_473
timestamp 1677622389
transform -1 0 4120 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7474
timestamp 1677622389
transform 1 0 4120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7476
timestamp 1677622389
transform 1 0 4128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7488
timestamp 1677622389
transform 1 0 4136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7489
timestamp 1677622389
transform 1 0 4144 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_406
timestamp 1677622389
transform 1 0 4152 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7490
timestamp 1677622389
transform 1 0 4248 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_475
timestamp 1677622389
transform -1 0 4272 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7491
timestamp 1677622389
transform 1 0 4272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7492
timestamp 1677622389
transform 1 0 4280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7493
timestamp 1677622389
transform 1 0 4288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7494
timestamp 1677622389
transform 1 0 4296 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_273
timestamp 1677622389
transform 1 0 4304 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7495
timestamp 1677622389
transform 1 0 4344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7496
timestamp 1677622389
transform 1 0 4352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7497
timestamp 1677622389
transform 1 0 4360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7498
timestamp 1677622389
transform 1 0 4368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7500
timestamp 1677622389
transform 1 0 4376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7502
timestamp 1677622389
transform 1 0 4384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7504
timestamp 1677622389
transform 1 0 4392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7508
timestamp 1677622389
transform 1 0 4400 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_477
timestamp 1677622389
transform -1 0 4424 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7509
timestamp 1677622389
transform 1 0 4424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7510
timestamp 1677622389
transform 1 0 4432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7512
timestamp 1677622389
transform 1 0 4440 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_274
timestamp 1677622389
transform 1 0 4448 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7514
timestamp 1677622389
transform 1 0 4488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7515
timestamp 1677622389
transform 1 0 4496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7516
timestamp 1677622389
transform 1 0 4504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7517
timestamp 1677622389
transform 1 0 4512 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_478
timestamp 1677622389
transform -1 0 4536 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7518
timestamp 1677622389
transform 1 0 4536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7519
timestamp 1677622389
transform 1 0 4544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7521
timestamp 1677622389
transform 1 0 4552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7523
timestamp 1677622389
transform 1 0 4560 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_276
timestamp 1677622389
transform 1 0 4568 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7525
timestamp 1677622389
transform 1 0 4608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7527
timestamp 1677622389
transform 1 0 4616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7528
timestamp 1677622389
transform 1 0 4624 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_278
timestamp 1677622389
transform 1 0 4632 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7529
timestamp 1677622389
transform 1 0 4672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7530
timestamp 1677622389
transform 1 0 4680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7531
timestamp 1677622389
transform 1 0 4688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7532
timestamp 1677622389
transform 1 0 4696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7533
timestamp 1677622389
transform 1 0 4704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7534
timestamp 1677622389
transform 1 0 4712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7535
timestamp 1677622389
transform 1 0 4720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7536
timestamp 1677622389
transform 1 0 4728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7537
timestamp 1677622389
transform 1 0 4736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7538
timestamp 1677622389
transform 1 0 4744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7539
timestamp 1677622389
transform 1 0 4752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7540
timestamp 1677622389
transform 1 0 4760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7541
timestamp 1677622389
transform 1 0 4768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7542
timestamp 1677622389
transform 1 0 4776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7543
timestamp 1677622389
transform 1 0 4784 0 -1 1770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_61
timestamp 1677622389
transform 1 0 4843 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_6383
timestamp 1677622389
transform 1 0 116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1677622389
transform 1 0 148 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5650
timestamp 1677622389
transform 1 0 188 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1677622389
transform 1 0 228 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1677622389
transform 1 0 164 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1677622389
transform 1 0 180 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1677622389
transform 1 0 196 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6385
timestamp 1677622389
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1677622389
transform 1 0 180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1677622389
transform 1 0 196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1677622389
transform 1 0 164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1677622389
transform 1 0 172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1677622389
transform 1 0 188 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5723
timestamp 1677622389
transform 1 0 212 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6388
timestamp 1677622389
transform 1 0 244 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5724
timestamp 1677622389
transform 1 0 284 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6487
timestamp 1677622389
transform 1 0 212 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5691
timestamp 1677622389
transform 1 0 308 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6389
timestamp 1677622389
transform 1 0 300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1677622389
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5747
timestamp 1677622389
transform 1 0 300 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1677622389
transform 1 0 324 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6391
timestamp 1677622389
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1677622389
transform 1 0 324 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5748
timestamp 1677622389
transform 1 0 332 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1677622389
transform 1 0 444 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6392
timestamp 1677622389
transform 1 0 356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1677622389
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1677622389
transform 1 0 340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1677622389
transform 1 0 348 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5726
timestamp 1677622389
transform 1 0 380 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6394
timestamp 1677622389
transform 1 0 420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1677622389
transform 1 0 444 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5768
timestamp 1677622389
transform 1 0 444 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1677622389
transform 1 0 508 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1677622389
transform 1 0 468 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6395
timestamp 1677622389
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1677622389
transform 1 0 548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1677622389
transform 1 0 468 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5769
timestamp 1677622389
transform 1 0 468 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1677622389
transform 1 0 548 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1677622389
transform 1 0 572 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6493
timestamp 1677622389
transform 1 0 596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1677622389
transform 1 0 612 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5771
timestamp 1677622389
transform 1 0 612 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1677622389
transform 1 0 628 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6397
timestamp 1677622389
transform 1 0 620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1677622389
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1677622389
transform 1 0 692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1677622389
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5749
timestamp 1677622389
transform 1 0 692 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6496
timestamp 1677622389
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1677622389
transform 1 0 708 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5772
timestamp 1677622389
transform 1 0 676 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1677622389
transform 1 0 684 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1677622389
transform 1 0 708 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1677622389
transform 1 0 732 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1677622389
transform 1 0 836 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6400
timestamp 1677622389
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1677622389
transform 1 0 820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1677622389
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5751
timestamp 1677622389
transform 1 0 804 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1677622389
transform 1 0 836 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6586
timestamp 1677622389
transform 1 0 844 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5789
timestamp 1677622389
transform 1 0 844 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1677622389
transform 1 0 860 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6498
timestamp 1677622389
transform 1 0 860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1677622389
transform 1 0 964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1677622389
transform 1 0 956 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1677622389
transform 1 0 1012 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5729
timestamp 1677622389
transform 1 0 1020 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6500
timestamp 1677622389
transform 1 0 1036 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5636
timestamp 1677622389
transform 1 0 1100 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1677622389
transform 1 0 1100 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6404
timestamp 1677622389
transform 1 0 1092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1677622389
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1677622389
transform 1 0 1116 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5753
timestamp 1677622389
transform 1 0 1092 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6501
timestamp 1677622389
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5790
timestamp 1677622389
transform 1 0 1084 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6502
timestamp 1677622389
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1677622389
transform 1 0 1180 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5670
timestamp 1677622389
transform 1 0 1196 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1677622389
transform 1 0 1252 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1677622389
transform 1 0 1236 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6408
timestamp 1677622389
transform 1 0 1236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1677622389
transform 1 0 1260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1677622389
transform 1 0 1228 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5754
timestamp 1677622389
transform 1 0 1236 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6504
timestamp 1677622389
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5696
timestamp 1677622389
transform 1 0 1308 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6505
timestamp 1677622389
transform 1 0 1300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1677622389
transform 1 0 1324 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5671
timestamp 1677622389
transform 1 0 1356 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1677622389
transform 1 0 1372 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1677622389
transform 1 0 1348 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6410
timestamp 1677622389
transform 1 0 1356 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5730
timestamp 1677622389
transform 1 0 1364 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6411
timestamp 1677622389
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1677622389
transform 1 0 1364 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5791
timestamp 1677622389
transform 1 0 1348 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1677622389
transform 1 0 1420 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1677622389
transform 1 0 1436 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1677622389
transform 1 0 1492 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6412
timestamp 1677622389
transform 1 0 1436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1677622389
transform 1 0 1492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1677622389
transform 1 0 1516 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5699
timestamp 1677622389
transform 1 0 1532 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6414
timestamp 1677622389
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1677622389
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5792
timestamp 1677622389
transform 1 0 1636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1677622389
transform 1 0 1692 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6415
timestamp 1677622389
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1677622389
transform 1 0 1732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1677622389
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1677622389
transform 1 0 1716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1677622389
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1677622389
transform 1 0 1748 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5793
timestamp 1677622389
transform 1 0 1740 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1677622389
transform 1 0 1764 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6418
timestamp 1677622389
transform 1 0 1764 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5639
timestamp 1677622389
transform 1 0 1836 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6419
timestamp 1677622389
transform 1 0 1844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1677622389
transform 1 0 1868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1677622389
transform 1 0 1892 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5700
timestamp 1677622389
transform 1 0 1940 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6420
timestamp 1677622389
transform 1 0 1924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1677622389
transform 1 0 1940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1677622389
transform 1 0 1956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1677622389
transform 1 0 1932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1677622389
transform 1 0 1948 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5654
timestamp 1677622389
transform 1 0 1996 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6517
timestamp 1677622389
transform 1 0 1996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1677622389
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1677622389
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5701
timestamp 1677622389
transform 1 0 2076 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6519
timestamp 1677622389
transform 1 0 2076 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5640
timestamp 1677622389
transform 1 0 2100 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1677622389
transform 1 0 2092 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6424
timestamp 1677622389
transform 1 0 2100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1677622389
transform 1 0 2132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1677622389
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5794
timestamp 1677622389
transform 1 0 2140 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1677622389
transform 1 0 2180 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6426
timestamp 1677622389
transform 1 0 2204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1677622389
transform 1 0 2236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1677622389
transform 1 0 2284 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5796
timestamp 1677622389
transform 1 0 2284 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1677622389
transform 1 0 2388 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1677622389
transform 1 0 2388 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6428
timestamp 1677622389
transform 1 0 2308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1677622389
transform 1 0 2364 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5755
timestamp 1677622389
transform 1 0 2364 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6522
timestamp 1677622389
transform 1 0 2388 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5774
timestamp 1677622389
transform 1 0 2340 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1677622389
transform 1 0 2388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1677622389
transform 1 0 2412 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6430
timestamp 1677622389
transform 1 0 2412 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5704
timestamp 1677622389
transform 1 0 2436 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1677622389
transform 1 0 2468 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6431
timestamp 1677622389
transform 1 0 2468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1677622389
transform 1 0 2500 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5798
timestamp 1677622389
transform 1 0 2500 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1677622389
transform 1 0 2532 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6524
timestamp 1677622389
transform 1 0 2524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1677622389
transform 1 0 2540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1677622389
transform 1 0 2548 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5756
timestamp 1677622389
transform 1 0 2548 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6525
timestamp 1677622389
transform 1 0 2556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1677622389
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1677622389
transform 1 0 2660 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5757
timestamp 1677622389
transform 1 0 2644 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6526
timestamp 1677622389
transform 1 0 2684 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5799
timestamp 1677622389
transform 1 0 2684 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6371
timestamp 1677622389
transform 1 0 2700 0 1 1655
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1677622389
transform 1 0 2716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1677622389
transform 1 0 2732 0 1 1655
box -2 -2 2 2
use M3_M2  M3_M2_5775
timestamp 1677622389
transform 1 0 2748 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1677622389
transform 1 0 2748 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1677622389
transform 1 0 2780 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6436
timestamp 1677622389
transform 1 0 2804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1677622389
transform 1 0 2852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1677622389
transform 1 0 2868 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1677622389
transform 1 0 2900 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1677622389
transform 1 0 2908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1677622389
transform 1 0 2932 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1677622389
transform 1 0 3028 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1677622389
transform 1 0 3012 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5731
timestamp 1677622389
transform 1 0 3012 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6379
timestamp 1677622389
transform 1 0 3036 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1677622389
transform 1 0 3020 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5732
timestamp 1677622389
transform 1 0 3044 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6529
timestamp 1677622389
transform 1 0 3044 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5641
timestamp 1677622389
transform 1 0 3108 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1677622389
transform 1 0 3140 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1677622389
transform 1 0 3100 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6439
timestamp 1677622389
transform 1 0 3100 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5677
timestamp 1677622389
transform 1 0 3132 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6440
timestamp 1677622389
transform 1 0 3204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1677622389
transform 1 0 3116 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1677622389
transform 1 0 3236 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5678
timestamp 1677622389
transform 1 0 3244 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6441
timestamp 1677622389
transform 1 0 3236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1677622389
transform 1 0 3252 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1677622389
transform 1 0 3244 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5707
timestamp 1677622389
transform 1 0 3260 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6381
timestamp 1677622389
transform 1 0 3276 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1677622389
transform 1 0 3260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1677622389
transform 1 0 3284 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5758
timestamp 1677622389
transform 1 0 3268 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6444
timestamp 1677622389
transform 1 0 3300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1677622389
transform 1 0 3292 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5776
timestamp 1677622389
transform 1 0 3276 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1677622389
transform 1 0 3300 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1677622389
transform 1 0 3308 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1677622389
transform 1 0 3332 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1677622389
transform 1 0 3340 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1677622389
transform 1 0 3356 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6445
timestamp 1677622389
transform 1 0 3364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1677622389
transform 1 0 3332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1677622389
transform 1 0 3348 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5777
timestamp 1677622389
transform 1 0 3324 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1677622389
transform 1 0 3324 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1677622389
transform 1 0 3364 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6534
timestamp 1677622389
transform 1 0 3372 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5679
timestamp 1677622389
transform 1 0 3396 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1677622389
transform 1 0 3412 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1677622389
transform 1 0 3404 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6535
timestamp 1677622389
transform 1 0 3396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1677622389
transform 1 0 3404 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5803
timestamp 1677622389
transform 1 0 3404 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6446
timestamp 1677622389
transform 1 0 3420 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5643
timestamp 1677622389
transform 1 0 3444 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1677622389
transform 1 0 3492 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1677622389
transform 1 0 3508 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1677622389
transform 1 0 3460 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1677622389
transform 1 0 3516 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1677622389
transform 1 0 3532 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1677622389
transform 1 0 3580 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1677622389
transform 1 0 3452 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6536
timestamp 1677622389
transform 1 0 3436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1677622389
transform 1 0 3452 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5680
timestamp 1677622389
transform 1 0 3476 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1677622389
transform 1 0 3572 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1677622389
transform 1 0 3564 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6448
timestamp 1677622389
transform 1 0 3556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1677622389
transform 1 0 3564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1677622389
transform 1 0 3572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1677622389
transform 1 0 3580 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5761
timestamp 1677622389
transform 1 0 3468 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6537
timestamp 1677622389
transform 1 0 3572 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1677622389
transform 1 0 3468 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5662
timestamp 1677622389
transform 1 0 3620 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6452
timestamp 1677622389
transform 1 0 3604 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5735
timestamp 1677622389
transform 1 0 3612 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6453
timestamp 1677622389
transform 1 0 3620 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5736
timestamp 1677622389
transform 1 0 3636 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6538
timestamp 1677622389
transform 1 0 3612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1677622389
transform 1 0 3628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1677622389
transform 1 0 3644 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5778
timestamp 1677622389
transform 1 0 3612 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1677622389
transform 1 0 3644 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1677622389
transform 1 0 3668 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6541
timestamp 1677622389
transform 1 0 3676 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5779
timestamp 1677622389
transform 1 0 3684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1677622389
transform 1 0 3692 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1677622389
transform 1 0 3716 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1677622389
transform 1 0 3708 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6454
timestamp 1677622389
transform 1 0 3716 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5738
timestamp 1677622389
transform 1 0 3724 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6455
timestamp 1677622389
transform 1 0 3732 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5712
timestamp 1677622389
transform 1 0 3748 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6456
timestamp 1677622389
transform 1 0 3748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1677622389
transform 1 0 3708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1677622389
transform 1 0 3724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1677622389
transform 1 0 3740 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5780
timestamp 1677622389
transform 1 0 3708 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1677622389
transform 1 0 3748 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6545
timestamp 1677622389
transform 1 0 3756 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5645
timestamp 1677622389
transform 1 0 3812 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1677622389
transform 1 0 3804 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1677622389
transform 1 0 3796 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6457
timestamp 1677622389
transform 1 0 3804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1677622389
transform 1 0 3796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1677622389
transform 1 0 3812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1677622389
transform 1 0 3820 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5781
timestamp 1677622389
transform 1 0 3820 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1677622389
transform 1 0 3860 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1677622389
transform 1 0 3868 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6458
timestamp 1677622389
transform 1 0 3852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1677622389
transform 1 0 3868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1677622389
transform 1 0 3860 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5763
timestamp 1677622389
transform 1 0 3868 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1677622389
transform 1 0 3884 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1677622389
transform 1 0 3884 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6550
timestamp 1677622389
transform 1 0 3876 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5646
timestamp 1677622389
transform 1 0 3900 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6382
timestamp 1677622389
transform 1 0 3908 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1677622389
transform 1 0 3900 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5713
timestamp 1677622389
transform 1 0 3924 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6461
timestamp 1677622389
transform 1 0 3924 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5684
timestamp 1677622389
transform 1 0 3940 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1677622389
transform 1 0 3940 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1677622389
transform 1 0 3956 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6462
timestamp 1677622389
transform 1 0 3964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1677622389
transform 1 0 3932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1677622389
transform 1 0 3940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1677622389
transform 1 0 3956 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5715
timestamp 1677622389
transform 1 0 3980 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6463
timestamp 1677622389
transform 1 0 3980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1677622389
transform 1 0 4028 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5741
timestamp 1677622389
transform 1 0 4036 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6554
timestamp 1677622389
transform 1 0 3996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1677622389
transform 1 0 4004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1677622389
transform 1 0 4020 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1677622389
transform 1 0 4036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1677622389
transform 1 0 4044 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5782
timestamp 1677622389
transform 1 0 3996 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1677622389
transform 1 0 4060 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1677622389
transform 1 0 4076 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1677622389
transform 1 0 4100 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1677622389
transform 1 0 4084 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1677622389
transform 1 0 4116 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6465
timestamp 1677622389
transform 1 0 4060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1677622389
transform 1 0 4076 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5742
timestamp 1677622389
transform 1 0 4092 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6467
timestamp 1677622389
transform 1 0 4100 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5648
timestamp 1677622389
transform 1 0 4132 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6559
timestamp 1677622389
transform 1 0 4068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1677622389
transform 1 0 4084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1677622389
transform 1 0 4092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1677622389
transform 1 0 4108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1677622389
transform 1 0 4124 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5783
timestamp 1677622389
transform 1 0 4044 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1677622389
transform 1 0 4004 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1677622389
transform 1 0 4028 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1677622389
transform 1 0 4124 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1677622389
transform 1 0 4148 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1677622389
transform 1 0 4156 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6468
timestamp 1677622389
transform 1 0 4156 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5743
timestamp 1677622389
transform 1 0 4164 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6469
timestamp 1677622389
transform 1 0 4172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1677622389
transform 1 0 4148 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1677622389
transform 1 0 4164 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5764
timestamp 1677622389
transform 1 0 4172 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1677622389
transform 1 0 4148 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1677622389
transform 1 0 4196 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6566
timestamp 1677622389
transform 1 0 4212 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5631
timestamp 1677622389
transform 1 0 4228 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1677622389
transform 1 0 4244 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6470
timestamp 1677622389
transform 1 0 4228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1677622389
transform 1 0 4244 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5686
timestamp 1677622389
transform 1 0 4260 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6472
timestamp 1677622389
transform 1 0 4260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1677622389
transform 1 0 4236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1677622389
transform 1 0 4252 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5785
timestamp 1677622389
transform 1 0 4252 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1677622389
transform 1 0 4308 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6473
timestamp 1677622389
transform 1 0 4308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1677622389
transform 1 0 4284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1677622389
transform 1 0 4300 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5765
timestamp 1677622389
transform 1 0 4308 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1677622389
transform 1 0 4324 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6474
timestamp 1677622389
transform 1 0 4324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1677622389
transform 1 0 4316 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5786
timestamp 1677622389
transform 1 0 4284 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6572
timestamp 1677622389
transform 1 0 4332 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5787
timestamp 1677622389
transform 1 0 4332 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1677622389
transform 1 0 4388 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6475
timestamp 1677622389
transform 1 0 4388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1677622389
transform 1 0 4364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1677622389
transform 1 0 4380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1677622389
transform 1 0 4396 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5668
timestamp 1677622389
transform 1 0 4420 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6476
timestamp 1677622389
transform 1 0 4420 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5633
timestamp 1677622389
transform 1 0 4452 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6477
timestamp 1677622389
transform 1 0 4452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1677622389
transform 1 0 4428 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5766
timestamp 1677622389
transform 1 0 4436 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6577
timestamp 1677622389
transform 1 0 4444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1677622389
transform 1 0 4460 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5634
timestamp 1677622389
transform 1 0 4500 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1677622389
transform 1 0 4532 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1677622389
transform 1 0 4516 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6478
timestamp 1677622389
transform 1 0 4516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1677622389
transform 1 0 4532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1677622389
transform 1 0 4524 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5767
timestamp 1677622389
transform 1 0 4532 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6580
timestamp 1677622389
transform 1 0 4540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1677622389
transform 1 0 4564 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5720
timestamp 1677622389
transform 1 0 4604 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1677622389
transform 1 0 4580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6480
timestamp 1677622389
transform 1 0 4604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1677622389
transform 1 0 4580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1677622389
transform 1 0 4596 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5669
timestamp 1677622389
transform 1 0 4628 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1677622389
transform 1 0 4620 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1677622389
transform 1 0 4668 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1677622389
transform 1 0 4676 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6591
timestamp 1677622389
transform 1 0 4676 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5722
timestamp 1677622389
transform 1 0 4780 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6481
timestamp 1677622389
transform 1 0 4732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1677622389
transform 1 0 4772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1677622389
transform 1 0 4780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1677622389
transform 1 0 4692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1677622389
transform 1 0 4788 0 1 1605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_62
timestamp 1677622389
transform 1 0 48 0 1 1570
box -10 -3 10 3
use FILL  FILL_7544
timestamp 1677622389
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_7545
timestamp 1677622389
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_7546
timestamp 1677622389
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_7547
timestamp 1677622389
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_7548
timestamp 1677622389
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_7549
timestamp 1677622389
transform 1 0 112 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_481
timestamp 1677622389
transform -1 0 136 0 1 1570
box -9 -3 26 105
use FILL  FILL_7550
timestamp 1677622389
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7551
timestamp 1677622389
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_7552
timestamp 1677622389
transform 1 0 152 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_280
timestamp 1677622389
transform -1 0 200 0 1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_409
timestamp 1677622389
transform 1 0 200 0 1 1570
box -8 -3 104 105
use FILL  FILL_7553
timestamp 1677622389
transform 1 0 296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7554
timestamp 1677622389
transform 1 0 304 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_281
timestamp 1677622389
transform 1 0 312 0 1 1570
box -8 -3 46 105
use FILL  FILL_7559
timestamp 1677622389
transform 1 0 352 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5810
timestamp 1677622389
transform 1 0 388 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_412
timestamp 1677622389
transform -1 0 456 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_413
timestamp 1677622389
transform 1 0 456 0 1 1570
box -8 -3 104 105
use FILL  FILL_7560
timestamp 1677622389
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7573
timestamp 1677622389
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7575
timestamp 1677622389
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_7577
timestamp 1677622389
transform 1 0 576 0 1 1570
box -8 -3 16 105
use FILL  FILL_7579
timestamp 1677622389
transform 1 0 584 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_485
timestamp 1677622389
transform 1 0 592 0 1 1570
box -9 -3 26 105
use FILL  FILL_7580
timestamp 1677622389
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_7581
timestamp 1677622389
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7582
timestamp 1677622389
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7583
timestamp 1677622389
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_7584
timestamp 1677622389
transform 1 0 640 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5811
timestamp 1677622389
transform 1 0 660 0 1 1575
box -3 -3 3 3
use FILL  FILL_7585
timestamp 1677622389
transform 1 0 648 0 1 1570
box -8 -3 16 105
use FILL  FILL_7586
timestamp 1677622389
transform 1 0 656 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_280
timestamp 1677622389
transform 1 0 664 0 1 1570
box -8 -3 46 105
use FILL  FILL_7587
timestamp 1677622389
transform 1 0 704 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5812
timestamp 1677622389
transform 1 0 724 0 1 1575
box -3 -3 3 3
use FILL  FILL_7588
timestamp 1677622389
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_7589
timestamp 1677622389
transform 1 0 720 0 1 1570
box -8 -3 16 105
use FILL  FILL_7590
timestamp 1677622389
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_7591
timestamp 1677622389
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_7592
timestamp 1677622389
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7597
timestamp 1677622389
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7599
timestamp 1677622389
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_7601
timestamp 1677622389
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_7603
timestamp 1677622389
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_7605
timestamp 1677622389
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7606
timestamp 1677622389
transform 1 0 792 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_284
timestamp 1677622389
transform -1 0 840 0 1 1570
box -8 -3 46 105
use FILL  FILL_7607
timestamp 1677622389
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_7611
timestamp 1677622389
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_7613
timestamp 1677622389
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_7615
timestamp 1677622389
transform 1 0 864 0 1 1570
box -8 -3 16 105
use FILL  FILL_7617
timestamp 1677622389
transform 1 0 872 0 1 1570
box -8 -3 16 105
use FILL  FILL_7618
timestamp 1677622389
transform 1 0 880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7619
timestamp 1677622389
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_7620
timestamp 1677622389
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_7622
timestamp 1677622389
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_7624
timestamp 1677622389
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_7626
timestamp 1677622389
transform 1 0 920 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5813
timestamp 1677622389
transform 1 0 956 0 1 1575
box -3 -3 3 3
use NOR2X1  NOR2X1_78
timestamp 1677622389
transform 1 0 928 0 1 1570
box -8 -3 32 105
use FILL  FILL_7628
timestamp 1677622389
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7629
timestamp 1677622389
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7630
timestamp 1677622389
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_7631
timestamp 1677622389
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7632
timestamp 1677622389
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7633
timestamp 1677622389
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_7634
timestamp 1677622389
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_79
timestamp 1677622389
transform 1 0 1008 0 1 1570
box -8 -3 32 105
use FILL  FILL_7635
timestamp 1677622389
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_7638
timestamp 1677622389
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_7640
timestamp 1677622389
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_7641
timestamp 1677622389
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_7642
timestamp 1677622389
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_7643
timestamp 1677622389
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_7646
timestamp 1677622389
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7648
timestamp 1677622389
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_286
timestamp 1677622389
transform 1 0 1096 0 1 1570
box -8 -3 46 105
use FILL  FILL_7650
timestamp 1677622389
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7651
timestamp 1677622389
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_7652
timestamp 1677622389
transform 1 0 1152 0 1 1570
box -8 -3 16 105
use FILL  FILL_7653
timestamp 1677622389
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_7654
timestamp 1677622389
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_7655
timestamp 1677622389
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7662
timestamp 1677622389
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7664
timestamp 1677622389
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5814
timestamp 1677622389
transform 1 0 1212 0 1 1575
box -3 -3 3 3
use FILL  FILL_7666
timestamp 1677622389
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_7668
timestamp 1677622389
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_7670
timestamp 1677622389
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5815
timestamp 1677622389
transform 1 0 1244 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_282
timestamp 1677622389
transform -1 0 1264 0 1 1570
box -8 -3 46 105
use FILL  FILL_7671
timestamp 1677622389
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_7672
timestamp 1677622389
transform 1 0 1272 0 1 1570
box -8 -3 16 105
use FILL  FILL_7673
timestamp 1677622389
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_7674
timestamp 1677622389
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_7680
timestamp 1677622389
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7682
timestamp 1677622389
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7684
timestamp 1677622389
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_7686
timestamp 1677622389
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_7688
timestamp 1677622389
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use FILL  FILL_7689
timestamp 1677622389
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_283
timestamp 1677622389
transform -1 0 1384 0 1 1570
box -8 -3 46 105
use FILL  FILL_7690
timestamp 1677622389
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_7691
timestamp 1677622389
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_7692
timestamp 1677622389
transform 1 0 1400 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5816
timestamp 1677622389
transform 1 0 1420 0 1 1575
box -3 -3 3 3
use FILL  FILL_7693
timestamp 1677622389
transform 1 0 1408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7694
timestamp 1677622389
transform 1 0 1416 0 1 1570
box -8 -3 16 105
use FILL  FILL_7695
timestamp 1677622389
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5817
timestamp 1677622389
transform 1 0 1516 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_416
timestamp 1677622389
transform -1 0 1528 0 1 1570
box -8 -3 104 105
use FILL  FILL_7696
timestamp 1677622389
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_7706
timestamp 1677622389
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5818
timestamp 1677622389
transform 1 0 1572 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_487
timestamp 1677622389
transform 1 0 1544 0 1 1570
box -9 -3 26 105
use FILL  FILL_7708
timestamp 1677622389
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7709
timestamp 1677622389
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_7710
timestamp 1677622389
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_7711
timestamp 1677622389
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_7712
timestamp 1677622389
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_7713
timestamp 1677622389
transform 1 0 1600 0 1 1570
box -8 -3 16 105
use FILL  FILL_7714
timestamp 1677622389
transform 1 0 1608 0 1 1570
box -8 -3 16 105
use FILL  FILL_7715
timestamp 1677622389
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7716
timestamp 1677622389
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7717
timestamp 1677622389
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_7718
timestamp 1677622389
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_7719
timestamp 1677622389
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_7720
timestamp 1677622389
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_7721
timestamp 1677622389
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7724
timestamp 1677622389
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_7726
timestamp 1677622389
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_7728
timestamp 1677622389
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_7730
timestamp 1677622389
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_7732
timestamp 1677622389
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_290
timestamp 1677622389
transform 1 0 1712 0 1 1570
box -8 -3 46 105
use FILL  FILL_7734
timestamp 1677622389
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7735
timestamp 1677622389
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_7736
timestamp 1677622389
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_7737
timestamp 1677622389
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_419
timestamp 1677622389
transform -1 0 1880 0 1 1570
box -8 -3 104 105
use FILL  FILL_7738
timestamp 1677622389
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7739
timestamp 1677622389
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use FILL  FILL_7740
timestamp 1677622389
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_7741
timestamp 1677622389
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_284
timestamp 1677622389
transform -1 0 1952 0 1 1570
box -8 -3 46 105
use FILL  FILL_7742
timestamp 1677622389
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7743
timestamp 1677622389
transform 1 0 1960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7744
timestamp 1677622389
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_94
timestamp 1677622389
transform 1 0 1976 0 1 1570
box -5 -3 28 105
use FILL  FILL_7745
timestamp 1677622389
transform 1 0 2000 0 1 1570
box -8 -3 16 105
use FILL  FILL_7766
timestamp 1677622389
transform 1 0 2008 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_95
timestamp 1677622389
transform -1 0 2040 0 1 1570
box -5 -3 28 105
use FILL  FILL_7767
timestamp 1677622389
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use FILL  FILL_7773
timestamp 1677622389
transform 1 0 2048 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_96
timestamp 1677622389
transform 1 0 2056 0 1 1570
box -5 -3 28 105
use FILL  FILL_7775
timestamp 1677622389
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7778
timestamp 1677622389
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_420
timestamp 1677622389
transform -1 0 2192 0 1 1570
box -8 -3 104 105
use FILL  FILL_7779
timestamp 1677622389
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5819
timestamp 1677622389
transform 1 0 2276 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_421
timestamp 1677622389
transform -1 0 2296 0 1 1570
box -8 -3 104 105
use FILL  FILL_7780
timestamp 1677622389
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5820
timestamp 1677622389
transform 1 0 2316 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_422
timestamp 1677622389
transform -1 0 2400 0 1 1570
box -8 -3 104 105
use FILL  FILL_7781
timestamp 1677622389
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_7782
timestamp 1677622389
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_423
timestamp 1677622389
transform -1 0 2512 0 1 1570
box -8 -3 104 105
use FILL  FILL_7783
timestamp 1677622389
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use FILL  FILL_7784
timestamp 1677622389
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_491
timestamp 1677622389
transform 1 0 2528 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_492
timestamp 1677622389
transform -1 0 2560 0 1 1570
box -9 -3 26 105
use FILL  FILL_7806
timestamp 1677622389
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7807
timestamp 1677622389
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_7808
timestamp 1677622389
transform 1 0 2576 0 1 1570
box -8 -3 16 105
use FILL  FILL_7809
timestamp 1677622389
transform 1 0 2584 0 1 1570
box -8 -3 16 105
use FILL  FILL_7810
timestamp 1677622389
transform 1 0 2592 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_426
timestamp 1677622389
transform -1 0 2696 0 1 1570
box -8 -3 104 105
use FILL  FILL_7811
timestamp 1677622389
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use FILL  FILL_7812
timestamp 1677622389
transform 1 0 2704 0 1 1570
box -8 -3 16 105
use FILL  FILL_7813
timestamp 1677622389
transform 1 0 2712 0 1 1570
box -8 -3 16 105
use FILL  FILL_7814
timestamp 1677622389
transform 1 0 2720 0 1 1570
box -8 -3 16 105
use FILL  FILL_7815
timestamp 1677622389
transform 1 0 2728 0 1 1570
box -8 -3 16 105
use FILL  FILL_7816
timestamp 1677622389
transform 1 0 2736 0 1 1570
box -8 -3 16 105
use FILL  FILL_7817
timestamp 1677622389
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7818
timestamp 1677622389
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7819
timestamp 1677622389
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_7820
timestamp 1677622389
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_7821
timestamp 1677622389
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use FILL  FILL_7822
timestamp 1677622389
transform 1 0 2784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7823
timestamp 1677622389
transform 1 0 2792 0 1 1570
box -8 -3 16 105
use FILL  FILL_7831
timestamp 1677622389
transform 1 0 2800 0 1 1570
box -8 -3 16 105
use FILL  FILL_7833
timestamp 1677622389
transform 1 0 2808 0 1 1570
box -8 -3 16 105
use FILL  FILL_7835
timestamp 1677622389
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_80
timestamp 1677622389
transform -1 0 2848 0 1 1570
box -8 -3 32 105
use INVX2  INVX2_493
timestamp 1677622389
transform 1 0 2848 0 1 1570
box -9 -3 26 105
use FILL  FILL_7836
timestamp 1677622389
transform 1 0 2864 0 1 1570
box -8 -3 16 105
use FILL  FILL_7844
timestamp 1677622389
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_7846
timestamp 1677622389
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7848
timestamp 1677622389
transform 1 0 2888 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_59
timestamp 1677622389
transform 1 0 2896 0 1 1570
box -8 -3 40 105
use FILL  FILL_7850
timestamp 1677622389
transform 1 0 2928 0 1 1570
box -8 -3 16 105
use FILL  FILL_7852
timestamp 1677622389
transform 1 0 2936 0 1 1570
box -8 -3 16 105
use FILL  FILL_7854
timestamp 1677622389
transform 1 0 2944 0 1 1570
box -8 -3 16 105
use FILL  FILL_7856
timestamp 1677622389
transform 1 0 2952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7858
timestamp 1677622389
transform 1 0 2960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7860
timestamp 1677622389
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_7862
timestamp 1677622389
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7864
timestamp 1677622389
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7866
timestamp 1677622389
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use FILL  FILL_7867
timestamp 1677622389
transform 1 0 3000 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_60
timestamp 1677622389
transform 1 0 3008 0 1 1570
box -8 -3 40 105
use FILL  FILL_7868
timestamp 1677622389
transform 1 0 3040 0 1 1570
box -8 -3 16 105
use FILL  FILL_7870
timestamp 1677622389
transform 1 0 3048 0 1 1570
box -8 -3 16 105
use FILL  FILL_7872
timestamp 1677622389
transform 1 0 3056 0 1 1570
box -8 -3 16 105
use FILL  FILL_7874
timestamp 1677622389
transform 1 0 3064 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_495
timestamp 1677622389
transform 1 0 3072 0 1 1570
box -9 -3 26 105
use FILL  FILL_7876
timestamp 1677622389
transform 1 0 3088 0 1 1570
box -8 -3 16 105
use FILL  FILL_7877
timestamp 1677622389
transform 1 0 3096 0 1 1570
box -8 -3 16 105
use FAX1  FAX1_1
timestamp 1677622389
transform -1 0 3224 0 1 1570
box -5 -3 126 105
use FILL  FILL_7878
timestamp 1677622389
transform 1 0 3224 0 1 1570
box -8 -3 16 105
use FILL  FILL_7879
timestamp 1677622389
transform 1 0 3232 0 1 1570
box -8 -3 16 105
use FILL  FILL_7880
timestamp 1677622389
transform 1 0 3240 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_61
timestamp 1677622389
transform 1 0 3248 0 1 1570
box -8 -3 40 105
use INVX2  INVX2_496
timestamp 1677622389
transform -1 0 3296 0 1 1570
box -9 -3 26 105
use FILL  FILL_7881
timestamp 1677622389
transform 1 0 3296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7882
timestamp 1677622389
transform 1 0 3304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7894
timestamp 1677622389
transform 1 0 3312 0 1 1570
box -8 -3 16 105
use FILL  FILL_7896
timestamp 1677622389
transform 1 0 3320 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1677622389
transform -1 0 3360 0 1 1570
box -7 -3 39 105
use FILL  FILL_7897
timestamp 1677622389
transform 1 0 3360 0 1 1570
box -8 -3 16 105
use FILL  FILL_7898
timestamp 1677622389
transform 1 0 3368 0 1 1570
box -8 -3 16 105
use FILL  FILL_7899
timestamp 1677622389
transform 1 0 3376 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_497
timestamp 1677622389
transform -1 0 3400 0 1 1570
box -9 -3 26 105
use FILL  FILL_7900
timestamp 1677622389
transform 1 0 3400 0 1 1570
box -8 -3 16 105
use FILL  FILL_7907
timestamp 1677622389
transform 1 0 3408 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1677622389
transform -1 0 3448 0 1 1570
box -7 -3 39 105
use FILL  FILL_7908
timestamp 1677622389
transform 1 0 3448 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5821
timestamp 1677622389
transform 1 0 3564 0 1 1575
box -3 -3 3 3
use FAX1  FAX1_2
timestamp 1677622389
transform -1 0 3576 0 1 1570
box -5 -3 126 105
use INVX2  INVX2_498
timestamp 1677622389
transform 1 0 3576 0 1 1570
box -9 -3 26 105
use FILL  FILL_7915
timestamp 1677622389
transform 1 0 3592 0 1 1570
box -8 -3 16 105
use FILL  FILL_7916
timestamp 1677622389
transform 1 0 3600 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_286
timestamp 1677622389
transform -1 0 3648 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_499
timestamp 1677622389
transform -1 0 3664 0 1 1570
box -9 -3 26 105
use FILL  FILL_7917
timestamp 1677622389
transform 1 0 3664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7918
timestamp 1677622389
transform 1 0 3672 0 1 1570
box -8 -3 16 105
use FILL  FILL_7919
timestamp 1677622389
transform 1 0 3680 0 1 1570
box -8 -3 16 105
use FILL  FILL_7922
timestamp 1677622389
transform 1 0 3688 0 1 1570
box -8 -3 16 105
use FILL  FILL_7924
timestamp 1677622389
transform 1 0 3696 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_287
timestamp 1677622389
transform 1 0 3704 0 1 1570
box -8 -3 46 105
use FILL  FILL_7926
timestamp 1677622389
transform 1 0 3744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7928
timestamp 1677622389
transform 1 0 3752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7930
timestamp 1677622389
transform 1 0 3760 0 1 1570
box -8 -3 16 105
use FILL  FILL_7932
timestamp 1677622389
transform 1 0 3768 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_288
timestamp 1677622389
transform 1 0 3776 0 1 1570
box -8 -3 46 105
use FILL  FILL_7934
timestamp 1677622389
transform 1 0 3816 0 1 1570
box -8 -3 16 105
use FILL  FILL_7937
timestamp 1677622389
transform 1 0 3824 0 1 1570
box -8 -3 16 105
use FILL  FILL_7939
timestamp 1677622389
transform 1 0 3832 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_289
timestamp 1677622389
transform 1 0 3840 0 1 1570
box -8 -3 46 105
use FILL  FILL_7941
timestamp 1677622389
transform 1 0 3880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7948
timestamp 1677622389
transform 1 0 3888 0 1 1570
box -8 -3 16 105
use FILL  FILL_7949
timestamp 1677622389
transform 1 0 3896 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1677622389
transform -1 0 3928 0 1 1570
box -8 -3 32 105
use FILL  FILL_7950
timestamp 1677622389
transform 1 0 3928 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_290
timestamp 1677622389
transform 1 0 3936 0 1 1570
box -8 -3 46 105
use FILL  FILL_7953
timestamp 1677622389
transform 1 0 3976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7954
timestamp 1677622389
transform 1 0 3984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7955
timestamp 1677622389
transform 1 0 3992 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_291
timestamp 1677622389
transform 1 0 4000 0 1 1570
box -8 -3 46 105
use FILL  FILL_7960
timestamp 1677622389
transform 1 0 4040 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_292
timestamp 1677622389
transform -1 0 4088 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_293
timestamp 1677622389
transform -1 0 4128 0 1 1570
box -8 -3 46 105
use FILL  FILL_7961
timestamp 1677622389
transform 1 0 4128 0 1 1570
box -8 -3 16 105
use FILL  FILL_7970
timestamp 1677622389
transform 1 0 4136 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5822
timestamp 1677622389
transform 1 0 4180 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_294
timestamp 1677622389
transform 1 0 4144 0 1 1570
box -8 -3 46 105
use FILL  FILL_7971
timestamp 1677622389
transform 1 0 4184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7972
timestamp 1677622389
transform 1 0 4192 0 1 1570
box -8 -3 16 105
use FILL  FILL_7974
timestamp 1677622389
transform 1 0 4200 0 1 1570
box -8 -3 16 105
use FILL  FILL_7976
timestamp 1677622389
transform 1 0 4208 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_295
timestamp 1677622389
transform -1 0 4256 0 1 1570
box -8 -3 46 105
use FILL  FILL_7977
timestamp 1677622389
transform 1 0 4256 0 1 1570
box -8 -3 16 105
use FILL  FILL_7980
timestamp 1677622389
transform 1 0 4264 0 1 1570
box -8 -3 16 105
use FILL  FILL_7982
timestamp 1677622389
transform 1 0 4272 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_296
timestamp 1677622389
transform 1 0 4280 0 1 1570
box -8 -3 46 105
use FILL  FILL_7984
timestamp 1677622389
transform 1 0 4320 0 1 1570
box -8 -3 16 105
use FILL  FILL_7987
timestamp 1677622389
transform 1 0 4328 0 1 1570
box -8 -3 16 105
use FILL  FILL_7988
timestamp 1677622389
transform 1 0 4336 0 1 1570
box -8 -3 16 105
use FILL  FILL_7989
timestamp 1677622389
transform 1 0 4344 0 1 1570
box -8 -3 16 105
use FILL  FILL_7990
timestamp 1677622389
transform 1 0 4352 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_297
timestamp 1677622389
transform 1 0 4360 0 1 1570
box -8 -3 46 105
use FILL  FILL_7991
timestamp 1677622389
transform 1 0 4400 0 1 1570
box -8 -3 16 105
use FILL  FILL_7996
timestamp 1677622389
transform 1 0 4408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7998
timestamp 1677622389
transform 1 0 4416 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_298
timestamp 1677622389
transform 1 0 4424 0 1 1570
box -8 -3 46 105
use FILL  FILL_7999
timestamp 1677622389
transform 1 0 4464 0 1 1570
box -8 -3 16 105
use FILL  FILL_8003
timestamp 1677622389
transform 1 0 4472 0 1 1570
box -8 -3 16 105
use FILL  FILL_8004
timestamp 1677622389
transform 1 0 4480 0 1 1570
box -8 -3 16 105
use FILL  FILL_8005
timestamp 1677622389
transform 1 0 4488 0 1 1570
box -8 -3 16 105
use FILL  FILL_8006
timestamp 1677622389
transform 1 0 4496 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_299
timestamp 1677622389
transform -1 0 4544 0 1 1570
box -8 -3 46 105
use FILL  FILL_8007
timestamp 1677622389
transform 1 0 4544 0 1 1570
box -8 -3 16 105
use FILL  FILL_8008
timestamp 1677622389
transform 1 0 4552 0 1 1570
box -8 -3 16 105
use FILL  FILL_8009
timestamp 1677622389
transform 1 0 4560 0 1 1570
box -8 -3 16 105
use FILL  FILL_8010
timestamp 1677622389
transform 1 0 4568 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_300
timestamp 1677622389
transform 1 0 4576 0 1 1570
box -8 -3 46 105
use FILL  FILL_8011
timestamp 1677622389
transform 1 0 4616 0 1 1570
box -8 -3 16 105
use FILL  FILL_8023
timestamp 1677622389
transform 1 0 4624 0 1 1570
box -8 -3 16 105
use FILL  FILL_8025
timestamp 1677622389
transform 1 0 4632 0 1 1570
box -8 -3 16 105
use FILL  FILL_8027
timestamp 1677622389
transform 1 0 4640 0 1 1570
box -8 -3 16 105
use FILL  FILL_8028
timestamp 1677622389
transform 1 0 4648 0 1 1570
box -8 -3 16 105
use FILL  FILL_8029
timestamp 1677622389
transform 1 0 4656 0 1 1570
box -8 -3 16 105
use FILL  FILL_8030
timestamp 1677622389
transform 1 0 4664 0 1 1570
box -8 -3 16 105
use FILL  FILL_8031
timestamp 1677622389
transform 1 0 4672 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_429
timestamp 1677622389
transform 1 0 4680 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_504
timestamp 1677622389
transform -1 0 4792 0 1 1570
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_63
timestamp 1677622389
transform 1 0 4819 0 1 1570
box -10 -3 10 3
use M2_M1  M2_M1_6599
timestamp 1677622389
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1677622389
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5926
timestamp 1677622389
transform 1 0 132 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1677622389
transform 1 0 172 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6695
timestamp 1677622389
transform 1 0 196 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5928
timestamp 1677622389
transform 1 0 196 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1677622389
transform 1 0 188 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6600
timestamp 1677622389
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5879
timestamp 1677622389
transform 1 0 292 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6601
timestamp 1677622389
transform 1 0 316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1677622389
transform 1 0 324 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5899
timestamp 1677622389
transform 1 0 236 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1677622389
transform 1 0 332 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6603
timestamp 1677622389
transform 1 0 340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1677622389
transform 1 0 348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1677622389
transform 1 0 356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1677622389
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1677622389
transform 1 0 292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1677622389
transform 1 0 300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1677622389
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1677622389
transform 1 0 332 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5929
timestamp 1677622389
transform 1 0 236 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1677622389
transform 1 0 260 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1677622389
transform 1 0 300 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1677622389
transform 1 0 316 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1677622389
transform 1 0 332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1677622389
transform 1 0 252 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1677622389
transform 1 0 292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1677622389
transform 1 0 252 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1677622389
transform 1 0 356 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1677622389
transform 1 0 364 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6606
timestamp 1677622389
transform 1 0 404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5881
timestamp 1677622389
transform 1 0 412 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6607
timestamp 1677622389
transform 1 0 420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1677622389
transform 1 0 396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1677622389
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1677622389
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1677622389
transform 1 0 468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1677622389
transform 1 0 476 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5901
timestamp 1677622389
transform 1 0 468 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1677622389
transform 1 0 484 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6704
timestamp 1677622389
transform 1 0 492 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5835
timestamp 1677622389
transform 1 0 508 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6593
timestamp 1677622389
transform 1 0 508 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1677622389
transform 1 0 516 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5883
timestamp 1677622389
transform 1 0 532 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6611
timestamp 1677622389
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5902
timestamp 1677622389
transform 1 0 524 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6705
timestamp 1677622389
transform 1 0 532 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5935
timestamp 1677622389
transform 1 0 532 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6706
timestamp 1677622389
transform 1 0 556 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5823
timestamp 1677622389
transform 1 0 596 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6612
timestamp 1677622389
transform 1 0 596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1677622389
transform 1 0 620 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5988
timestamp 1677622389
transform 1 0 588 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1677622389
transform 1 0 596 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1677622389
transform 1 0 652 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6613
timestamp 1677622389
transform 1 0 684 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5936
timestamp 1677622389
transform 1 0 684 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1677622389
transform 1 0 700 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6614
timestamp 1677622389
transform 1 0 724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1677622389
transform 1 0 700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1677622389
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1677622389
transform 1 0 732 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5836
timestamp 1677622389
transform 1 0 748 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6711
timestamp 1677622389
transform 1 0 748 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1677622389
transform 1 0 756 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5999
timestamp 1677622389
transform 1 0 772 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1677622389
transform 1 0 804 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1677622389
transform 1 0 796 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1677622389
transform 1 0 820 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6616
timestamp 1677622389
transform 1 0 796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1677622389
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1677622389
transform 1 0 788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1677622389
transform 1 0 804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1677622389
transform 1 0 820 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5937
timestamp 1677622389
transform 1 0 788 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6715
timestamp 1677622389
transform 1 0 836 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5838
timestamp 1677622389
transform 1 0 860 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6618
timestamp 1677622389
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5854
timestamp 1677622389
transform 1 0 900 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6619
timestamp 1677622389
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5959
timestamp 1677622389
transform 1 0 908 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1677622389
transform 1 0 948 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6620
timestamp 1677622389
transform 1 0 948 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5884
timestamp 1677622389
transform 1 0 980 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5885
timestamp 1677622389
transform 1 0 996 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6716
timestamp 1677622389
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5903
timestamp 1677622389
transform 1 0 1020 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6717
timestamp 1677622389
transform 1 0 1028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1677622389
transform 1 0 1036 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5938
timestamp 1677622389
transform 1 0 996 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1677622389
transform 1 0 940 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1677622389
transform 1 0 1036 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6621
timestamp 1677622389
transform 1 0 1076 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5940
timestamp 1677622389
transform 1 0 1076 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6719
timestamp 1677622389
transform 1 0 1084 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5961
timestamp 1677622389
transform 1 0 1084 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6592
timestamp 1677622389
transform 1 0 1100 0 1 1555
box -2 -2 2 2
use M3_M2  M3_M2_5856
timestamp 1677622389
transform 1 0 1100 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1677622389
transform 1 0 1132 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6622
timestamp 1677622389
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5857
timestamp 1677622389
transform 1 0 1148 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6623
timestamp 1677622389
transform 1 0 1164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1677622389
transform 1 0 1140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1677622389
transform 1 0 1156 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5904
timestamp 1677622389
transform 1 0 1164 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1677622389
transform 1 0 1156 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1677622389
transform 1 0 1140 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6722
timestamp 1677622389
transform 1 0 1180 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5942
timestamp 1677622389
transform 1 0 1188 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6723
timestamp 1677622389
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5825
timestamp 1677622389
transform 1 0 1236 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6624
timestamp 1677622389
transform 1 0 1228 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5826
timestamp 1677622389
transform 1 0 1276 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1677622389
transform 1 0 1276 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6625
timestamp 1677622389
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1677622389
transform 1 0 1276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1677622389
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1677622389
transform 1 0 1284 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5943
timestamp 1677622389
transform 1 0 1276 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6726
timestamp 1677622389
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5905
timestamp 1677622389
transform 1 0 1324 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6627
timestamp 1677622389
transform 1 0 1420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1677622389
transform 1 0 1340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1677622389
transform 1 0 1396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1677622389
transform 1 0 1436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1677622389
transform 1 0 1444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5858
timestamp 1677622389
transform 1 0 1468 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1677622389
transform 1 0 1500 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5886
timestamp 1677622389
transform 1 0 1484 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6629
timestamp 1677622389
transform 1 0 1492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1677622389
transform 1 0 1468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6731
timestamp 1677622389
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6732
timestamp 1677622389
transform 1 0 1500 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5944
timestamp 1677622389
transform 1 0 1492 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1677622389
transform 1 0 1532 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6630
timestamp 1677622389
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5906
timestamp 1677622389
transform 1 0 1556 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1677622389
transform 1 0 1580 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6733
timestamp 1677622389
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5908
timestamp 1677622389
transform 1 0 1628 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6734
timestamp 1677622389
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1677622389
transform 1 0 1644 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5945
timestamp 1677622389
transform 1 0 1604 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1677622389
transform 1 0 1628 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1677622389
transform 1 0 1644 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6736
timestamp 1677622389
transform 1 0 1708 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5964
timestamp 1677622389
transform 1 0 1716 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6631
timestamp 1677622389
transform 1 0 1732 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5827
timestamp 1677622389
transform 1 0 1748 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1677622389
transform 1 0 1748 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1677622389
transform 1 0 1756 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6632
timestamp 1677622389
transform 1 0 1748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1677622389
transform 1 0 1764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6737
timestamp 1677622389
transform 1 0 1756 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5965
timestamp 1677622389
transform 1 0 1756 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1677622389
transform 1 0 1756 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1677622389
transform 1 0 1788 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1677622389
transform 1 0 1780 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6634
timestamp 1677622389
transform 1 0 1780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6738
timestamp 1677622389
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6739
timestamp 1677622389
transform 1 0 1836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6740
timestamp 1677622389
transform 1 0 1844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6741
timestamp 1677622389
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5843
timestamp 1677622389
transform 1 0 1900 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1677622389
transform 1 0 1876 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1677622389
transform 1 0 1892 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6635
timestamp 1677622389
transform 1 0 1876 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5966
timestamp 1677622389
transform 1 0 1868 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1677622389
transform 1 0 1892 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6636
timestamp 1677622389
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6742
timestamp 1677622389
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5909
timestamp 1677622389
transform 1 0 1900 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1677622389
transform 1 0 1924 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1677622389
transform 1 0 1916 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6743
timestamp 1677622389
transform 1 0 1908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1677622389
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6744
timestamp 1677622389
transform 1 0 1924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1677622389
transform 1 0 1916 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6821
timestamp 1677622389
transform 1 0 1932 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1677622389
transform 1 0 1948 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1677622389
transform 1 0 1972 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6745
timestamp 1677622389
transform 1 0 1948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1677622389
transform 1 0 1964 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5947
timestamp 1677622389
transform 1 0 1956 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1677622389
transform 1 0 1956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1677622389
transform 1 0 1972 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6640
timestamp 1677622389
transform 1 0 1996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6747
timestamp 1677622389
transform 1 0 1988 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5910
timestamp 1677622389
transform 1 0 1996 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1677622389
transform 1 0 1988 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1677622389
transform 1 0 2068 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6641
timestamp 1677622389
transform 1 0 2076 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6000
timestamp 1677622389
transform 1 0 2076 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6642
timestamp 1677622389
transform 1 0 2140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6748
timestamp 1677622389
transform 1 0 2172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1677622389
transform 1 0 2220 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5968
timestamp 1677622389
transform 1 0 2172 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6750
timestamp 1677622389
transform 1 0 2244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1677622389
transform 1 0 2236 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6822
timestamp 1677622389
transform 1 0 2228 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_5969
timestamp 1677622389
transform 1 0 2244 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6751
timestamp 1677622389
transform 1 0 2268 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5948
timestamp 1677622389
transform 1 0 2268 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6802
timestamp 1677622389
transform 1 0 2276 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5970
timestamp 1677622389
transform 1 0 2276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1677622389
transform 1 0 2300 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6752
timestamp 1677622389
transform 1 0 2316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1677622389
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6753
timestamp 1677622389
transform 1 0 2340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5829
timestamp 1677622389
transform 1 0 2380 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6754
timestamp 1677622389
transform 1 0 2380 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5992
timestamp 1677622389
transform 1 0 2388 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6644
timestamp 1677622389
transform 1 0 2404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5865
timestamp 1677622389
transform 1 0 2484 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1677622389
transform 1 0 2476 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6645
timestamp 1677622389
transform 1 0 2508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6755
timestamp 1677622389
transform 1 0 2428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6756
timestamp 1677622389
transform 1 0 2460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6757
timestamp 1677622389
transform 1 0 2484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5949
timestamp 1677622389
transform 1 0 2484 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1677622389
transform 1 0 2524 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1677622389
transform 1 0 2540 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6594
timestamp 1677622389
transform 1 0 2548 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_5868
timestamp 1677622389
transform 1 0 2596 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1677622389
transform 1 0 2548 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6646
timestamp 1677622389
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5911
timestamp 1677622389
transform 1 0 2604 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6758
timestamp 1677622389
transform 1 0 2636 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5950
timestamp 1677622389
transform 1 0 2636 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1677622389
transform 1 0 2684 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6647
timestamp 1677622389
transform 1 0 2780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6759
timestamp 1677622389
transform 1 0 2756 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5830
timestamp 1677622389
transform 1 0 2836 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1677622389
transform 1 0 2860 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6648
timestamp 1677622389
transform 1 0 2900 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5972
timestamp 1677622389
transform 1 0 2892 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6760
timestamp 1677622389
transform 1 0 2908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1677622389
transform 1 0 2924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6803
timestamp 1677622389
transform 1 0 2932 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5844
timestamp 1677622389
transform 1 0 3020 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6595
timestamp 1677622389
transform 1 0 3020 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1677622389
transform 1 0 3004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6762
timestamp 1677622389
transform 1 0 2996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6763
timestamp 1677622389
transform 1 0 3020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6764
timestamp 1677622389
transform 1 0 3028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1677622389
transform 1 0 3036 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5831
timestamp 1677622389
transform 1 0 3052 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1677622389
transform 1 0 3084 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6765
timestamp 1677622389
transform 1 0 3084 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5845
timestamp 1677622389
transform 1 0 3108 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6596
timestamp 1677622389
transform 1 0 3108 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1677622389
transform 1 0 3108 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5893
timestamp 1677622389
transform 1 0 3116 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6766
timestamp 1677622389
transform 1 0 3116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6767
timestamp 1677622389
transform 1 0 3124 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5951
timestamp 1677622389
transform 1 0 3116 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1677622389
transform 1 0 3148 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6652
timestamp 1677622389
transform 1 0 3148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6804
timestamp 1677622389
transform 1 0 3156 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5832
timestamp 1677622389
transform 1 0 3204 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1677622389
transform 1 0 3188 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6597
timestamp 1677622389
transform 1 0 3212 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1677622389
transform 1 0 3196 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1677622389
transform 1 0 3204 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5913
timestamp 1677622389
transform 1 0 3196 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1677622389
transform 1 0 3212 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6768
timestamp 1677622389
transform 1 0 3212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5952
timestamp 1677622389
transform 1 0 3204 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6655
timestamp 1677622389
transform 1 0 3244 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5914
timestamp 1677622389
transform 1 0 3244 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6805
timestamp 1677622389
transform 1 0 3268 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1677622389
transform 1 0 3284 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1677622389
transform 1 0 3308 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5869
timestamp 1677622389
transform 1 0 3332 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6656
timestamp 1677622389
transform 1 0 3332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6823
timestamp 1677622389
transform 1 0 3324 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_5973
timestamp 1677622389
transform 1 0 3332 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6657
timestamp 1677622389
transform 1 0 3364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1677622389
transform 1 0 3356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6771
timestamp 1677622389
transform 1 0 3372 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5847
timestamp 1677622389
transform 1 0 3396 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1677622389
transform 1 0 3396 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6658
timestamp 1677622389
transform 1 0 3404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5915
timestamp 1677622389
transform 1 0 3396 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1677622389
transform 1 0 3580 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1677622389
transform 1 0 3460 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6598
timestamp 1677622389
transform 1 0 3468 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_5872
timestamp 1677622389
transform 1 0 3556 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1677622389
transform 1 0 3572 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6659
timestamp 1677622389
transform 1 0 3460 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5974
timestamp 1677622389
transform 1 0 3452 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1677622389
transform 1 0 3468 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6772
timestamp 1677622389
transform 1 0 3556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1677622389
transform 1 0 3564 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5975
timestamp 1677622389
transform 1 0 3524 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1677622389
transform 1 0 3548 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6660
timestamp 1677622389
transform 1 0 3580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1677622389
transform 1 0 3596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1677622389
transform 1 0 3692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6774
timestamp 1677622389
transform 1 0 3628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6775
timestamp 1677622389
transform 1 0 3676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6776
timestamp 1677622389
transform 1 0 3684 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5896
timestamp 1677622389
transform 1 0 3724 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6777
timestamp 1677622389
transform 1 0 3716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6778
timestamp 1677622389
transform 1 0 3724 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5977
timestamp 1677622389
transform 1 0 3724 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6663
timestamp 1677622389
transform 1 0 3748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1677622389
transform 1 0 3756 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5953
timestamp 1677622389
transform 1 0 3748 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1677622389
transform 1 0 3788 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6779
timestamp 1677622389
transform 1 0 3796 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5918
timestamp 1677622389
transform 1 0 3812 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6807
timestamp 1677622389
transform 1 0 3812 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1677622389
transform 1 0 3836 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5897
timestamp 1677622389
transform 1 0 3876 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1677622389
transform 1 0 3900 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6666
timestamp 1677622389
transform 1 0 3892 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6780
timestamp 1677622389
transform 1 0 3884 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1677622389
transform 1 0 3916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1677622389
transform 1 0 3916 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5978
timestamp 1677622389
transform 1 0 3916 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1677622389
transform 1 0 3932 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6668
timestamp 1677622389
transform 1 0 3924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6781
timestamp 1677622389
transform 1 0 3956 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5954
timestamp 1677622389
transform 1 0 3948 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1677622389
transform 1 0 3988 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6809
timestamp 1677622389
transform 1 0 3988 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5993
timestamp 1677622389
transform 1 0 3972 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5994
timestamp 1677622389
transform 1 0 3988 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6782
timestamp 1677622389
transform 1 0 4020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1677622389
transform 1 0 4060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1677622389
transform 1 0 4076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6783
timestamp 1677622389
transform 1 0 4068 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5955
timestamp 1677622389
transform 1 0 4060 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6671
timestamp 1677622389
transform 1 0 4100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1677622389
transform 1 0 4124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6784
timestamp 1677622389
transform 1 0 4108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6785
timestamp 1677622389
transform 1 0 4116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1677622389
transform 1 0 4100 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5979
timestamp 1677622389
transform 1 0 4100 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5995
timestamp 1677622389
transform 1 0 4108 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1677622389
transform 1 0 4116 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6786
timestamp 1677622389
transform 1 0 4148 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5874
timestamp 1677622389
transform 1 0 4188 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6787
timestamp 1677622389
transform 1 0 4180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6788
timestamp 1677622389
transform 1 0 4188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6811
timestamp 1677622389
transform 1 0 4164 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5996
timestamp 1677622389
transform 1 0 4164 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6812
timestamp 1677622389
transform 1 0 4188 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5850
timestamp 1677622389
transform 1 0 4204 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6673
timestamp 1677622389
transform 1 0 4220 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5920
timestamp 1677622389
transform 1 0 4220 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1677622389
transform 1 0 4236 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1677622389
transform 1 0 4236 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6674
timestamp 1677622389
transform 1 0 4236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6789
timestamp 1677622389
transform 1 0 4236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6790
timestamp 1677622389
transform 1 0 4252 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5980
timestamp 1677622389
transform 1 0 4236 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1677622389
transform 1 0 4252 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6675
timestamp 1677622389
transform 1 0 4276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1677622389
transform 1 0 4292 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5898
timestamp 1677622389
transform 1 0 4308 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1677622389
transform 1 0 4324 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6677
timestamp 1677622389
transform 1 0 4316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6791
timestamp 1677622389
transform 1 0 4300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6813
timestamp 1677622389
transform 1 0 4316 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1677622389
transform 1 0 4324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6814
timestamp 1677622389
transform 1 0 4324 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5982
timestamp 1677622389
transform 1 0 4324 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1677622389
transform 1 0 4316 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6679
timestamp 1677622389
transform 1 0 4364 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5876
timestamp 1677622389
transform 1 0 4396 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6680
timestamp 1677622389
transform 1 0 4388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1677622389
transform 1 0 4396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1677622389
transform 1 0 4372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6793
timestamp 1677622389
transform 1 0 4380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6815
timestamp 1677622389
transform 1 0 4396 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5983
timestamp 1677622389
transform 1 0 4396 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6794
timestamp 1677622389
transform 1 0 4444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6816
timestamp 1677622389
transform 1 0 4428 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1677622389
transform 1 0 4460 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5921
timestamp 1677622389
transform 1 0 4460 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6817
timestamp 1677622389
transform 1 0 4460 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6004
timestamp 1677622389
transform 1 0 4460 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6795
timestamp 1677622389
transform 1 0 4476 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5922
timestamp 1677622389
transform 1 0 4484 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1677622389
transform 1 0 4500 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6818
timestamp 1677622389
transform 1 0 4484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1677622389
transform 1 0 4516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1677622389
transform 1 0 4524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1677622389
transform 1 0 4532 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5924
timestamp 1677622389
transform 1 0 4524 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6819
timestamp 1677622389
transform 1 0 4524 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5956
timestamp 1677622389
transform 1 0 4532 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1677622389
transform 1 0 4524 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6686
timestamp 1677622389
transform 1 0 4588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6796
timestamp 1677622389
transform 1 0 4572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6797
timestamp 1677622389
transform 1 0 4580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6798
timestamp 1677622389
transform 1 0 4628 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5985
timestamp 1677622389
transform 1 0 4628 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6687
timestamp 1677622389
transform 1 0 4660 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1677622389
transform 1 0 4676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1677622389
transform 1 0 4668 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5877
timestamp 1677622389
transform 1 0 4716 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6689
timestamp 1677622389
transform 1 0 4716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1677622389
transform 1 0 4732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1677622389
transform 1 0 4748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1677622389
transform 1 0 4740 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5878
timestamp 1677622389
transform 1 0 4772 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6692
timestamp 1677622389
transform 1 0 4764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1677622389
transform 1 0 4772 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5925
timestamp 1677622389
transform 1 0 4804 0 1 1525
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_64
timestamp 1677622389
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_410
timestamp 1677622389
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7555
timestamp 1677622389
transform 1 0 168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7556
timestamp 1677622389
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7557
timestamp 1677622389
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7558
timestamp 1677622389
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_411
timestamp 1677622389
transform 1 0 200 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_482
timestamp 1677622389
transform -1 0 312 0 -1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_282
timestamp 1677622389
transform 1 0 312 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7561
timestamp 1677622389
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7562
timestamp 1677622389
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7563
timestamp 1677622389
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7564
timestamp 1677622389
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_279
timestamp 1677622389
transform -1 0 424 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7565
timestamp 1677622389
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7566
timestamp 1677622389
transform 1 0 432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7567
timestamp 1677622389
transform 1 0 440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7568
timestamp 1677622389
transform 1 0 448 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_483
timestamp 1677622389
transform -1 0 472 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_484
timestamp 1677622389
transform 1 0 472 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7569
timestamp 1677622389
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7570
timestamp 1677622389
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7571
timestamp 1677622389
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_283
timestamp 1677622389
transform 1 0 512 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7572
timestamp 1677622389
transform 1 0 552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7574
timestamp 1677622389
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7576
timestamp 1677622389
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7578
timestamp 1677622389
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_414
timestamp 1677622389
transform 1 0 584 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7593
timestamp 1677622389
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7594
timestamp 1677622389
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7595
timestamp 1677622389
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_281
timestamp 1677622389
transform 1 0 704 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7596
timestamp 1677622389
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7598
timestamp 1677622389
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7600
timestamp 1677622389
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7602
timestamp 1677622389
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7604
timestamp 1677622389
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_285
timestamp 1677622389
transform 1 0 784 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7608
timestamp 1677622389
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7609
timestamp 1677622389
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7610
timestamp 1677622389
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7612
timestamp 1677622389
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7614
timestamp 1677622389
transform 1 0 856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7616
timestamp 1677622389
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_93
timestamp 1677622389
transform 1 0 872 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7621
timestamp 1677622389
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7623
timestamp 1677622389
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7625
timestamp 1677622389
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7627
timestamp 1677622389
transform 1 0 920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7636
timestamp 1677622389
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_415
timestamp 1677622389
transform 1 0 936 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7637
timestamp 1677622389
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7639
timestamp 1677622389
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7644
timestamp 1677622389
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_486
timestamp 1677622389
transform -1 0 1072 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7645
timestamp 1677622389
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7647
timestamp 1677622389
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7649
timestamp 1677622389
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7656
timestamp 1677622389
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7657
timestamp 1677622389
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7658
timestamp 1677622389
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7659
timestamp 1677622389
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7660
timestamp 1677622389
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_287
timestamp 1677622389
transform 1 0 1136 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7661
timestamp 1677622389
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7663
timestamp 1677622389
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7665
timestamp 1677622389
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7667
timestamp 1677622389
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7669
timestamp 1677622389
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7675
timestamp 1677622389
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7676
timestamp 1677622389
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7677
timestamp 1677622389
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7678
timestamp 1677622389
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_288
timestamp 1677622389
transform -1 0 1288 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7679
timestamp 1677622389
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7681
timestamp 1677622389
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7683
timestamp 1677622389
transform 1 0 1304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7685
timestamp 1677622389
transform 1 0 1312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7687
timestamp 1677622389
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7697
timestamp 1677622389
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_417
timestamp 1677622389
transform -1 0 1432 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7698
timestamp 1677622389
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7699
timestamp 1677622389
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7700
timestamp 1677622389
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7701
timestamp 1677622389
transform 1 0 1456 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_289
timestamp 1677622389
transform -1 0 1504 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7702
timestamp 1677622389
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7703
timestamp 1677622389
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7704
timestamp 1677622389
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7705
timestamp 1677622389
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7707
timestamp 1677622389
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_418
timestamp 1677622389
transform 1 0 1544 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7722
timestamp 1677622389
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_488
timestamp 1677622389
transform -1 0 1664 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7723
timestamp 1677622389
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7725
timestamp 1677622389
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7727
timestamp 1677622389
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7729
timestamp 1677622389
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7731
timestamp 1677622389
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7733
timestamp 1677622389
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7746
timestamp 1677622389
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7747
timestamp 1677622389
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7748
timestamp 1677622389
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_291
timestamp 1677622389
transform 1 0 1736 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7749
timestamp 1677622389
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7750
timestamp 1677622389
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7751
timestamp 1677622389
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7752
timestamp 1677622389
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7753
timestamp 1677622389
transform 1 0 1808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7754
timestamp 1677622389
transform 1 0 1816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7755
timestamp 1677622389
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_489
timestamp 1677622389
transform 1 0 1832 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7756
timestamp 1677622389
transform 1 0 1848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7757
timestamp 1677622389
transform 1 0 1856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7758
timestamp 1677622389
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_292
timestamp 1677622389
transform -1 0 1912 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7759
timestamp 1677622389
transform 1 0 1912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7760
timestamp 1677622389
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7761
timestamp 1677622389
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7762
timestamp 1677622389
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_293
timestamp 1677622389
transform -1 0 1984 0 -1 1570
box -8 -3 46 105
use M3_M2  M3_M2_6005
timestamp 1677622389
transform 1 0 1996 0 1 1475
box -3 -3 3 3
use FILL  FILL_7763
timestamp 1677622389
transform 1 0 1984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7764
timestamp 1677622389
transform 1 0 1992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7765
timestamp 1677622389
transform 1 0 2000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7768
timestamp 1677622389
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7769
timestamp 1677622389
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7770
timestamp 1677622389
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7771
timestamp 1677622389
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7772
timestamp 1677622389
transform 1 0 2040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7774
timestamp 1677622389
transform 1 0 2048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7776
timestamp 1677622389
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_490
timestamp 1677622389
transform -1 0 2080 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7777
timestamp 1677622389
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7785
timestamp 1677622389
transform 1 0 2088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7786
timestamp 1677622389
transform 1 0 2096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7787
timestamp 1677622389
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7788
timestamp 1677622389
transform 1 0 2112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7789
timestamp 1677622389
transform 1 0 2120 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_424
timestamp 1677622389
transform 1 0 2128 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7790
timestamp 1677622389
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_58
timestamp 1677622389
transform 1 0 2232 0 -1 1570
box -8 -3 40 105
use M3_M2  M3_M2_6006
timestamp 1677622389
transform 1 0 2276 0 1 1475
box -3 -3 3 3
use FILL  FILL_7791
timestamp 1677622389
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7792
timestamp 1677622389
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7793
timestamp 1677622389
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7794
timestamp 1677622389
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7795
timestamp 1677622389
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7796
timestamp 1677622389
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_97
timestamp 1677622389
transform 1 0 2312 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7797
timestamp 1677622389
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7798
timestamp 1677622389
transform 1 0 2344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7799
timestamp 1677622389
transform 1 0 2352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7800
timestamp 1677622389
transform 1 0 2360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7801
timestamp 1677622389
transform 1 0 2368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7802
timestamp 1677622389
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_98
timestamp 1677622389
transform 1 0 2384 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7803
timestamp 1677622389
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7804
timestamp 1677622389
transform 1 0 2416 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_425
timestamp 1677622389
transform -1 0 2520 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7805
timestamp 1677622389
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7824
timestamp 1677622389
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FAX1  FAX1_0
timestamp 1677622389
transform -1 0 2656 0 -1 1570
box -5 -3 126 105
use FILL  FILL_7825
timestamp 1677622389
transform 1 0 2656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7826
timestamp 1677622389
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7827
timestamp 1677622389
transform 1 0 2672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7828
timestamp 1677622389
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7829
timestamp 1677622389
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_427
timestamp 1677622389
transform -1 0 2792 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7830
timestamp 1677622389
transform 1 0 2792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7832
timestamp 1677622389
transform 1 0 2800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7834
timestamp 1677622389
transform 1 0 2808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7837
timestamp 1677622389
transform 1 0 2816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7838
timestamp 1677622389
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7839
timestamp 1677622389
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7840
timestamp 1677622389
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7841
timestamp 1677622389
transform 1 0 2848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7842
timestamp 1677622389
transform 1 0 2856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7843
timestamp 1677622389
transform 1 0 2864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7845
timestamp 1677622389
transform 1 0 2872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7847
timestamp 1677622389
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7849
timestamp 1677622389
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_130
timestamp 1677622389
transform 1 0 2896 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7851
timestamp 1677622389
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7853
timestamp 1677622389
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7855
timestamp 1677622389
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7857
timestamp 1677622389
transform 1 0 2952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7859
timestamp 1677622389
transform 1 0 2960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7861
timestamp 1677622389
transform 1 0 2968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7863
timestamp 1677622389
transform 1 0 2976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7865
timestamp 1677622389
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1677622389
transform 1 0 2992 0 -1 1570
box -7 -3 39 105
use INVX2  INVX2_494
timestamp 1677622389
transform -1 0 3040 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7869
timestamp 1677622389
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7871
timestamp 1677622389
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7873
timestamp 1677622389
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7875
timestamp 1677622389
transform 1 0 3064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7883
timestamp 1677622389
transform 1 0 3072 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1677622389
transform 1 0 3080 0 -1 1570
box -7 -3 39 105
use FILL  FILL_7884
timestamp 1677622389
transform 1 0 3112 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_131
timestamp 1677622389
transform 1 0 3120 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7885
timestamp 1677622389
transform 1 0 3152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7886
timestamp 1677622389
transform 1 0 3160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7887
timestamp 1677622389
transform 1 0 3168 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1677622389
transform -1 0 3208 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7888
timestamp 1677622389
transform 1 0 3208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7889
timestamp 1677622389
transform 1 0 3216 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1677622389
transform 1 0 3224 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7890
timestamp 1677622389
transform 1 0 3248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7891
timestamp 1677622389
transform 1 0 3256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7892
timestamp 1677622389
transform 1 0 3264 0 -1 1570
box -8 -3 16 105
use AND2X1  AND2X1_0
timestamp 1677622389
transform 1 0 3272 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7893
timestamp 1677622389
transform 1 0 3304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7895
timestamp 1677622389
transform 1 0 3312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7901
timestamp 1677622389
transform 1 0 3320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7902
timestamp 1677622389
transform 1 0 3328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7903
timestamp 1677622389
transform 1 0 3336 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_285
timestamp 1677622389
transform 1 0 3344 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7904
timestamp 1677622389
transform 1 0 3384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7905
timestamp 1677622389
transform 1 0 3392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7906
timestamp 1677622389
transform 1 0 3400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7909
timestamp 1677622389
transform 1 0 3408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7910
timestamp 1677622389
transform 1 0 3416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7911
timestamp 1677622389
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7912
timestamp 1677622389
transform 1 0 3432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7913
timestamp 1677622389
transform 1 0 3440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7914
timestamp 1677622389
transform 1 0 3448 0 -1 1570
box -8 -3 16 105
use FAX1  FAX1_3
timestamp 1677622389
transform -1 0 3576 0 -1 1570
box -5 -3 126 105
use FILL  FILL_7920
timestamp 1677622389
transform 1 0 3576 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_428
timestamp 1677622389
transform 1 0 3584 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7921
timestamp 1677622389
transform 1 0 3680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7923
timestamp 1677622389
transform 1 0 3688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7925
timestamp 1677622389
transform 1 0 3696 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_500
timestamp 1677622389
transform 1 0 3704 0 -1 1570
box -9 -3 26 105
use BUFX2  BUFX2_99
timestamp 1677622389
transform 1 0 3720 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7927
timestamp 1677622389
transform 1 0 3744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7929
timestamp 1677622389
transform 1 0 3752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7931
timestamp 1677622389
transform 1 0 3760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7933
timestamp 1677622389
transform 1 0 3768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7935
timestamp 1677622389
transform 1 0 3776 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_132
timestamp 1677622389
transform 1 0 3784 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7936
timestamp 1677622389
transform 1 0 3816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7938
timestamp 1677622389
transform 1 0 3824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7940
timestamp 1677622389
transform 1 0 3832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7942
timestamp 1677622389
transform 1 0 3840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7943
timestamp 1677622389
transform 1 0 3848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7944
timestamp 1677622389
transform 1 0 3856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7945
timestamp 1677622389
transform 1 0 3864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7946
timestamp 1677622389
transform 1 0 3872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7947
timestamp 1677622389
transform 1 0 3880 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_133
timestamp 1677622389
transform 1 0 3888 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7951
timestamp 1677622389
transform 1 0 3920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7952
timestamp 1677622389
transform 1 0 3928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7956
timestamp 1677622389
transform 1 0 3936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7957
timestamp 1677622389
transform 1 0 3944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7958
timestamp 1677622389
transform 1 0 3952 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_134
timestamp 1677622389
transform 1 0 3960 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7959
timestamp 1677622389
transform 1 0 3992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7962
timestamp 1677622389
transform 1 0 4000 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1677622389
transform -1 0 4032 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7963
timestamp 1677622389
transform 1 0 4032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7964
timestamp 1677622389
transform 1 0 4040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7965
timestamp 1677622389
transform 1 0 4048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7966
timestamp 1677622389
transform 1 0 4056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7967
timestamp 1677622389
transform 1 0 4064 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_135
timestamp 1677622389
transform 1 0 4072 0 -1 1570
box -8 -3 34 105
use INVX2  INVX2_501
timestamp 1677622389
transform -1 0 4120 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7968
timestamp 1677622389
transform 1 0 4120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7969
timestamp 1677622389
transform 1 0 4128 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_136
timestamp 1677622389
transform 1 0 4136 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_8
timestamp 1677622389
transform -1 0 4192 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7973
timestamp 1677622389
transform 1 0 4192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7975
timestamp 1677622389
transform 1 0 4200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7978
timestamp 1677622389
transform 1 0 4208 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_9
timestamp 1677622389
transform -1 0 4240 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_502
timestamp 1677622389
transform -1 0 4256 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7979
timestamp 1677622389
transform 1 0 4256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7981
timestamp 1677622389
transform 1 0 4264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7983
timestamp 1677622389
transform 1 0 4272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7985
timestamp 1677622389
transform 1 0 4280 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_137
timestamp 1677622389
transform 1 0 4288 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7986
timestamp 1677622389
transform 1 0 4320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7992
timestamp 1677622389
transform 1 0 4328 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_138
timestamp 1677622389
transform -1 0 4368 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7993
timestamp 1677622389
transform 1 0 4368 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_503
timestamp 1677622389
transform -1 0 4392 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7994
timestamp 1677622389
transform 1 0 4392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7995
timestamp 1677622389
transform 1 0 4400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7997
timestamp 1677622389
transform 1 0 4408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8000
timestamp 1677622389
transform 1 0 4416 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_139
timestamp 1677622389
transform -1 0 4456 0 -1 1570
box -8 -3 34 105
use FILL  FILL_8001
timestamp 1677622389
transform 1 0 4456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8002
timestamp 1677622389
transform 1 0 4464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8012
timestamp 1677622389
transform 1 0 4472 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_140
timestamp 1677622389
transform -1 0 4512 0 -1 1570
box -8 -3 34 105
use FILL  FILL_8013
timestamp 1677622389
transform 1 0 4512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8014
timestamp 1677622389
transform 1 0 4520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8015
timestamp 1677622389
transform 1 0 4528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8016
timestamp 1677622389
transform 1 0 4536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8017
timestamp 1677622389
transform 1 0 4544 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_141
timestamp 1677622389
transform -1 0 4584 0 -1 1570
box -8 -3 34 105
use FILL  FILL_8018
timestamp 1677622389
transform 1 0 4584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8019
timestamp 1677622389
transform 1 0 4592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8020
timestamp 1677622389
transform 1 0 4600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8021
timestamp 1677622389
transform 1 0 4608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8022
timestamp 1677622389
transform 1 0 4616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8024
timestamp 1677622389
transform 1 0 4624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8026
timestamp 1677622389
transform 1 0 4632 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_301
timestamp 1677622389
transform 1 0 4640 0 -1 1570
box -8 -3 46 105
use FILL  FILL_8032
timestamp 1677622389
transform 1 0 4680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8033
timestamp 1677622389
transform 1 0 4688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8034
timestamp 1677622389
transform 1 0 4696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8035
timestamp 1677622389
transform 1 0 4704 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_302
timestamp 1677622389
transform 1 0 4712 0 -1 1570
box -8 -3 46 105
use FILL  FILL_8036
timestamp 1677622389
transform 1 0 4752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8037
timestamp 1677622389
transform 1 0 4760 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_505
timestamp 1677622389
transform 1 0 4768 0 -1 1570
box -9 -3 26 105
use FILL  FILL_8038
timestamp 1677622389
transform 1 0 4784 0 -1 1570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_65
timestamp 1677622389
transform 1 0 4843 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_6025
timestamp 1677622389
transform 1 0 148 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6045
timestamp 1677622389
transform 1 0 68 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1677622389
transform 1 0 148 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6075
timestamp 1677622389
transform 1 0 68 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1677622389
transform 1 0 84 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1677622389
transform 1 0 188 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1677622389
transform 1 0 180 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6832
timestamp 1677622389
transform 1 0 108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6833
timestamp 1677622389
transform 1 0 164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1677622389
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6929
timestamp 1677622389
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6115
timestamp 1677622389
transform 1 0 84 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1677622389
transform 1 0 156 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1677622389
transform 1 0 228 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6048
timestamp 1677622389
transform 1 0 244 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6835
timestamp 1677622389
transform 1 0 188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6836
timestamp 1677622389
transform 1 0 204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6837
timestamp 1677622389
transform 1 0 220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6838
timestamp 1677622389
transform 1 0 228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6839
timestamp 1677622389
transform 1 0 244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6930
timestamp 1677622389
transform 1 0 180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6931
timestamp 1677622389
transform 1 0 188 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6117
timestamp 1677622389
transform 1 0 188 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6932
timestamp 1677622389
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6933
timestamp 1677622389
transform 1 0 236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6934
timestamp 1677622389
transform 1 0 252 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6140
timestamp 1677622389
transform 1 0 220 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6141
timestamp 1677622389
transform 1 0 252 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1677622389
transform 1 0 268 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6840
timestamp 1677622389
transform 1 0 268 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6014
timestamp 1677622389
transform 1 0 308 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6841
timestamp 1677622389
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6842
timestamp 1677622389
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6935
timestamp 1677622389
transform 1 0 292 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6101
timestamp 1677622389
transform 1 0 372 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6936
timestamp 1677622389
transform 1 0 380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6118
timestamp 1677622389
transform 1 0 380 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1677622389
transform 1 0 404 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6843
timestamp 1677622389
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6844
timestamp 1677622389
transform 1 0 420 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6077
timestamp 1677622389
transform 1 0 428 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6845
timestamp 1677622389
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6937
timestamp 1677622389
transform 1 0 412 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6102
timestamp 1677622389
transform 1 0 420 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6938
timestamp 1677622389
transform 1 0 428 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6119
timestamp 1677622389
transform 1 0 412 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1677622389
transform 1 0 452 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6846
timestamp 1677622389
transform 1 0 452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6939
timestamp 1677622389
transform 1 0 484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7005
timestamp 1677622389
transform 1 0 476 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1677622389
transform 1 0 524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6940
timestamp 1677622389
transform 1 0 516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6941
timestamp 1677622389
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6078
timestamp 1677622389
transform 1 0 548 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6942
timestamp 1677622389
transform 1 0 548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6848
timestamp 1677622389
transform 1 0 564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6943
timestamp 1677622389
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1677622389
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6016
timestamp 1677622389
transform 1 0 668 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1677622389
transform 1 0 700 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6850
timestamp 1677622389
transform 1 0 700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6944
timestamp 1677622389
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6050
timestamp 1677622389
transform 1 0 748 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6824
timestamp 1677622389
transform 1 0 756 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6851
timestamp 1677622389
transform 1 0 748 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6079
timestamp 1677622389
transform 1 0 756 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1677622389
transform 1 0 804 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6852
timestamp 1677622389
transform 1 0 796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6945
timestamp 1677622389
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6825
timestamp 1677622389
transform 1 0 820 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6080
timestamp 1677622389
transform 1 0 820 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6946
timestamp 1677622389
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6017
timestamp 1677622389
transform 1 0 860 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1677622389
transform 1 0 844 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6853
timestamp 1677622389
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6854
timestamp 1677622389
transform 1 0 860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6947
timestamp 1677622389
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6120
timestamp 1677622389
transform 1 0 860 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7006
timestamp 1677622389
transform 1 0 868 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6121
timestamp 1677622389
transform 1 0 900 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1677622389
transform 1 0 924 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6948
timestamp 1677622389
transform 1 0 916 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6029
timestamp 1677622389
transform 1 0 956 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_7007
timestamp 1677622389
transform 1 0 956 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6082
timestamp 1677622389
transform 1 0 996 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6855
timestamp 1677622389
transform 1 0 1004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6949
timestamp 1677622389
transform 1 0 996 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6083
timestamp 1677622389
transform 1 0 1028 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6856
timestamp 1677622389
transform 1 0 1036 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6103
timestamp 1677622389
transform 1 0 1036 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6142
timestamp 1677622389
transform 1 0 1028 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1677622389
transform 1 0 1068 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6857
timestamp 1677622389
transform 1 0 1092 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6085
timestamp 1677622389
transform 1 0 1140 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6950
timestamp 1677622389
transform 1 0 1068 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6122
timestamp 1677622389
transform 1 0 1068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6123
timestamp 1677622389
transform 1 0 1084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6124
timestamp 1677622389
transform 1 0 1140 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6143
timestamp 1677622389
transform 1 0 1068 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6144
timestamp 1677622389
transform 1 0 1140 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6858
timestamp 1677622389
transform 1 0 1156 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6053
timestamp 1677622389
transform 1 0 1220 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6086
timestamp 1677622389
transform 1 0 1172 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1677622389
transform 1 0 1260 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6859
timestamp 1677622389
transform 1 0 1220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6860
timestamp 1677622389
transform 1 0 1252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6861
timestamp 1677622389
transform 1 0 1260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6951
timestamp 1677622389
transform 1 0 1172 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6125
timestamp 1677622389
transform 1 0 1172 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6952
timestamp 1677622389
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6018
timestamp 1677622389
transform 1 0 1284 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1677622389
transform 1 0 1340 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1677622389
transform 1 0 1396 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1677622389
transform 1 0 1436 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6862
timestamp 1677622389
transform 1 0 1372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6863
timestamp 1677622389
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6953
timestamp 1677622389
transform 1 0 1348 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6126
timestamp 1677622389
transform 1 0 1348 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6954
timestamp 1677622389
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6019
timestamp 1677622389
transform 1 0 1492 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1677622389
transform 1 0 1484 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1677622389
transform 1 0 1508 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6864
timestamp 1677622389
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6865
timestamp 1677622389
transform 1 0 1484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6866
timestamp 1677622389
transform 1 0 1500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6867
timestamp 1677622389
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6955
timestamp 1677622389
transform 1 0 1492 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6145
timestamp 1677622389
transform 1 0 1500 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1677622389
transform 1 0 1660 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1677622389
transform 1 0 1564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6057
timestamp 1677622389
transform 1 0 1628 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1677622389
transform 1 0 1668 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6868
timestamp 1677622389
transform 1 0 1628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6869
timestamp 1677622389
transform 1 0 1660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6870
timestamp 1677622389
transform 1 0 1668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6956
timestamp 1677622389
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6957
timestamp 1677622389
transform 1 0 1580 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6104
timestamp 1677622389
transform 1 0 1700 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6146
timestamp 1677622389
transform 1 0 1708 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1677622389
transform 1 0 1764 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6033
timestamp 1677622389
transform 1 0 1740 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6871
timestamp 1677622389
transform 1 0 1732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6872
timestamp 1677622389
transform 1 0 1748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6873
timestamp 1677622389
transform 1 0 1764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6958
timestamp 1677622389
transform 1 0 1732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6959
timestamp 1677622389
transform 1 0 1740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6960
timestamp 1677622389
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6127
timestamp 1677622389
transform 1 0 1756 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6128
timestamp 1677622389
transform 1 0 1788 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6874
timestamp 1677622389
transform 1 0 1868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6961
timestamp 1677622389
transform 1 0 1820 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6129
timestamp 1677622389
transform 1 0 1820 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6130
timestamp 1677622389
transform 1 0 1868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1677622389
transform 1 0 2004 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1677622389
transform 1 0 1996 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6059
timestamp 1677622389
transform 1 0 1972 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6875
timestamp 1677622389
transform 1 0 1908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6876
timestamp 1677622389
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6131
timestamp 1677622389
transform 1 0 1908 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1677622389
transform 1 0 1964 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6877
timestamp 1677622389
transform 1 0 1972 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6105
timestamp 1677622389
transform 1 0 1948 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1677622389
transform 1 0 1972 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6962
timestamp 1677622389
transform 1 0 1996 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6132
timestamp 1677622389
transform 1 0 1996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1677622389
transform 1 0 2020 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1677622389
transform 1 0 2012 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6878
timestamp 1677622389
transform 1 0 2012 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6147
timestamp 1677622389
transform 1 0 2004 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1677622389
transform 1 0 2028 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6963
timestamp 1677622389
transform 1 0 2028 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6148
timestamp 1677622389
transform 1 0 2036 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6879
timestamp 1677622389
transform 1 0 2052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6880
timestamp 1677622389
transform 1 0 2108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6964
timestamp 1677622389
transform 1 0 2148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6133
timestamp 1677622389
transform 1 0 2124 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6134
timestamp 1677622389
transform 1 0 2148 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1677622389
transform 1 0 2220 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1677622389
transform 1 0 2252 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6881
timestamp 1677622389
transform 1 0 2212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6882
timestamp 1677622389
transform 1 0 2228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6965
timestamp 1677622389
transform 1 0 2188 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6135
timestamp 1677622389
transform 1 0 2188 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6883
timestamp 1677622389
transform 1 0 2324 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6010
timestamp 1677622389
transform 1 0 2404 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6884
timestamp 1677622389
transform 1 0 2412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6885
timestamp 1677622389
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6966
timestamp 1677622389
transform 1 0 2388 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6136
timestamp 1677622389
transform 1 0 2468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1677622389
transform 1 0 2604 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1677622389
transform 1 0 2644 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6036
timestamp 1677622389
transform 1 0 2540 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1677622389
transform 1 0 2596 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6886
timestamp 1677622389
transform 1 0 2580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6967
timestamp 1677622389
transform 1 0 2484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7008
timestamp 1677622389
transform 1 0 2492 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6038
timestamp 1677622389
transform 1 0 2636 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1677622389
transform 1 0 2668 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6040
timestamp 1677622389
transform 1 0 2764 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6061
timestamp 1677622389
transform 1 0 2628 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1677622389
transform 1 0 2660 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1677622389
transform 1 0 2724 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6887
timestamp 1677622389
transform 1 0 2628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6888
timestamp 1677622389
transform 1 0 2636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6889
timestamp 1677622389
transform 1 0 2660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6890
timestamp 1677622389
transform 1 0 2724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6891
timestamp 1677622389
transform 1 0 2764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6968
timestamp 1677622389
transform 1 0 2604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6969
timestamp 1677622389
transform 1 0 2612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6970
timestamp 1677622389
transform 1 0 2660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6971
timestamp 1677622389
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6972
timestamp 1677622389
transform 1 0 2764 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6137
timestamp 1677622389
transform 1 0 2660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6149
timestamp 1677622389
transform 1 0 2604 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6150
timestamp 1677622389
transform 1 0 2636 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1677622389
transform 1 0 2764 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6151
timestamp 1677622389
transform 1 0 2748 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1677622389
transform 1 0 2884 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1677622389
transform 1 0 2924 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6892
timestamp 1677622389
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6107
timestamp 1677622389
transform 1 0 2876 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1677622389
transform 1 0 2900 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6893
timestamp 1677622389
transform 1 0 2900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6894
timestamp 1677622389
transform 1 0 2908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6973
timestamp 1677622389
transform 1 0 2892 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6139
timestamp 1677622389
transform 1 0 2852 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7009
timestamp 1677622389
transform 1 0 2876 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6152
timestamp 1677622389
transform 1 0 2828 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_7010
timestamp 1677622389
transform 1 0 2996 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6895
timestamp 1677622389
transform 1 0 3012 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6089
timestamp 1677622389
transform 1 0 3020 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1677622389
transform 1 0 3012 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6974
timestamp 1677622389
transform 1 0 3052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6975
timestamp 1677622389
transform 1 0 3060 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6896
timestamp 1677622389
transform 1 0 3084 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6041
timestamp 1677622389
transform 1 0 3092 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6897
timestamp 1677622389
transform 1 0 3100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7011
timestamp 1677622389
transform 1 0 3092 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6153
timestamp 1677622389
transform 1 0 3092 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6042
timestamp 1677622389
transform 1 0 3116 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6976
timestamp 1677622389
transform 1 0 3108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6977
timestamp 1677622389
transform 1 0 3116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6898
timestamp 1677622389
transform 1 0 3124 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6090
timestamp 1677622389
transform 1 0 3132 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6978
timestamp 1677622389
transform 1 0 3132 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6154
timestamp 1677622389
transform 1 0 3148 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1677622389
transform 1 0 3196 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6826
timestamp 1677622389
transform 1 0 3252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6899
timestamp 1677622389
transform 1 0 3236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6900
timestamp 1677622389
transform 1 0 3244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6901
timestamp 1677622389
transform 1 0 3268 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6043
timestamp 1677622389
transform 1 0 3300 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6979
timestamp 1677622389
transform 1 0 3292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6980
timestamp 1677622389
transform 1 0 3300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6981
timestamp 1677622389
transform 1 0 3316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7012
timestamp 1677622389
transform 1 0 3332 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6982
timestamp 1677622389
transform 1 0 3348 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6044
timestamp 1677622389
transform 1 0 3364 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6902
timestamp 1677622389
transform 1 0 3396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6903
timestamp 1677622389
transform 1 0 3404 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6109
timestamp 1677622389
transform 1 0 3404 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6983
timestamp 1677622389
transform 1 0 3428 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6066
timestamp 1677622389
transform 1 0 3540 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6904
timestamp 1677622389
transform 1 0 3540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6905
timestamp 1677622389
transform 1 0 3548 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6067
timestamp 1677622389
transform 1 0 3564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1677622389
transform 1 0 3564 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1677622389
transform 1 0 3580 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6906
timestamp 1677622389
transform 1 0 3604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6907
timestamp 1677622389
transform 1 0 3660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6984
timestamp 1677622389
transform 1 0 3564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6985
timestamp 1677622389
transform 1 0 3580 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6093
timestamp 1677622389
transform 1 0 3692 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6908
timestamp 1677622389
transform 1 0 3724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6986
timestamp 1677622389
transform 1 0 3692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6909
timestamp 1677622389
transform 1 0 3780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6910
timestamp 1677622389
transform 1 0 3788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6987
timestamp 1677622389
transform 1 0 3788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6827
timestamp 1677622389
transform 1 0 3812 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6068
timestamp 1677622389
transform 1 0 3820 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6911
timestamp 1677622389
transform 1 0 3820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6988
timestamp 1677622389
transform 1 0 3820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6828
timestamp 1677622389
transform 1 0 3836 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6912
timestamp 1677622389
transform 1 0 3860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6989
timestamp 1677622389
transform 1 0 3876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6990
timestamp 1677622389
transform 1 0 3884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6991
timestamp 1677622389
transform 1 0 3908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6829
timestamp 1677622389
transform 1 0 3916 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6069
timestamp 1677622389
transform 1 0 3948 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6913
timestamp 1677622389
transform 1 0 3980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6992
timestamp 1677622389
transform 1 0 3948 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6110
timestamp 1677622389
transform 1 0 4020 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6914
timestamp 1677622389
transform 1 0 4036 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6915
timestamp 1677622389
transform 1 0 4044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6830
timestamp 1677622389
transform 1 0 4092 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6831
timestamp 1677622389
transform 1 0 4108 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6993
timestamp 1677622389
transform 1 0 4140 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6094
timestamp 1677622389
transform 1 0 4148 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6994
timestamp 1677622389
transform 1 0 4148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6095
timestamp 1677622389
transform 1 0 4188 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6995
timestamp 1677622389
transform 1 0 4180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6916
timestamp 1677622389
transform 1 0 4204 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6070
timestamp 1677622389
transform 1 0 4220 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1677622389
transform 1 0 4220 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6917
timestamp 1677622389
transform 1 0 4268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6996
timestamp 1677622389
transform 1 0 4220 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6111
timestamp 1677622389
transform 1 0 4268 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6918
timestamp 1677622389
transform 1 0 4324 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6112
timestamp 1677622389
transform 1 0 4332 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6997
timestamp 1677622389
transform 1 0 4356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6919
timestamp 1677622389
transform 1 0 4380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6998
timestamp 1677622389
transform 1 0 4388 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6113
timestamp 1677622389
transform 1 0 4396 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6999
timestamp 1677622389
transform 1 0 4420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6071
timestamp 1677622389
transform 1 0 4436 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6920
timestamp 1677622389
transform 1 0 4436 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6155
timestamp 1677622389
transform 1 0 4428 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1677622389
transform 1 0 4540 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1677622389
transform 1 0 4452 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6921
timestamp 1677622389
transform 1 0 4476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6922
timestamp 1677622389
transform 1 0 4532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6923
timestamp 1677622389
transform 1 0 4540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7000
timestamp 1677622389
transform 1 0 4452 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6114
timestamp 1677622389
transform 1 0 4476 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7001
timestamp 1677622389
transform 1 0 4548 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6073
timestamp 1677622389
transform 1 0 4604 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6074
timestamp 1677622389
transform 1 0 4660 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6098
timestamp 1677622389
transform 1 0 4572 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6924
timestamp 1677622389
transform 1 0 4620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6925
timestamp 1677622389
transform 1 0 4652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7002
timestamp 1677622389
transform 1 0 4572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6926
timestamp 1677622389
transform 1 0 4676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7003
timestamp 1677622389
transform 1 0 4668 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6156
timestamp 1677622389
transform 1 0 4564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6157
timestamp 1677622389
transform 1 0 4636 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6158
timestamp 1677622389
transform 1 0 4660 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1677622389
transform 1 0 4692 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1677622389
transform 1 0 4708 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6927
timestamp 1677622389
transform 1 0 4732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6928
timestamp 1677622389
transform 1 0 4788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7004
timestamp 1677622389
transform 1 0 4708 0 1 1405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_66
timestamp 1677622389
transform 1 0 48 0 1 1370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_430
timestamp 1677622389
transform 1 0 72 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_506
timestamp 1677622389
transform -1 0 184 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6159
timestamp 1677622389
transform 1 0 212 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_294
timestamp 1677622389
transform -1 0 224 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_295
timestamp 1677622389
transform -1 0 264 0 1 1370
box -8 -3 46 105
use FILL  FILL_8039
timestamp 1677622389
transform 1 0 264 0 1 1370
box -8 -3 16 105
use FILL  FILL_8040
timestamp 1677622389
transform 1 0 272 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6160
timestamp 1677622389
transform 1 0 300 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_431
timestamp 1677622389
transform 1 0 280 0 1 1370
box -8 -3 104 105
use FILL  FILL_8041
timestamp 1677622389
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_8042
timestamp 1677622389
transform 1 0 384 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_303
timestamp 1677622389
transform -1 0 432 0 1 1370
box -8 -3 46 105
use FILL  FILL_8043
timestamp 1677622389
transform 1 0 432 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_507
timestamp 1677622389
transform -1 0 456 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6161
timestamp 1677622389
transform 1 0 468 0 1 1375
box -3 -3 3 3
use FILL  FILL_8044
timestamp 1677622389
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_8045
timestamp 1677622389
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_8046
timestamp 1677622389
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_8047
timestamp 1677622389
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_8048
timestamp 1677622389
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8049
timestamp 1677622389
transform 1 0 496 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_296
timestamp 1677622389
transform 1 0 504 0 1 1370
box -8 -3 46 105
use FILL  FILL_8050
timestamp 1677622389
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_8051
timestamp 1677622389
transform 1 0 552 0 1 1370
box -8 -3 16 105
use FILL  FILL_8052
timestamp 1677622389
transform 1 0 560 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_100
timestamp 1677622389
transform -1 0 592 0 1 1370
box -5 -3 28 105
use FILL  FILL_8053
timestamp 1677622389
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_8054
timestamp 1677622389
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_8055
timestamp 1677622389
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_8056
timestamp 1677622389
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_8057
timestamp 1677622389
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_8058
timestamp 1677622389
transform 1 0 632 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_434
timestamp 1677622389
transform 1 0 640 0 1 1370
box -8 -3 104 105
use FILL  FILL_8082
timestamp 1677622389
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_8083
timestamp 1677622389
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_8084
timestamp 1677622389
transform 1 0 752 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_510
timestamp 1677622389
transform -1 0 776 0 1 1370
box -9 -3 26 105
use FILL  FILL_8085
timestamp 1677622389
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8086
timestamp 1677622389
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_8092
timestamp 1677622389
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_8094
timestamp 1677622389
transform 1 0 800 0 1 1370
box -8 -3 16 105
use FILL  FILL_8096
timestamp 1677622389
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_8097
timestamp 1677622389
transform 1 0 816 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_300
timestamp 1677622389
transform -1 0 864 0 1 1370
box -8 -3 46 105
use FILL  FILL_8098
timestamp 1677622389
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_8102
timestamp 1677622389
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_8104
timestamp 1677622389
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_8106
timestamp 1677622389
transform 1 0 888 0 1 1370
box -8 -3 16 105
use FILL  FILL_8107
timestamp 1677622389
transform 1 0 896 0 1 1370
box -8 -3 16 105
use FILL  FILL_8108
timestamp 1677622389
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_8109
timestamp 1677622389
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_8111
timestamp 1677622389
transform 1 0 920 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_82
timestamp 1677622389
transform 1 0 928 0 1 1370
box -8 -3 32 105
use FILL  FILL_8113
timestamp 1677622389
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_8118
timestamp 1677622389
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_8119
timestamp 1677622389
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8120
timestamp 1677622389
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8121
timestamp 1677622389
transform 1 0 984 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6162
timestamp 1677622389
transform 1 0 1004 0 1 1375
box -3 -3 3 3
use FILL  FILL_8123
timestamp 1677622389
transform 1 0 992 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_84
timestamp 1677622389
transform 1 0 1000 0 1 1370
box -8 -3 32 105
use FILL  FILL_8125
timestamp 1677622389
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8130
timestamp 1677622389
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use FILL  FILL_8132
timestamp 1677622389
transform 1 0 1040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8134
timestamp 1677622389
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_436
timestamp 1677622389
transform 1 0 1056 0 1 1370
box -8 -3 104 105
use FILL  FILL_8136
timestamp 1677622389
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_437
timestamp 1677622389
transform 1 0 1160 0 1 1370
box -8 -3 104 105
use FILL  FILL_8137
timestamp 1677622389
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_8138
timestamp 1677622389
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_8139
timestamp 1677622389
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_513
timestamp 1677622389
transform 1 0 1280 0 1 1370
box -9 -3 26 105
use FILL  FILL_8156
timestamp 1677622389
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_8160
timestamp 1677622389
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8161
timestamp 1677622389
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8162
timestamp 1677622389
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8163
timestamp 1677622389
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_438
timestamp 1677622389
transform 1 0 1336 0 1 1370
box -8 -3 104 105
use FILL  FILL_8164
timestamp 1677622389
transform 1 0 1432 0 1 1370
box -8 -3 16 105
use FILL  FILL_8165
timestamp 1677622389
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_8175
timestamp 1677622389
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use FILL  FILL_8177
timestamp 1677622389
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_304
timestamp 1677622389
transform -1 0 1504 0 1 1370
box -8 -3 46 105
use FILL  FILL_8178
timestamp 1677622389
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_8179
timestamp 1677622389
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_8183
timestamp 1677622389
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_8185
timestamp 1677622389
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_8186
timestamp 1677622389
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_8187
timestamp 1677622389
transform 1 0 1544 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_516
timestamp 1677622389
transform -1 0 1568 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6163
timestamp 1677622389
transform 1 0 1612 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_439
timestamp 1677622389
transform 1 0 1568 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_517
timestamp 1677622389
transform -1 0 1680 0 1 1370
box -9 -3 26 105
use FILL  FILL_8188
timestamp 1677622389
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8189
timestamp 1677622389
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_8190
timestamp 1677622389
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_8191
timestamp 1677622389
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_8192
timestamp 1677622389
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_8193
timestamp 1677622389
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6164
timestamp 1677622389
transform 1 0 1740 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6165
timestamp 1677622389
transform 1 0 1764 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_306
timestamp 1677622389
transform -1 0 1768 0 1 1370
box -8 -3 46 105
use FILL  FILL_8194
timestamp 1677622389
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8195
timestamp 1677622389
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8196
timestamp 1677622389
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_8210
timestamp 1677622389
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_8212
timestamp 1677622389
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_440
timestamp 1677622389
transform 1 0 1808 0 1 1370
box -8 -3 104 105
use FILL  FILL_8213
timestamp 1677622389
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_441
timestamp 1677622389
transform -1 0 2008 0 1 1370
box -8 -3 104 105
use FILL  FILL_8214
timestamp 1677622389
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_518
timestamp 1677622389
transform -1 0 2032 0 1 1370
box -9 -3 26 105
use FILL  FILL_8215
timestamp 1677622389
transform 1 0 2032 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6166
timestamp 1677622389
transform 1 0 2052 0 1 1375
box -3 -3 3 3
use FILL  FILL_8216
timestamp 1677622389
transform 1 0 2040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8217
timestamp 1677622389
transform 1 0 2048 0 1 1370
box -8 -3 16 105
use FILL  FILL_8218
timestamp 1677622389
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_442
timestamp 1677622389
transform -1 0 2160 0 1 1370
box -8 -3 104 105
use FILL  FILL_8219
timestamp 1677622389
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use FILL  FILL_8236
timestamp 1677622389
transform 1 0 2168 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_445
timestamp 1677622389
transform 1 0 2176 0 1 1370
box -8 -3 104 105
use FILL  FILL_8237
timestamp 1677622389
transform 1 0 2272 0 1 1370
box -8 -3 16 105
use FILL  FILL_8238
timestamp 1677622389
transform 1 0 2280 0 1 1370
box -8 -3 16 105
use FILL  FILL_8239
timestamp 1677622389
transform 1 0 2288 0 1 1370
box -8 -3 16 105
use FILL  FILL_8240
timestamp 1677622389
transform 1 0 2296 0 1 1370
box -8 -3 16 105
use FILL  FILL_8241
timestamp 1677622389
transform 1 0 2304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8242
timestamp 1677622389
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8243
timestamp 1677622389
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8244
timestamp 1677622389
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8245
timestamp 1677622389
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8246
timestamp 1677622389
transform 1 0 2344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8247
timestamp 1677622389
transform 1 0 2352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8248
timestamp 1677622389
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_8249
timestamp 1677622389
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_446
timestamp 1677622389
transform 1 0 2376 0 1 1370
box -8 -3 104 105
use FILL  FILL_8250
timestamp 1677622389
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_4
timestamp 1677622389
transform -1 0 2600 0 1 1370
box -5 -3 126 105
use FILL  FILL_8251
timestamp 1677622389
transform 1 0 2600 0 1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1677622389
transform -1 0 2664 0 1 1370
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_447
timestamp 1677622389
transform -1 0 2760 0 1 1370
box -8 -3 104 105
use FILL  FILL_8252
timestamp 1677622389
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1677622389
transform 1 0 2768 0 1 1370
box -5 -3 126 105
use FAX1  FAX1_6
timestamp 1677622389
transform 1 0 2888 0 1 1370
box -5 -3 126 105
use FILL  FILL_8253
timestamp 1677622389
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8284
timestamp 1677622389
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_8286
timestamp 1677622389
transform 1 0 3024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8288
timestamp 1677622389
transform 1 0 3032 0 1 1370
box -8 -3 16 105
use FILL  FILL_8289
timestamp 1677622389
transform 1 0 3040 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1677622389
transform 1 0 3048 0 1 1370
box -7 -3 39 105
use FILL  FILL_8290
timestamp 1677622389
transform 1 0 3080 0 1 1370
box -8 -3 16 105
use FILL  FILL_8291
timestamp 1677622389
transform 1 0 3088 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_521
timestamp 1677622389
transform -1 0 3112 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_522
timestamp 1677622389
transform 1 0 3112 0 1 1370
box -9 -3 26 105
use FILL  FILL_8292
timestamp 1677622389
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8293
timestamp 1677622389
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_8294
timestamp 1677622389
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_8299
timestamp 1677622389
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use FILL  FILL_8300
timestamp 1677622389
transform 1 0 3160 0 1 1370
box -8 -3 16 105
use FILL  FILL_8301
timestamp 1677622389
transform 1 0 3168 0 1 1370
box -8 -3 16 105
use FILL  FILL_8302
timestamp 1677622389
transform 1 0 3176 0 1 1370
box -8 -3 16 105
use FILL  FILL_8303
timestamp 1677622389
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_8304
timestamp 1677622389
transform 1 0 3192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8307
timestamp 1677622389
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use FILL  FILL_8309
timestamp 1677622389
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_8311
timestamp 1677622389
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_12
timestamp 1677622389
transform 1 0 3224 0 1 1370
box -8 -3 32 105
use FILL  FILL_8312
timestamp 1677622389
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_523
timestamp 1677622389
transform -1 0 3272 0 1 1370
box -9 -3 26 105
use FILL  FILL_8313
timestamp 1677622389
transform 1 0 3272 0 1 1370
box -8 -3 16 105
use FILL  FILL_8314
timestamp 1677622389
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use FILL  FILL_8315
timestamp 1677622389
transform 1 0 3288 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1677622389
transform -1 0 3328 0 1 1370
box -7 -3 39 105
use FILL  FILL_8316
timestamp 1677622389
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8325
timestamp 1677622389
transform 1 0 3336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8326
timestamp 1677622389
transform 1 0 3344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8327
timestamp 1677622389
transform 1 0 3352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8328
timestamp 1677622389
transform 1 0 3360 0 1 1370
box -8 -3 16 105
use FILL  FILL_8329
timestamp 1677622389
transform 1 0 3368 0 1 1370
box -8 -3 16 105
use FILL  FILL_8330
timestamp 1677622389
transform 1 0 3376 0 1 1370
box -8 -3 16 105
use FILL  FILL_8333
timestamp 1677622389
transform 1 0 3384 0 1 1370
box -8 -3 16 105
use FILL  FILL_8335
timestamp 1677622389
transform 1 0 3392 0 1 1370
box -8 -3 16 105
use FILL  FILL_8336
timestamp 1677622389
transform 1 0 3400 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_9
timestamp 1677622389
transform -1 0 3440 0 1 1370
box -7 -3 39 105
use FILL  FILL_8337
timestamp 1677622389
transform 1 0 3440 0 1 1370
box -8 -3 16 105
use FILL  FILL_8338
timestamp 1677622389
transform 1 0 3448 0 1 1370
box -8 -3 16 105
use FILL  FILL_8339
timestamp 1677622389
transform 1 0 3456 0 1 1370
box -8 -3 16 105
use FILL  FILL_8340
timestamp 1677622389
transform 1 0 3464 0 1 1370
box -8 -3 16 105
use FILL  FILL_8341
timestamp 1677622389
transform 1 0 3472 0 1 1370
box -8 -3 16 105
use FILL  FILL_8342
timestamp 1677622389
transform 1 0 3480 0 1 1370
box -8 -3 16 105
use FILL  FILL_8343
timestamp 1677622389
transform 1 0 3488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8344
timestamp 1677622389
transform 1 0 3496 0 1 1370
box -8 -3 16 105
use FILL  FILL_8345
timestamp 1677622389
transform 1 0 3504 0 1 1370
box -8 -3 16 105
use FILL  FILL_8346
timestamp 1677622389
transform 1 0 3512 0 1 1370
box -8 -3 16 105
use FILL  FILL_8348
timestamp 1677622389
transform 1 0 3520 0 1 1370
box -8 -3 16 105
use FILL  FILL_8349
timestamp 1677622389
transform 1 0 3528 0 1 1370
box -8 -3 16 105
use FILL  FILL_8350
timestamp 1677622389
transform 1 0 3536 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_102
timestamp 1677622389
transform 1 0 3544 0 1 1370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_451
timestamp 1677622389
transform 1 0 3568 0 1 1370
box -8 -3 104 105
use FILL  FILL_8351
timestamp 1677622389
transform 1 0 3664 0 1 1370
box -8 -3 16 105
use FILL  FILL_8352
timestamp 1677622389
transform 1 0 3672 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_452
timestamp 1677622389
transform 1 0 3680 0 1 1370
box -8 -3 104 105
use FILL  FILL_8363
timestamp 1677622389
transform 1 0 3776 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_144
timestamp 1677622389
transform 1 0 3784 0 1 1370
box -8 -3 34 105
use FILL  FILL_8364
timestamp 1677622389
transform 1 0 3816 0 1 1370
box -8 -3 16 105
use FILL  FILL_8365
timestamp 1677622389
transform 1 0 3824 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1677622389
transform -1 0 3856 0 1 1370
box -8 -3 32 105
use FILL  FILL_8366
timestamp 1677622389
transform 1 0 3856 0 1 1370
box -8 -3 16 105
use FILL  FILL_8380
timestamp 1677622389
transform 1 0 3864 0 1 1370
box -8 -3 16 105
use FILL  FILL_8382
timestamp 1677622389
transform 1 0 3872 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_145
timestamp 1677622389
transform 1 0 3880 0 1 1370
box -8 -3 34 105
use FILL  FILL_8384
timestamp 1677622389
transform 1 0 3912 0 1 1370
box -8 -3 16 105
use FILL  FILL_8390
timestamp 1677622389
transform 1 0 3920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8392
timestamp 1677622389
transform 1 0 3928 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_453
timestamp 1677622389
transform 1 0 3936 0 1 1370
box -8 -3 104 105
use FILL  FILL_8394
timestamp 1677622389
transform 1 0 4032 0 1 1370
box -8 -3 16 105
use FILL  FILL_8395
timestamp 1677622389
transform 1 0 4040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8396
timestamp 1677622389
transform 1 0 4048 0 1 1370
box -8 -3 16 105
use FILL  FILL_8397
timestamp 1677622389
transform 1 0 4056 0 1 1370
box -8 -3 16 105
use FILL  FILL_8398
timestamp 1677622389
transform 1 0 4064 0 1 1370
box -8 -3 16 105
use FILL  FILL_8399
timestamp 1677622389
transform 1 0 4072 0 1 1370
box -8 -3 16 105
use FILL  FILL_8400
timestamp 1677622389
transform 1 0 4080 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1677622389
transform -1 0 4112 0 1 1370
box -8 -3 32 105
use FILL  FILL_8401
timestamp 1677622389
transform 1 0 4112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8415
timestamp 1677622389
transform 1 0 4120 0 1 1370
box -8 -3 16 105
use FILL  FILL_8417
timestamp 1677622389
transform 1 0 4128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8419
timestamp 1677622389
transform 1 0 4136 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_146
timestamp 1677622389
transform -1 0 4176 0 1 1370
box -8 -3 34 105
use FILL  FILL_8420
timestamp 1677622389
transform 1 0 4176 0 1 1370
box -8 -3 16 105
use FILL  FILL_8421
timestamp 1677622389
transform 1 0 4184 0 1 1370
box -8 -3 16 105
use FILL  FILL_8422
timestamp 1677622389
transform 1 0 4192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8423
timestamp 1677622389
transform 1 0 4200 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_454
timestamp 1677622389
transform 1 0 4208 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6167
timestamp 1677622389
transform 1 0 4316 0 1 1375
box -3 -3 3 3
use FILL  FILL_8424
timestamp 1677622389
transform 1 0 4304 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_528
timestamp 1677622389
transform 1 0 4312 0 1 1370
box -9 -3 26 105
use FILL  FILL_8433
timestamp 1677622389
transform 1 0 4328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8434
timestamp 1677622389
transform 1 0 4336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8435
timestamp 1677622389
transform 1 0 4344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8436
timestamp 1677622389
transform 1 0 4352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8438
timestamp 1677622389
transform 1 0 4360 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_314
timestamp 1677622389
transform -1 0 4408 0 1 1370
box -8 -3 46 105
use M3_M2  M3_M2_6168
timestamp 1677622389
transform 1 0 4420 0 1 1375
box -3 -3 3 3
use FILL  FILL_8439
timestamp 1677622389
transform 1 0 4408 0 1 1370
box -8 -3 16 105
use FILL  FILL_8440
timestamp 1677622389
transform 1 0 4416 0 1 1370
box -8 -3 16 105
use FILL  FILL_8441
timestamp 1677622389
transform 1 0 4424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8442
timestamp 1677622389
transform 1 0 4432 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_456
timestamp 1677622389
transform 1 0 4440 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_529
timestamp 1677622389
transform -1 0 4552 0 1 1370
box -9 -3 26 105
use FILL  FILL_8443
timestamp 1677622389
transform 1 0 4552 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_457
timestamp 1677622389
transform 1 0 4560 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_530
timestamp 1677622389
transform -1 0 4672 0 1 1370
box -9 -3 26 105
use FILL  FILL_8444
timestamp 1677622389
transform 1 0 4672 0 1 1370
box -8 -3 16 105
use FILL  FILL_8458
timestamp 1677622389
transform 1 0 4680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8460
timestamp 1677622389
transform 1 0 4688 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_459
timestamp 1677622389
transform 1 0 4696 0 1 1370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_67
timestamp 1677622389
transform 1 0 4819 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_7127
timestamp 1677622389
transform 1 0 108 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6169
timestamp 1677622389
transform 1 0 180 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7019
timestamp 1677622389
transform 1 0 180 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6259
timestamp 1677622389
transform 1 0 180 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6170
timestamp 1677622389
transform 1 0 204 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6202
timestamp 1677622389
transform 1 0 236 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7020
timestamp 1677622389
transform 1 0 196 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6233
timestamp 1677622389
transform 1 0 228 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6203
timestamp 1677622389
transform 1 0 292 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7021
timestamp 1677622389
transform 1 0 284 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6234
timestamp 1677622389
transform 1 0 292 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7022
timestamp 1677622389
transform 1 0 300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7128
timestamp 1677622389
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7129
timestamp 1677622389
transform 1 0 284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7130
timestamp 1677622389
transform 1 0 308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7023
timestamp 1677622389
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6235
timestamp 1677622389
transform 1 0 332 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7131
timestamp 1677622389
transform 1 0 332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7132
timestamp 1677622389
transform 1 0 348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7024
timestamp 1677622389
transform 1 0 364 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6260
timestamp 1677622389
transform 1 0 364 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7025
timestamp 1677622389
transform 1 0 380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7026
timestamp 1677622389
transform 1 0 468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7027
timestamp 1677622389
transform 1 0 476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7028
timestamp 1677622389
transform 1 0 492 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6171
timestamp 1677622389
transform 1 0 508 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7133
timestamp 1677622389
transform 1 0 428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7134
timestamp 1677622389
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7135
timestamp 1677622389
transform 1 0 484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7136
timestamp 1677622389
transform 1 0 500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7137
timestamp 1677622389
transform 1 0 508 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6278
timestamp 1677622389
transform 1 0 460 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6279
timestamp 1677622389
transform 1 0 492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6323
timestamp 1677622389
transform 1 0 468 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6324
timestamp 1677622389
transform 1 0 500 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7029
timestamp 1677622389
transform 1 0 516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7030
timestamp 1677622389
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7031
timestamp 1677622389
transform 1 0 572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7138
timestamp 1677622389
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7139
timestamp 1677622389
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7140
timestamp 1677622389
transform 1 0 580 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6280
timestamp 1677622389
transform 1 0 572 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6325
timestamp 1677622389
transform 1 0 564 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7032
timestamp 1677622389
transform 1 0 612 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6236
timestamp 1677622389
transform 1 0 620 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7141
timestamp 1677622389
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6326
timestamp 1677622389
transform 1 0 604 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6204
timestamp 1677622389
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7033
timestamp 1677622389
transform 1 0 660 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6327
timestamp 1677622389
transform 1 0 660 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6186
timestamp 1677622389
transform 1 0 756 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6205
timestamp 1677622389
transform 1 0 676 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6206
timestamp 1677622389
transform 1 0 748 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7034
timestamp 1677622389
transform 1 0 676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7142
timestamp 1677622389
transform 1 0 724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7143
timestamp 1677622389
transform 1 0 756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7144
timestamp 1677622389
transform 1 0 764 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6281
timestamp 1677622389
transform 1 0 724 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6282
timestamp 1677622389
transform 1 0 764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6328
timestamp 1677622389
transform 1 0 764 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7035
timestamp 1677622389
transform 1 0 804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7145
timestamp 1677622389
transform 1 0 796 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6283
timestamp 1677622389
transform 1 0 804 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6172
timestamp 1677622389
transform 1 0 844 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6187
timestamp 1677622389
transform 1 0 820 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6207
timestamp 1677622389
transform 1 0 844 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7036
timestamp 1677622389
transform 1 0 820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7013
timestamp 1677622389
transform 1 0 860 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7037
timestamp 1677622389
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6237
timestamp 1677622389
transform 1 0 860 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7038
timestamp 1677622389
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7146
timestamp 1677622389
transform 1 0 836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7147
timestamp 1677622389
transform 1 0 852 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6284
timestamp 1677622389
transform 1 0 836 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6285
timestamp 1677622389
transform 1 0 852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6329
timestamp 1677622389
transform 1 0 884 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7014
timestamp 1677622389
transform 1 0 908 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6261
timestamp 1677622389
transform 1 0 908 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6286
timestamp 1677622389
transform 1 0 900 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6350
timestamp 1677622389
transform 1 0 916 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7039
timestamp 1677622389
transform 1 0 932 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6330
timestamp 1677622389
transform 1 0 932 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7148
timestamp 1677622389
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6287
timestamp 1677622389
transform 1 0 964 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7040
timestamp 1677622389
transform 1 0 980 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6288
timestamp 1677622389
transform 1 0 980 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6238
timestamp 1677622389
transform 1 0 1012 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6331
timestamp 1677622389
transform 1 0 1020 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7149
timestamp 1677622389
transform 1 0 1036 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6289
timestamp 1677622389
transform 1 0 1044 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6351
timestamp 1677622389
transform 1 0 1036 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7041
timestamp 1677622389
transform 1 0 1060 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6290
timestamp 1677622389
transform 1 0 1060 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6332
timestamp 1677622389
transform 1 0 1060 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7150
timestamp 1677622389
transform 1 0 1092 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6188
timestamp 1677622389
transform 1 0 1132 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6189
timestamp 1677622389
transform 1 0 1164 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6208
timestamp 1677622389
transform 1 0 1124 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6209
timestamp 1677622389
transform 1 0 1140 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6210
timestamp 1677622389
transform 1 0 1156 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7042
timestamp 1677622389
transform 1 0 1124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7043
timestamp 1677622389
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7044
timestamp 1677622389
transform 1 0 1156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7045
timestamp 1677622389
transform 1 0 1164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7151
timestamp 1677622389
transform 1 0 1140 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6291
timestamp 1677622389
transform 1 0 1140 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7152
timestamp 1677622389
transform 1 0 1164 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6333
timestamp 1677622389
transform 1 0 1164 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6173
timestamp 1677622389
transform 1 0 1188 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7046
timestamp 1677622389
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7153
timestamp 1677622389
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6334
timestamp 1677622389
transform 1 0 1212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6190
timestamp 1677622389
transform 1 0 1260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6211
timestamp 1677622389
transform 1 0 1268 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7047
timestamp 1677622389
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7048
timestamp 1677622389
transform 1 0 1268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7154
timestamp 1677622389
transform 1 0 1236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7155
timestamp 1677622389
transform 1 0 1252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7156
timestamp 1677622389
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6292
timestamp 1677622389
transform 1 0 1252 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6335
timestamp 1677622389
transform 1 0 1268 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6359
timestamp 1677622389
transform 1 0 1308 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6174
timestamp 1677622389
transform 1 0 1332 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6239
timestamp 1677622389
transform 1 0 1324 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7049
timestamp 1677622389
transform 1 0 1332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7050
timestamp 1677622389
transform 1 0 1348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7051
timestamp 1677622389
transform 1 0 1356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7157
timestamp 1677622389
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7158
timestamp 1677622389
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6293
timestamp 1677622389
transform 1 0 1356 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6336
timestamp 1677622389
transform 1 0 1348 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6360
timestamp 1677622389
transform 1 0 1324 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7159
timestamp 1677622389
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6191
timestamp 1677622389
transform 1 0 1428 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7160
timestamp 1677622389
transform 1 0 1428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7052
timestamp 1677622389
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7053
timestamp 1677622389
transform 1 0 1484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7054
timestamp 1677622389
transform 1 0 1500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7055
timestamp 1677622389
transform 1 0 1508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7161
timestamp 1677622389
transform 1 0 1468 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6294
timestamp 1677622389
transform 1 0 1468 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7162
timestamp 1677622389
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6337
timestamp 1677622389
transform 1 0 1484 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6192
timestamp 1677622389
transform 1 0 1524 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7056
timestamp 1677622389
transform 1 0 1524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7057
timestamp 1677622389
transform 1 0 1556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7163
timestamp 1677622389
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6262
timestamp 1677622389
transform 1 0 1556 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6295
timestamp 1677622389
transform 1 0 1556 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6361
timestamp 1677622389
transform 1 0 1548 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1677622389
transform 1 0 1580 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7058
timestamp 1677622389
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7059
timestamp 1677622389
transform 1 0 1596 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6240
timestamp 1677622389
transform 1 0 1604 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7060
timestamp 1677622389
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7164
timestamp 1677622389
transform 1 0 1604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7165
timestamp 1677622389
transform 1 0 1620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6296
timestamp 1677622389
transform 1 0 1604 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6362
timestamp 1677622389
transform 1 0 1620 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7166
timestamp 1677622389
transform 1 0 1636 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6297
timestamp 1677622389
transform 1 0 1636 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7061
timestamp 1677622389
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7062
timestamp 1677622389
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6263
timestamp 1677622389
transform 1 0 1652 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6193
timestamp 1677622389
transform 1 0 1708 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7063
timestamp 1677622389
transform 1 0 1700 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6264
timestamp 1677622389
transform 1 0 1684 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7167
timestamp 1677622389
transform 1 0 1692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7168
timestamp 1677622389
transform 1 0 1708 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6363
timestamp 1677622389
transform 1 0 1708 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6212
timestamp 1677622389
transform 1 0 1748 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6213
timestamp 1677622389
transform 1 0 1780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7064
timestamp 1677622389
transform 1 0 1748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7065
timestamp 1677622389
transform 1 0 1756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7066
timestamp 1677622389
transform 1 0 1780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7067
timestamp 1677622389
transform 1 0 1788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7169
timestamp 1677622389
transform 1 0 1740 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6352
timestamp 1677622389
transform 1 0 1740 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7170
timestamp 1677622389
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6298
timestamp 1677622389
transform 1 0 1764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6299
timestamp 1677622389
transform 1 0 1788 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6353
timestamp 1677622389
transform 1 0 1756 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6354
timestamp 1677622389
transform 1 0 1780 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6364
timestamp 1677622389
transform 1 0 1748 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7171
timestamp 1677622389
transform 1 0 1804 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6214
timestamp 1677622389
transform 1 0 1828 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7068
timestamp 1677622389
transform 1 0 1908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7172
timestamp 1677622389
transform 1 0 1820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7173
timestamp 1677622389
transform 1 0 1828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7174
timestamp 1677622389
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6300
timestamp 1677622389
transform 1 0 1820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6301
timestamp 1677622389
transform 1 0 1860 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6241
timestamp 1677622389
transform 1 0 1932 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7175
timestamp 1677622389
transform 1 0 1932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7230
timestamp 1677622389
transform 1 0 1964 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6176
timestamp 1677622389
transform 1 0 1980 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6177
timestamp 1677622389
transform 1 0 2020 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7069
timestamp 1677622389
transform 1 0 2076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7176
timestamp 1677622389
transform 1 0 2036 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6338
timestamp 1677622389
transform 1 0 2076 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6242
timestamp 1677622389
transform 1 0 2116 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6265
timestamp 1677622389
transform 1 0 2124 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7231
timestamp 1677622389
transform 1 0 2100 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6302
timestamp 1677622389
transform 1 0 2108 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6339
timestamp 1677622389
transform 1 0 2100 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7243
timestamp 1677622389
transform 1 0 2108 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_6178
timestamp 1677622389
transform 1 0 2140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6215
timestamp 1677622389
transform 1 0 2148 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7232
timestamp 1677622389
transform 1 0 2140 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7244
timestamp 1677622389
transform 1 0 2132 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_6266
timestamp 1677622389
transform 1 0 2156 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7233
timestamp 1677622389
transform 1 0 2164 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6179
timestamp 1677622389
transform 1 0 2236 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6194
timestamp 1677622389
transform 1 0 2260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6216
timestamp 1677622389
transform 1 0 2180 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7070
timestamp 1677622389
transform 1 0 2180 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6243
timestamp 1677622389
transform 1 0 2212 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7177
timestamp 1677622389
transform 1 0 2212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7178
timestamp 1677622389
transform 1 0 2260 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6303
timestamp 1677622389
transform 1 0 2180 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6304
timestamp 1677622389
transform 1 0 2204 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6305
timestamp 1677622389
transform 1 0 2220 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7179
timestamp 1677622389
transform 1 0 2276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6217
timestamp 1677622389
transform 1 0 2364 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6244
timestamp 1677622389
transform 1 0 2300 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6245
timestamp 1677622389
transform 1 0 2340 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7071
timestamp 1677622389
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7180
timestamp 1677622389
transform 1 0 2340 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6267
timestamp 1677622389
transform 1 0 2364 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7072
timestamp 1677622389
transform 1 0 2388 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6246
timestamp 1677622389
transform 1 0 2396 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7073
timestamp 1677622389
transform 1 0 2412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7181
timestamp 1677622389
transform 1 0 2396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7234
timestamp 1677622389
transform 1 0 2436 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7074
timestamp 1677622389
transform 1 0 2468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7182
timestamp 1677622389
transform 1 0 2476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7075
timestamp 1677622389
transform 1 0 2500 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6247
timestamp 1677622389
transform 1 0 2556 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7183
timestamp 1677622389
transform 1 0 2556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7076
timestamp 1677622389
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7077
timestamp 1677622389
transform 1 0 2636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7184
timestamp 1677622389
transform 1 0 2612 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7185
timestamp 1677622389
transform 1 0 2628 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6306
timestamp 1677622389
transform 1 0 2604 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7078
timestamp 1677622389
transform 1 0 2676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7186
timestamp 1677622389
transform 1 0 2668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7079
timestamp 1677622389
transform 1 0 2708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7187
timestamp 1677622389
transform 1 0 2700 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6307
timestamp 1677622389
transform 1 0 2700 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6268
timestamp 1677622389
transform 1 0 2740 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7080
timestamp 1677622389
transform 1 0 2828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7188
timestamp 1677622389
transform 1 0 2804 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6308
timestamp 1677622389
transform 1 0 2804 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6195
timestamp 1677622389
transform 1 0 2852 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7081
timestamp 1677622389
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7189
timestamp 1677622389
transform 1 0 2844 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6269
timestamp 1677622389
transform 1 0 2852 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7015
timestamp 1677622389
transform 1 0 2964 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6248
timestamp 1677622389
transform 1 0 2908 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6249
timestamp 1677622389
transform 1 0 2964 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7082
timestamp 1677622389
transform 1 0 2972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7083
timestamp 1677622389
transform 1 0 2980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7190
timestamp 1677622389
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6218
timestamp 1677622389
transform 1 0 3028 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7235
timestamp 1677622389
transform 1 0 3020 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7191
timestamp 1677622389
transform 1 0 3036 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6219
timestamp 1677622389
transform 1 0 3060 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7192
timestamp 1677622389
transform 1 0 3060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7236
timestamp 1677622389
transform 1 0 3036 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7237
timestamp 1677622389
transform 1 0 3044 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7238
timestamp 1677622389
transform 1 0 3068 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6340
timestamp 1677622389
transform 1 0 3068 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6220
timestamp 1677622389
transform 1 0 3084 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6221
timestamp 1677622389
transform 1 0 3100 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7016
timestamp 1677622389
transform 1 0 3116 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7084
timestamp 1677622389
transform 1 0 3084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7193
timestamp 1677622389
transform 1 0 3084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7245
timestamp 1677622389
transform 1 0 3076 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_7194
timestamp 1677622389
transform 1 0 3108 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7195
timestamp 1677622389
transform 1 0 3124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7085
timestamp 1677622389
transform 1 0 3140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7086
timestamp 1677622389
transform 1 0 3148 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6270
timestamp 1677622389
transform 1 0 3140 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7239
timestamp 1677622389
transform 1 0 3156 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6355
timestamp 1677622389
transform 1 0 3188 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6196
timestamp 1677622389
transform 1 0 3220 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7087
timestamp 1677622389
transform 1 0 3212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7088
timestamp 1677622389
transform 1 0 3220 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6309
timestamp 1677622389
transform 1 0 3212 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6356
timestamp 1677622389
transform 1 0 3212 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7089
timestamp 1677622389
transform 1 0 3300 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6250
timestamp 1677622389
transform 1 0 3308 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7090
timestamp 1677622389
transform 1 0 3316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7196
timestamp 1677622389
transform 1 0 3276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7197
timestamp 1677622389
transform 1 0 3292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7198
timestamp 1677622389
transform 1 0 3308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7199
timestamp 1677622389
transform 1 0 3316 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6341
timestamp 1677622389
transform 1 0 3292 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7017
timestamp 1677622389
transform 1 0 3324 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6310
timestamp 1677622389
transform 1 0 3316 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6197
timestamp 1677622389
transform 1 0 3372 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6222
timestamp 1677622389
transform 1 0 3364 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7091
timestamp 1677622389
transform 1 0 3364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7092
timestamp 1677622389
transform 1 0 3372 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6198
timestamp 1677622389
transform 1 0 3516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6223
timestamp 1677622389
transform 1 0 3428 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6224
timestamp 1677622389
transform 1 0 3444 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7018
timestamp 1677622389
transform 1 0 3500 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6251
timestamp 1677622389
transform 1 0 3500 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7093
timestamp 1677622389
transform 1 0 3516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7200
timestamp 1677622389
transform 1 0 3404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7201
timestamp 1677622389
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6271
timestamp 1677622389
transform 1 0 3508 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7202
timestamp 1677622389
transform 1 0 3516 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6225
timestamp 1677622389
transform 1 0 3532 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6199
timestamp 1677622389
transform 1 0 3556 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6272
timestamp 1677622389
transform 1 0 3548 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7094
timestamp 1677622389
transform 1 0 3588 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6252
timestamp 1677622389
transform 1 0 3596 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7095
timestamp 1677622389
transform 1 0 3604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7203
timestamp 1677622389
transform 1 0 3564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7204
timestamp 1677622389
transform 1 0 3572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7205
timestamp 1677622389
transform 1 0 3580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7206
timestamp 1677622389
transform 1 0 3596 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6311
timestamp 1677622389
transform 1 0 3580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6342
timestamp 1677622389
transform 1 0 3596 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6357
timestamp 1677622389
transform 1 0 3572 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7207
timestamp 1677622389
transform 1 0 3612 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6312
timestamp 1677622389
transform 1 0 3612 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6343
timestamp 1677622389
transform 1 0 3628 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7096
timestamp 1677622389
transform 1 0 3660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7097
timestamp 1677622389
transform 1 0 3676 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6253
timestamp 1677622389
transform 1 0 3716 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7098
timestamp 1677622389
transform 1 0 3724 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6254
timestamp 1677622389
transform 1 0 3732 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7099
timestamp 1677622389
transform 1 0 3740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7208
timestamp 1677622389
transform 1 0 3708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7209
timestamp 1677622389
transform 1 0 3716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7210
timestamp 1677622389
transform 1 0 3732 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6313
timestamp 1677622389
transform 1 0 3716 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6344
timestamp 1677622389
transform 1 0 3732 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6358
timestamp 1677622389
transform 1 0 3708 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7211
timestamp 1677622389
transform 1 0 3748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6314
timestamp 1677622389
transform 1 0 3748 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7100
timestamp 1677622389
transform 1 0 3780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7212
timestamp 1677622389
transform 1 0 3796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7240
timestamp 1677622389
transform 1 0 3820 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6345
timestamp 1677622389
transform 1 0 3836 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6200
timestamp 1677622389
transform 1 0 3956 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7101
timestamp 1677622389
transform 1 0 3956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7102
timestamp 1677622389
transform 1 0 3964 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6255
timestamp 1677622389
transform 1 0 3972 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7103
timestamp 1677622389
transform 1 0 3980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7213
timestamp 1677622389
transform 1 0 3972 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6226
timestamp 1677622389
transform 1 0 4028 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7104
timestamp 1677622389
transform 1 0 4028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7214
timestamp 1677622389
transform 1 0 4028 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6180
timestamp 1677622389
transform 1 0 4044 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6227
timestamp 1677622389
transform 1 0 4068 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7105
timestamp 1677622389
transform 1 0 4044 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6315
timestamp 1677622389
transform 1 0 4036 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6346
timestamp 1677622389
transform 1 0 4036 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6256
timestamp 1677622389
transform 1 0 4052 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7106
timestamp 1677622389
transform 1 0 4060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7107
timestamp 1677622389
transform 1 0 4076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7215
timestamp 1677622389
transform 1 0 4052 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6273
timestamp 1677622389
transform 1 0 4060 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7216
timestamp 1677622389
transform 1 0 4068 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6316
timestamp 1677622389
transform 1 0 4052 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6347
timestamp 1677622389
transform 1 0 4084 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6181
timestamp 1677622389
transform 1 0 4140 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7124
timestamp 1677622389
transform 1 0 4268 0 1 1333
box -2 -2 2 2
use M2_M1  M2_M1_7217
timestamp 1677622389
transform 1 0 4228 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6274
timestamp 1677622389
transform 1 0 4268 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6317
timestamp 1677622389
transform 1 0 4228 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7108
timestamp 1677622389
transform 1 0 4284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7109
timestamp 1677622389
transform 1 0 4316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7110
timestamp 1677622389
transform 1 0 4332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7218
timestamp 1677622389
transform 1 0 4324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7219
timestamp 1677622389
transform 1 0 4340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7111
timestamp 1677622389
transform 1 0 4356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7220
timestamp 1677622389
transform 1 0 4356 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6318
timestamp 1677622389
transform 1 0 4380 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7112
timestamp 1677622389
transform 1 0 4396 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6201
timestamp 1677622389
transform 1 0 4500 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7125
timestamp 1677622389
transform 1 0 4412 0 1 1333
box -2 -2 2 2
use M2_M1  M2_M1_7113
timestamp 1677622389
transform 1 0 4500 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6275
timestamp 1677622389
transform 1 0 4412 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7221
timestamp 1677622389
transform 1 0 4436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7222
timestamp 1677622389
transform 1 0 4492 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6319
timestamp 1677622389
transform 1 0 4436 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7241
timestamp 1677622389
transform 1 0 4508 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6182
timestamp 1677622389
transform 1 0 4540 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7126
timestamp 1677622389
transform 1 0 4532 0 1 1333
box -2 -2 2 2
use M2_M1  M2_M1_7114
timestamp 1677622389
transform 1 0 4540 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6348
timestamp 1677622389
transform 1 0 4508 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6349
timestamp 1677622389
transform 1 0 4524 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6320
timestamp 1677622389
transform 1 0 4540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6228
timestamp 1677622389
transform 1 0 4556 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7223
timestamp 1677622389
transform 1 0 4556 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6257
timestamp 1677622389
transform 1 0 4580 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6229
timestamp 1677622389
transform 1 0 4596 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7115
timestamp 1677622389
transform 1 0 4588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7242
timestamp 1677622389
transform 1 0 4564 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6183
timestamp 1677622389
transform 1 0 4620 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7116
timestamp 1677622389
transform 1 0 4612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7117
timestamp 1677622389
transform 1 0 4620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7224
timestamp 1677622389
transform 1 0 4612 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6321
timestamp 1677622389
transform 1 0 4612 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6258
timestamp 1677622389
transform 1 0 4628 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7118
timestamp 1677622389
transform 1 0 4636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7225
timestamp 1677622389
transform 1 0 4644 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7226
timestamp 1677622389
transform 1 0 4668 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6322
timestamp 1677622389
transform 1 0 4676 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6184
timestamp 1677622389
transform 1 0 4700 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6230
timestamp 1677622389
transform 1 0 4692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6231
timestamp 1677622389
transform 1 0 4732 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7119
timestamp 1677622389
transform 1 0 4692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7120
timestamp 1677622389
transform 1 0 4700 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7121
timestamp 1677622389
transform 1 0 4716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7122
timestamp 1677622389
transform 1 0 4732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7227
timestamp 1677622389
transform 1 0 4708 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6276
timestamp 1677622389
transform 1 0 4716 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7228
timestamp 1677622389
transform 1 0 4724 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6277
timestamp 1677622389
transform 1 0 4732 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7229
timestamp 1677622389
transform 1 0 4740 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6232
timestamp 1677622389
transform 1 0 4748 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6185
timestamp 1677622389
transform 1 0 4772 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7123
timestamp 1677622389
transform 1 0 4788 0 1 1335
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_68
timestamp 1677622389
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_8059
timestamp 1677622389
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8060
timestamp 1677622389
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8061
timestamp 1677622389
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8062
timestamp 1677622389
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8063
timestamp 1677622389
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8064
timestamp 1677622389
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8065
timestamp 1677622389
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8066
timestamp 1677622389
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_508
timestamp 1677622389
transform -1 0 152 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8067
timestamp 1677622389
transform 1 0 152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8068
timestamp 1677622389
transform 1 0 160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8069
timestamp 1677622389
transform 1 0 168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8070
timestamp 1677622389
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_432
timestamp 1677622389
transform 1 0 184 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_509
timestamp 1677622389
transform 1 0 280 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8071
timestamp 1677622389
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8072
timestamp 1677622389
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_297
timestamp 1677622389
transform 1 0 312 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8073
timestamp 1677622389
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8074
timestamp 1677622389
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6365
timestamp 1677622389
transform 1 0 412 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_433
timestamp 1677622389
transform 1 0 368 0 -1 1370
box -8 -3 104 105
use AOI22X1  AOI22X1_298
timestamp 1677622389
transform 1 0 464 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8075
timestamp 1677622389
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8076
timestamp 1677622389
transform 1 0 512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8077
timestamp 1677622389
transform 1 0 520 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_299
timestamp 1677622389
transform 1 0 528 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8078
timestamp 1677622389
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8079
timestamp 1677622389
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8080
timestamp 1677622389
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6366
timestamp 1677622389
transform 1 0 620 0 1 1275
box -3 -3 3 3
use OAI22X1  OAI22X1_304
timestamp 1677622389
transform 1 0 592 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8081
timestamp 1677622389
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8087
timestamp 1677622389
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8088
timestamp 1677622389
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6367
timestamp 1677622389
transform 1 0 668 0 1 1275
box -3 -3 3 3
use FILL  FILL_8089
timestamp 1677622389
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_435
timestamp 1677622389
transform 1 0 664 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8090
timestamp 1677622389
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_511
timestamp 1677622389
transform -1 0 784 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8091
timestamp 1677622389
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8093
timestamp 1677622389
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8095
timestamp 1677622389
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8099
timestamp 1677622389
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_301
timestamp 1677622389
transform -1 0 856 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8100
timestamp 1677622389
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8101
timestamp 1677622389
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8103
timestamp 1677622389
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8105
timestamp 1677622389
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_81
timestamp 1677622389
transform 1 0 888 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8110
timestamp 1677622389
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8112
timestamp 1677622389
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8114
timestamp 1677622389
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8115
timestamp 1677622389
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8116
timestamp 1677622389
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8117
timestamp 1677622389
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_83
timestamp 1677622389
transform 1 0 960 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8122
timestamp 1677622389
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8124
timestamp 1677622389
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8126
timestamp 1677622389
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8127
timestamp 1677622389
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8128
timestamp 1677622389
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8129
timestamp 1677622389
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8131
timestamp 1677622389
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8133
timestamp 1677622389
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8135
timestamp 1677622389
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6368
timestamp 1677622389
transform 1 0 1084 0 1 1275
box -3 -3 3 3
use INVX2  INVX2_512
timestamp 1677622389
transform 1 0 1056 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8140
timestamp 1677622389
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8141
timestamp 1677622389
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8142
timestamp 1677622389
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8143
timestamp 1677622389
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8144
timestamp 1677622389
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8145
timestamp 1677622389
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_302
timestamp 1677622389
transform 1 0 1120 0 -1 1370
box -8 -3 46 105
use M3_M2  M3_M2_6369
timestamp 1677622389
transform 1 0 1172 0 1 1275
box -3 -3 3 3
use FILL  FILL_8146
timestamp 1677622389
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8147
timestamp 1677622389
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8148
timestamp 1677622389
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8149
timestamp 1677622389
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8150
timestamp 1677622389
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8151
timestamp 1677622389
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8152
timestamp 1677622389
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8153
timestamp 1677622389
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8154
timestamp 1677622389
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_303
timestamp 1677622389
transform 1 0 1232 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8155
timestamp 1677622389
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8157
timestamp 1677622389
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8158
timestamp 1677622389
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8159
timestamp 1677622389
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8166
timestamp 1677622389
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_305
timestamp 1677622389
transform -1 0 1352 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8167
timestamp 1677622389
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_514
timestamp 1677622389
transform 1 0 1360 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8168
timestamp 1677622389
transform 1 0 1376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8169
timestamp 1677622389
transform 1 0 1384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8170
timestamp 1677622389
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8171
timestamp 1677622389
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8172
timestamp 1677622389
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8173
timestamp 1677622389
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_515
timestamp 1677622389
transform -1 0 1440 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8174
timestamp 1677622389
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8176
timestamp 1677622389
transform 1 0 1448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8180
timestamp 1677622389
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8181
timestamp 1677622389
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_305
timestamp 1677622389
transform -1 0 1512 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8182
timestamp 1677622389
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8184
timestamp 1677622389
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8197
timestamp 1677622389
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_306
timestamp 1677622389
transform -1 0 1576 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8198
timestamp 1677622389
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8199
timestamp 1677622389
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_307
timestamp 1677622389
transform 1 0 1592 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8200
timestamp 1677622389
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8201
timestamp 1677622389
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8202
timestamp 1677622389
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8203
timestamp 1677622389
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8204
timestamp 1677622389
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8205
timestamp 1677622389
transform 1 0 1672 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_308
timestamp 1677622389
transform 1 0 1680 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8206
timestamp 1677622389
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8207
timestamp 1677622389
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8208
timestamp 1677622389
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_307
timestamp 1677622389
transform 1 0 1744 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8209
timestamp 1677622389
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8211
timestamp 1677622389
transform 1 0 1792 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_519
timestamp 1677622389
transform 1 0 1800 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8220
timestamp 1677622389
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_443
timestamp 1677622389
transform -1 0 1920 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8221
timestamp 1677622389
transform 1 0 1920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8222
timestamp 1677622389
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8223
timestamp 1677622389
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8224
timestamp 1677622389
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8225
timestamp 1677622389
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8226
timestamp 1677622389
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8227
timestamp 1677622389
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8228
timestamp 1677622389
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8229
timestamp 1677622389
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_444
timestamp 1677622389
transform -1 0 2088 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8230
timestamp 1677622389
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_62
timestamp 1677622389
transform -1 0 2128 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8231
timestamp 1677622389
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8232
timestamp 1677622389
transform 1 0 2136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8233
timestamp 1677622389
transform 1 0 2144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8234
timestamp 1677622389
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8235
timestamp 1677622389
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_448
timestamp 1677622389
transform 1 0 2168 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8254
timestamp 1677622389
transform 1 0 2264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8255
timestamp 1677622389
transform 1 0 2272 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6370
timestamp 1677622389
transform 1 0 2292 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_449
timestamp 1677622389
transform -1 0 2376 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8256
timestamp 1677622389
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_142
timestamp 1677622389
transform 1 0 2384 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8257
timestamp 1677622389
transform 1 0 2416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8258
timestamp 1677622389
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_10
timestamp 1677622389
transform -1 0 2456 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8259
timestamp 1677622389
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8260
timestamp 1677622389
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8261
timestamp 1677622389
transform 1 0 2472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8262
timestamp 1677622389
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8263
timestamp 1677622389
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8264
timestamp 1677622389
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8265
timestamp 1677622389
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8266
timestamp 1677622389
transform 1 0 2512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8267
timestamp 1677622389
transform 1 0 2520 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1677622389
transform 1 0 2528 0 -1 1370
box -7 -3 39 105
use FILL  FILL_8268
timestamp 1677622389
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8269
timestamp 1677622389
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8270
timestamp 1677622389
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_520
timestamp 1677622389
transform -1 0 2600 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8271
timestamp 1677622389
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_51
timestamp 1677622389
transform -1 0 2640 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8272
timestamp 1677622389
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8273
timestamp 1677622389
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8274
timestamp 1677622389
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8275
timestamp 1677622389
transform 1 0 2664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8276
timestamp 1677622389
transform 1 0 2672 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_308
timestamp 1677622389
transform 1 0 2680 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8277
timestamp 1677622389
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8278
timestamp 1677622389
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8279
timestamp 1677622389
transform 1 0 2736 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_450
timestamp 1677622389
transform -1 0 2840 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8280
timestamp 1677622389
transform 1 0 2840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8281
timestamp 1677622389
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_7
timestamp 1677622389
transform 1 0 2856 0 -1 1370
box -5 -3 126 105
use NAND2X1  NAND2X1_11
timestamp 1677622389
transform 1 0 2976 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8282
timestamp 1677622389
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8283
timestamp 1677622389
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8285
timestamp 1677622389
transform 1 0 3016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8287
timestamp 1677622389
transform 1 0 3024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8295
timestamp 1677622389
transform 1 0 3032 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_63
timestamp 1677622389
transform -1 0 3072 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8296
timestamp 1677622389
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_6
timestamp 1677622389
transform 1 0 3080 0 -1 1370
box -7 -3 39 105
use FILL  FILL_8297
timestamp 1677622389
transform 1 0 3112 0 -1 1370
box -8 -3 16 105
use BUFX2  BUFX2_101
timestamp 1677622389
transform 1 0 3120 0 -1 1370
box -5 -3 28 105
use FILL  FILL_8298
timestamp 1677622389
transform 1 0 3144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8305
timestamp 1677622389
transform 1 0 3152 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_143
timestamp 1677622389
transform -1 0 3192 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8306
timestamp 1677622389
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8308
timestamp 1677622389
transform 1 0 3200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8310
timestamp 1677622389
transform 1 0 3208 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_524
timestamp 1677622389
transform 1 0 3216 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8317
timestamp 1677622389
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8318
timestamp 1677622389
transform 1 0 3240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8319
timestamp 1677622389
transform 1 0 3248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8320
timestamp 1677622389
transform 1 0 3256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8321
timestamp 1677622389
transform 1 0 3264 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_309
timestamp 1677622389
transform 1 0 3272 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8322
timestamp 1677622389
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8323
timestamp 1677622389
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8324
timestamp 1677622389
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8331
timestamp 1677622389
transform 1 0 3336 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_8
timestamp 1677622389
transform -1 0 3376 0 -1 1370
box -7 -3 39 105
use M3_M2  M3_M2_6371
timestamp 1677622389
transform 1 0 3388 0 1 1275
box -3 -3 3 3
use FILL  FILL_8332
timestamp 1677622389
transform 1 0 3376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8334
timestamp 1677622389
transform 1 0 3384 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_8
timestamp 1677622389
transform 1 0 3392 0 -1 1370
box -5 -3 126 105
use FILL  FILL_8347
timestamp 1677622389
transform 1 0 3512 0 -1 1370
box -8 -3 16 105
use BUFX2  BUFX2_103
timestamp 1677622389
transform 1 0 3520 0 -1 1370
box -5 -3 28 105
use FILL  FILL_8353
timestamp 1677622389
transform 1 0 3544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8354
timestamp 1677622389
transform 1 0 3552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8355
timestamp 1677622389
transform 1 0 3560 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_309
timestamp 1677622389
transform 1 0 3568 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8356
timestamp 1677622389
transform 1 0 3608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8357
timestamp 1677622389
transform 1 0 3616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8358
timestamp 1677622389
transform 1 0 3624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8359
timestamp 1677622389
transform 1 0 3632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8360
timestamp 1677622389
transform 1 0 3640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8361
timestamp 1677622389
transform 1 0 3648 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_525
timestamp 1677622389
transform 1 0 3656 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8362
timestamp 1677622389
transform 1 0 3672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8367
timestamp 1677622389
transform 1 0 3680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8368
timestamp 1677622389
transform 1 0 3688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8369
timestamp 1677622389
transform 1 0 3696 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_310
timestamp 1677622389
transform 1 0 3704 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8370
timestamp 1677622389
transform 1 0 3744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8371
timestamp 1677622389
transform 1 0 3752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8372
timestamp 1677622389
transform 1 0 3760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8373
timestamp 1677622389
transform 1 0 3768 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_526
timestamp 1677622389
transform 1 0 3776 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8374
timestamp 1677622389
transform 1 0 3792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8375
timestamp 1677622389
transform 1 0 3800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8376
timestamp 1677622389
transform 1 0 3808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8377
timestamp 1677622389
transform 1 0 3816 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1677622389
transform -1 0 3848 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8378
timestamp 1677622389
transform 1 0 3848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8379
timestamp 1677622389
transform 1 0 3856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8381
timestamp 1677622389
transform 1 0 3864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8383
timestamp 1677622389
transform 1 0 3872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8385
timestamp 1677622389
transform 1 0 3880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8386
timestamp 1677622389
transform 1 0 3888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8387
timestamp 1677622389
transform 1 0 3896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8388
timestamp 1677622389
transform 1 0 3904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8389
timestamp 1677622389
transform 1 0 3912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8391
timestamp 1677622389
transform 1 0 3920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8393
timestamp 1677622389
transform 1 0 3928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8402
timestamp 1677622389
transform 1 0 3936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8403
timestamp 1677622389
transform 1 0 3944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8404
timestamp 1677622389
transform 1 0 3952 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_311
timestamp 1677622389
transform -1 0 4000 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8405
timestamp 1677622389
transform 1 0 4000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8406
timestamp 1677622389
transform 1 0 4008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8407
timestamp 1677622389
transform 1 0 4016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8408
timestamp 1677622389
transform 1 0 4024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8409
timestamp 1677622389
transform 1 0 4032 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_312
timestamp 1677622389
transform -1 0 4080 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8410
timestamp 1677622389
transform 1 0 4080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8411
timestamp 1677622389
transform 1 0 4088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8412
timestamp 1677622389
transform 1 0 4096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8413
timestamp 1677622389
transform 1 0 4104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8414
timestamp 1677622389
transform 1 0 4112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8416
timestamp 1677622389
transform 1 0 4120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8418
timestamp 1677622389
transform 1 0 4128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8425
timestamp 1677622389
transform 1 0 4136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8426
timestamp 1677622389
transform 1 0 4144 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_527
timestamp 1677622389
transform -1 0 4168 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8427
timestamp 1677622389
transform 1 0 4168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8428
timestamp 1677622389
transform 1 0 4176 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_455
timestamp 1677622389
transform -1 0 4280 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8429
timestamp 1677622389
transform 1 0 4280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8430
timestamp 1677622389
transform 1 0 4288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8431
timestamp 1677622389
transform 1 0 4296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8432
timestamp 1677622389
transform 1 0 4304 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_313
timestamp 1677622389
transform 1 0 4312 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8437
timestamp 1677622389
transform 1 0 4352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8445
timestamp 1677622389
transform 1 0 4360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8446
timestamp 1677622389
transform 1 0 4368 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_531
timestamp 1677622389
transform -1 0 4392 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8447
timestamp 1677622389
transform 1 0 4392 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_458
timestamp 1677622389
transform 1 0 4400 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8448
timestamp 1677622389
transform 1 0 4496 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_147
timestamp 1677622389
transform -1 0 4536 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8449
timestamp 1677622389
transform 1 0 4536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8450
timestamp 1677622389
transform 1 0 4544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8451
timestamp 1677622389
transform 1 0 4552 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_148
timestamp 1677622389
transform -1 0 4592 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8452
timestamp 1677622389
transform 1 0 4592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8453
timestamp 1677622389
transform 1 0 4600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8454
timestamp 1677622389
transform 1 0 4608 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_315
timestamp 1677622389
transform 1 0 4616 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8455
timestamp 1677622389
transform 1 0 4656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8456
timestamp 1677622389
transform 1 0 4664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8457
timestamp 1677622389
transform 1 0 4672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8459
timestamp 1677622389
transform 1 0 4680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8461
timestamp 1677622389
transform 1 0 4688 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_316
timestamp 1677622389
transform 1 0 4696 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8462
timestamp 1677622389
transform 1 0 4736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8463
timestamp 1677622389
transform 1 0 4744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8464
timestamp 1677622389
transform 1 0 4752 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_532
timestamp 1677622389
transform -1 0 4776 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8465
timestamp 1677622389
transform 1 0 4776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8466
timestamp 1677622389
transform 1 0 4784 0 -1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_69
timestamp 1677622389
transform 1 0 4843 0 1 1270
box -10 -3 10 3
use M3_M2  M3_M2_6414
timestamp 1677622389
transform 1 0 164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6435
timestamp 1677622389
transform 1 0 132 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6436
timestamp 1677622389
transform 1 0 172 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7258
timestamp 1677622389
transform 1 0 132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7259
timestamp 1677622389
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7260
timestamp 1677622389
transform 1 0 172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7371
timestamp 1677622389
transform 1 0 84 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6415
timestamp 1677622389
transform 1 0 196 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7261
timestamp 1677622389
transform 1 0 180 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6479
timestamp 1677622389
transform 1 0 188 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7262
timestamp 1677622389
transform 1 0 204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7372
timestamp 1677622389
transform 1 0 188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7373
timestamp 1677622389
transform 1 0 196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7374
timestamp 1677622389
transform 1 0 212 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6545
timestamp 1677622389
transform 1 0 204 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7263
timestamp 1677622389
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7264
timestamp 1677622389
transform 1 0 268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7375
timestamp 1677622389
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6500
timestamp 1677622389
transform 1 0 260 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6480
timestamp 1677622389
transform 1 0 284 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7265
timestamp 1677622389
transform 1 0 292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7376
timestamp 1677622389
transform 1 0 276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7377
timestamp 1677622389
transform 1 0 284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7378
timestamp 1677622389
transform 1 0 300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7266
timestamp 1677622389
transform 1 0 316 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6481
timestamp 1677622389
transform 1 0 324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6416
timestamp 1677622389
transform 1 0 380 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6437
timestamp 1677622389
transform 1 0 372 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7267
timestamp 1677622389
transform 1 0 348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7268
timestamp 1677622389
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7269
timestamp 1677622389
transform 1 0 372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7379
timestamp 1677622389
transform 1 0 364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7380
timestamp 1677622389
transform 1 0 380 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6519
timestamp 1677622389
transform 1 0 364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6438
timestamp 1677622389
transform 1 0 404 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7270
timestamp 1677622389
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7271
timestamp 1677622389
transform 1 0 436 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6501
timestamp 1677622389
transform 1 0 436 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6417
timestamp 1677622389
transform 1 0 460 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7272
timestamp 1677622389
transform 1 0 460 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6482
timestamp 1677622389
transform 1 0 468 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7273
timestamp 1677622389
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7381
timestamp 1677622389
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7382
timestamp 1677622389
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7383
timestamp 1677622389
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6520
timestamp 1677622389
transform 1 0 484 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7274
timestamp 1677622389
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6379
timestamp 1677622389
transform 1 0 516 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6380
timestamp 1677622389
transform 1 0 548 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6392
timestamp 1677622389
transform 1 0 556 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6393
timestamp 1677622389
transform 1 0 620 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6418
timestamp 1677622389
transform 1 0 540 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6439
timestamp 1677622389
transform 1 0 524 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6440
timestamp 1677622389
transform 1 0 564 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7275
timestamp 1677622389
transform 1 0 524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7276
timestamp 1677622389
transform 1 0 564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7384
timestamp 1677622389
transform 1 0 516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6483
timestamp 1677622389
transform 1 0 572 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7277
timestamp 1677622389
transform 1 0 620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7385
timestamp 1677622389
transform 1 0 540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7386
timestamp 1677622389
transform 1 0 628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6521
timestamp 1677622389
transform 1 0 628 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6441
timestamp 1677622389
transform 1 0 652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6442
timestamp 1677622389
transform 1 0 684 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7278
timestamp 1677622389
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7279
timestamp 1677622389
transform 1 0 668 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6484
timestamp 1677622389
transform 1 0 676 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7280
timestamp 1677622389
transform 1 0 684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7387
timestamp 1677622389
transform 1 0 660 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6546
timestamp 1677622389
transform 1 0 660 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7388
timestamp 1677622389
transform 1 0 684 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6394
timestamp 1677622389
transform 1 0 700 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7389
timestamp 1677622389
transform 1 0 700 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6485
timestamp 1677622389
transform 1 0 724 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7281
timestamp 1677622389
transform 1 0 732 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6502
timestamp 1677622389
transform 1 0 716 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7390
timestamp 1677622389
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6522
timestamp 1677622389
transform 1 0 724 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7282
timestamp 1677622389
transform 1 0 748 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6503
timestamp 1677622389
transform 1 0 748 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7391
timestamp 1677622389
transform 1 0 756 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6486
timestamp 1677622389
transform 1 0 764 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6419
timestamp 1677622389
transform 1 0 804 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6443
timestamp 1677622389
transform 1 0 796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6395
timestamp 1677622389
transform 1 0 836 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6444
timestamp 1677622389
transform 1 0 820 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6445
timestamp 1677622389
transform 1 0 836 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7283
timestamp 1677622389
transform 1 0 804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7284
timestamp 1677622389
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7285
timestamp 1677622389
transform 1 0 836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7392
timestamp 1677622389
transform 1 0 796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7393
timestamp 1677622389
transform 1 0 804 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6487
timestamp 1677622389
transform 1 0 844 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6420
timestamp 1677622389
transform 1 0 860 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7286
timestamp 1677622389
transform 1 0 860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7394
timestamp 1677622389
transform 1 0 836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7395
timestamp 1677622389
transform 1 0 844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6504
timestamp 1677622389
transform 1 0 852 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6381
timestamp 1677622389
transform 1 0 916 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7287
timestamp 1677622389
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7288
timestamp 1677622389
transform 1 0 900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7289
timestamp 1677622389
transform 1 0 916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7396
timestamp 1677622389
transform 1 0 908 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7469
timestamp 1677622389
transform 1 0 924 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6547
timestamp 1677622389
transform 1 0 924 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7397
timestamp 1677622389
transform 1 0 972 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6523
timestamp 1677622389
transform 1 0 964 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7470
timestamp 1677622389
transform 1 0 972 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7290
timestamp 1677622389
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6488
timestamp 1677622389
transform 1 0 1004 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7291
timestamp 1677622389
transform 1 0 1012 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6505
timestamp 1677622389
transform 1 0 996 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7398
timestamp 1677622389
transform 1 0 1004 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6489
timestamp 1677622389
transform 1 0 1052 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7292
timestamp 1677622389
transform 1 0 1076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7399
timestamp 1677622389
transform 1 0 1028 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6524
timestamp 1677622389
transform 1 0 1028 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7293
timestamp 1677622389
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6382
timestamp 1677622389
transform 1 0 1220 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6446
timestamp 1677622389
transform 1 0 1236 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7294
timestamp 1677622389
transform 1 0 1220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7295
timestamp 1677622389
transform 1 0 1236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7400
timestamp 1677622389
transform 1 0 1212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7401
timestamp 1677622389
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7402
timestamp 1677622389
transform 1 0 1236 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6525
timestamp 1677622389
transform 1 0 1212 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6526
timestamp 1677622389
transform 1 0 1236 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7296
timestamp 1677622389
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7297
timestamp 1677622389
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6506
timestamp 1677622389
transform 1 0 1324 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7403
timestamp 1677622389
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7404
timestamp 1677622389
transform 1 0 1372 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6447
timestamp 1677622389
transform 1 0 1468 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6383
timestamp 1677622389
transform 1 0 1492 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7298
timestamp 1677622389
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7299
timestamp 1677622389
transform 1 0 1484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7405
timestamp 1677622389
transform 1 0 1404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7406
timestamp 1677622389
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6448
timestamp 1677622389
transform 1 0 1524 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7300
timestamp 1677622389
transform 1 0 1508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7301
timestamp 1677622389
transform 1 0 1524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7407
timestamp 1677622389
transform 1 0 1516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7408
timestamp 1677622389
transform 1 0 1532 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6527
timestamp 1677622389
transform 1 0 1532 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6449
timestamp 1677622389
transform 1 0 1548 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7302
timestamp 1677622389
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7409
timestamp 1677622389
transform 1 0 1548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6450
timestamp 1677622389
transform 1 0 1572 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6451
timestamp 1677622389
transform 1 0 1612 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7303
timestamp 1677622389
transform 1 0 1572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7304
timestamp 1677622389
transform 1 0 1580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7305
timestamp 1677622389
transform 1 0 1612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7306
timestamp 1677622389
transform 1 0 1676 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7410
timestamp 1677622389
transform 1 0 1660 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6528
timestamp 1677622389
transform 1 0 1580 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7411
timestamp 1677622389
transform 1 0 1692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7307
timestamp 1677622389
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7308
timestamp 1677622389
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7412
timestamp 1677622389
transform 1 0 1724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7413
timestamp 1677622389
transform 1 0 1740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7309
timestamp 1677622389
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7310
timestamp 1677622389
transform 1 0 1844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7414
timestamp 1677622389
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7311
timestamp 1677622389
transform 1 0 1892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7312
timestamp 1677622389
transform 1 0 1956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7313
timestamp 1677622389
transform 1 0 1972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7415
timestamp 1677622389
transform 1 0 1948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7416
timestamp 1677622389
transform 1 0 1964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7417
timestamp 1677622389
transform 1 0 1972 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6529
timestamp 1677622389
transform 1 0 1948 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7314
timestamp 1677622389
transform 1 0 2012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7249
timestamp 1677622389
transform 1 0 2044 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7315
timestamp 1677622389
transform 1 0 2036 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6530
timestamp 1677622389
transform 1 0 2044 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7246
timestamp 1677622389
transform 1 0 2124 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_7247
timestamp 1677622389
transform 1 0 2140 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_7250
timestamp 1677622389
transform 1 0 2132 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7418
timestamp 1677622389
transform 1 0 2132 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6548
timestamp 1677622389
transform 1 0 2140 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7316
timestamp 1677622389
transform 1 0 2172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7419
timestamp 1677622389
transform 1 0 2204 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6372
timestamp 1677622389
transform 1 0 2252 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6452
timestamp 1677622389
transform 1 0 2276 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6421
timestamp 1677622389
transform 1 0 2332 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7251
timestamp 1677622389
transform 1 0 2332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7317
timestamp 1677622389
transform 1 0 2276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7318
timestamp 1677622389
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7420
timestamp 1677622389
transform 1 0 2228 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6490
timestamp 1677622389
transform 1 0 2324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6531
timestamp 1677622389
transform 1 0 2276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6532
timestamp 1677622389
transform 1 0 2308 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6549
timestamp 1677622389
transform 1 0 2220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6396
timestamp 1677622389
transform 1 0 2356 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6453
timestamp 1677622389
transform 1 0 2348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6491
timestamp 1677622389
transform 1 0 2356 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7421
timestamp 1677622389
transform 1 0 2348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7319
timestamp 1677622389
transform 1 0 2396 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6454
timestamp 1677622389
transform 1 0 2412 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7422
timestamp 1677622389
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6550
timestamp 1677622389
transform 1 0 2412 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6422
timestamp 1677622389
transform 1 0 2436 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7320
timestamp 1677622389
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6455
timestamp 1677622389
transform 1 0 2508 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7321
timestamp 1677622389
transform 1 0 2508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7423
timestamp 1677622389
transform 1 0 2492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7322
timestamp 1677622389
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6456
timestamp 1677622389
transform 1 0 2588 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7323
timestamp 1677622389
transform 1 0 2580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7424
timestamp 1677622389
transform 1 0 2580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7471
timestamp 1677622389
transform 1 0 2572 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6551
timestamp 1677622389
transform 1 0 2580 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6397
timestamp 1677622389
transform 1 0 2636 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6423
timestamp 1677622389
transform 1 0 2604 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6424
timestamp 1677622389
transform 1 0 2628 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6384
timestamp 1677622389
transform 1 0 2668 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6385
timestamp 1677622389
transform 1 0 2684 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6398
timestamp 1677622389
transform 1 0 2756 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6457
timestamp 1677622389
transform 1 0 2628 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6458
timestamp 1677622389
transform 1 0 2652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6459
timestamp 1677622389
transform 1 0 2716 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7324
timestamp 1677622389
transform 1 0 2628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7325
timestamp 1677622389
transform 1 0 2636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7326
timestamp 1677622389
transform 1 0 2660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7327
timestamp 1677622389
transform 1 0 2716 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7425
timestamp 1677622389
transform 1 0 2604 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6533
timestamp 1677622389
transform 1 0 2604 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6552
timestamp 1677622389
transform 1 0 2612 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6507
timestamp 1677622389
transform 1 0 2716 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7426
timestamp 1677622389
transform 1 0 2740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7427
timestamp 1677622389
transform 1 0 2756 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6534
timestamp 1677622389
transform 1 0 2676 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6386
timestamp 1677622389
transform 1 0 2868 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6399
timestamp 1677622389
transform 1 0 2772 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6400
timestamp 1677622389
transform 1 0 2844 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6425
timestamp 1677622389
transform 1 0 2788 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7328
timestamp 1677622389
transform 1 0 2772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7329
timestamp 1677622389
transform 1 0 2780 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6492
timestamp 1677622389
transform 1 0 2868 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6387
timestamp 1677622389
transform 1 0 2900 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6426
timestamp 1677622389
transform 1 0 2892 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7428
timestamp 1677622389
transform 1 0 2876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7429
timestamp 1677622389
transform 1 0 2884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7472
timestamp 1677622389
transform 1 0 2868 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6401
timestamp 1677622389
transform 1 0 3004 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7330
timestamp 1677622389
transform 1 0 2996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7331
timestamp 1677622389
transform 1 0 3004 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6508
timestamp 1677622389
transform 1 0 3004 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6402
timestamp 1677622389
transform 1 0 3036 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7252
timestamp 1677622389
transform 1 0 3036 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7430
timestamp 1677622389
transform 1 0 3012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7431
timestamp 1677622389
transform 1 0 3020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7473
timestamp 1677622389
transform 1 0 2908 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6553
timestamp 1677622389
transform 1 0 2908 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6554
timestamp 1677622389
transform 1 0 3020 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6403
timestamp 1677622389
transform 1 0 3060 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7253
timestamp 1677622389
transform 1 0 3052 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6373
timestamp 1677622389
transform 1 0 3092 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6427
timestamp 1677622389
transform 1 0 3084 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6460
timestamp 1677622389
transform 1 0 3076 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7332
timestamp 1677622389
transform 1 0 3076 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6374
timestamp 1677622389
transform 1 0 3124 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6404
timestamp 1677622389
transform 1 0 3116 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7248
timestamp 1677622389
transform 1 0 3108 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_6461
timestamp 1677622389
transform 1 0 3100 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7333
timestamp 1677622389
transform 1 0 3100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7254
timestamp 1677622389
transform 1 0 3116 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7432
timestamp 1677622389
transform 1 0 3124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7255
timestamp 1677622389
transform 1 0 3156 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6428
timestamp 1677622389
transform 1 0 3188 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7433
timestamp 1677622389
transform 1 0 3188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7434
timestamp 1677622389
transform 1 0 3196 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6535
timestamp 1677622389
transform 1 0 3196 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7435
timestamp 1677622389
transform 1 0 3212 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6375
timestamp 1677622389
transform 1 0 3244 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6388
timestamp 1677622389
transform 1 0 3236 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6376
timestamp 1677622389
transform 1 0 3276 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6389
timestamp 1677622389
transform 1 0 3276 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6405
timestamp 1677622389
transform 1 0 3260 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6462
timestamp 1677622389
transform 1 0 3228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6463
timestamp 1677622389
transform 1 0 3252 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7334
timestamp 1677622389
transform 1 0 3228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7335
timestamp 1677622389
transform 1 0 3236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7336
timestamp 1677622389
transform 1 0 3244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7337
timestamp 1677622389
transform 1 0 3260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7436
timestamp 1677622389
transform 1 0 3244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7437
timestamp 1677622389
transform 1 0 3252 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6555
timestamp 1677622389
transform 1 0 3236 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7438
timestamp 1677622389
transform 1 0 3300 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6390
timestamp 1677622389
transform 1 0 3340 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6406
timestamp 1677622389
transform 1 0 3332 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6429
timestamp 1677622389
transform 1 0 3316 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7338
timestamp 1677622389
transform 1 0 3308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7339
timestamp 1677622389
transform 1 0 3316 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6509
timestamp 1677622389
transform 1 0 3308 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6391
timestamp 1677622389
transform 1 0 3380 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6407
timestamp 1677622389
transform 1 0 3364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6430
timestamp 1677622389
transform 1 0 3356 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6431
timestamp 1677622389
transform 1 0 3412 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6464
timestamp 1677622389
transform 1 0 3348 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7439
timestamp 1677622389
transform 1 0 3316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7440
timestamp 1677622389
transform 1 0 3332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7340
timestamp 1677622389
transform 1 0 3348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6556
timestamp 1677622389
transform 1 0 3340 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6465
timestamp 1677622389
transform 1 0 3460 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7341
timestamp 1677622389
transform 1 0 3452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7342
timestamp 1677622389
transform 1 0 3460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7441
timestamp 1677622389
transform 1 0 3356 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6510
timestamp 1677622389
transform 1 0 3364 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7442
timestamp 1677622389
transform 1 0 3468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7474
timestamp 1677622389
transform 1 0 3364 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6536
timestamp 1677622389
transform 1 0 3468 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6408
timestamp 1677622389
transform 1 0 3572 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6466
timestamp 1677622389
transform 1 0 3540 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7343
timestamp 1677622389
transform 1 0 3484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7344
timestamp 1677622389
transform 1 0 3540 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6493
timestamp 1677622389
transform 1 0 3564 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6511
timestamp 1677622389
transform 1 0 3484 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6512
timestamp 1677622389
transform 1 0 3540 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7443
timestamp 1677622389
transform 1 0 3564 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6409
timestamp 1677622389
transform 1 0 3588 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6467
timestamp 1677622389
transform 1 0 3620 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7345
timestamp 1677622389
transform 1 0 3612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7346
timestamp 1677622389
transform 1 0 3628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7444
timestamp 1677622389
transform 1 0 3604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7445
timestamp 1677622389
transform 1 0 3620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6557
timestamp 1677622389
transform 1 0 3604 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6558
timestamp 1677622389
transform 1 0 3628 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6494
timestamp 1677622389
transform 1 0 3676 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7446
timestamp 1677622389
transform 1 0 3676 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6468
timestamp 1677622389
transform 1 0 3692 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7347
timestamp 1677622389
transform 1 0 3740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7447
timestamp 1677622389
transform 1 0 3692 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6513
timestamp 1677622389
transform 1 0 3740 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6559
timestamp 1677622389
transform 1 0 3764 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7348
timestamp 1677622389
transform 1 0 3780 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6432
timestamp 1677622389
transform 1 0 3796 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7349
timestamp 1677622389
transform 1 0 3804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7448
timestamp 1677622389
transform 1 0 3796 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6560
timestamp 1677622389
transform 1 0 3796 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6433
timestamp 1677622389
transform 1 0 3836 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7350
timestamp 1677622389
transform 1 0 3836 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6495
timestamp 1677622389
transform 1 0 3844 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7351
timestamp 1677622389
transform 1 0 3852 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6514
timestamp 1677622389
transform 1 0 3820 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7449
timestamp 1677622389
transform 1 0 3828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7450
timestamp 1677622389
transform 1 0 3844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6537
timestamp 1677622389
transform 1 0 3852 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6561
timestamp 1677622389
transform 1 0 3844 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6496
timestamp 1677622389
transform 1 0 3868 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7451
timestamp 1677622389
transform 1 0 3868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7256
timestamp 1677622389
transform 1 0 3908 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6538
timestamp 1677622389
transform 1 0 3916 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6469
timestamp 1677622389
transform 1 0 3940 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7352
timestamp 1677622389
transform 1 0 3964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7353
timestamp 1677622389
transform 1 0 4020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7354
timestamp 1677622389
transform 1 0 4028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7452
timestamp 1677622389
transform 1 0 3940 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6515
timestamp 1677622389
transform 1 0 3972 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6539
timestamp 1677622389
transform 1 0 3964 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6562
timestamp 1677622389
transform 1 0 3932 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7355
timestamp 1677622389
transform 1 0 4052 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6540
timestamp 1677622389
transform 1 0 4060 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6470
timestamp 1677622389
transform 1 0 4084 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7356
timestamp 1677622389
transform 1 0 4108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7357
timestamp 1677622389
transform 1 0 4164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7453
timestamp 1677622389
transform 1 0 4084 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6541
timestamp 1677622389
transform 1 0 4108 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6410
timestamp 1677622389
transform 1 0 4244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6471
timestamp 1677622389
transform 1 0 4196 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6472
timestamp 1677622389
transform 1 0 4268 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7358
timestamp 1677622389
transform 1 0 4236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7454
timestamp 1677622389
transform 1 0 4196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7359
timestamp 1677622389
transform 1 0 4300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7360
timestamp 1677622389
transform 1 0 4324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7455
timestamp 1677622389
transform 1 0 4316 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6411
timestamp 1677622389
transform 1 0 4340 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7456
timestamp 1677622389
transform 1 0 4332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6542
timestamp 1677622389
transform 1 0 4332 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6473
timestamp 1677622389
transform 1 0 4372 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7361
timestamp 1677622389
transform 1 0 4372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7362
timestamp 1677622389
transform 1 0 4388 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6516
timestamp 1677622389
transform 1 0 4372 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6377
timestamp 1677622389
transform 1 0 4412 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_7457
timestamp 1677622389
transform 1 0 4380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7458
timestamp 1677622389
transform 1 0 4396 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6517
timestamp 1677622389
transform 1 0 4404 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6474
timestamp 1677622389
transform 1 0 4420 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6412
timestamp 1677622389
transform 1 0 4444 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6518
timestamp 1677622389
transform 1 0 4436 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7363
timestamp 1677622389
transform 1 0 4468 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6475
timestamp 1677622389
transform 1 0 4476 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6413
timestamp 1677622389
transform 1 0 4500 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6476
timestamp 1677622389
transform 1 0 4516 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7364
timestamp 1677622389
transform 1 0 4508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7365
timestamp 1677622389
transform 1 0 4524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7459
timestamp 1677622389
transform 1 0 4492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7460
timestamp 1677622389
transform 1 0 4500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7461
timestamp 1677622389
transform 1 0 4516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6563
timestamp 1677622389
transform 1 0 4500 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7462
timestamp 1677622389
transform 1 0 4540 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6497
timestamp 1677622389
transform 1 0 4548 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7463
timestamp 1677622389
transform 1 0 4548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7257
timestamp 1677622389
transform 1 0 4564 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_6498
timestamp 1677622389
transform 1 0 4564 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7366
timestamp 1677622389
transform 1 0 4588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7367
timestamp 1677622389
transform 1 0 4596 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6564
timestamp 1677622389
transform 1 0 4588 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6499
timestamp 1677622389
transform 1 0 4612 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7464
timestamp 1677622389
transform 1 0 4604 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6434
timestamp 1677622389
transform 1 0 4644 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6477
timestamp 1677622389
transform 1 0 4636 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7368
timestamp 1677622389
transform 1 0 4644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7465
timestamp 1677622389
transform 1 0 4620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7466
timestamp 1677622389
transform 1 0 4636 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7467
timestamp 1677622389
transform 1 0 4652 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6543
timestamp 1677622389
transform 1 0 4652 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6378
timestamp 1677622389
transform 1 0 4700 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6478
timestamp 1677622389
transform 1 0 4724 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7369
timestamp 1677622389
transform 1 0 4724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7370
timestamp 1677622389
transform 1 0 4780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7468
timestamp 1677622389
transform 1 0 4700 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6544
timestamp 1677622389
transform 1 0 4716 0 1 1195
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_70
timestamp 1677622389
transform 1 0 48 0 1 1170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_460
timestamp 1677622389
transform 1 0 72 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_533
timestamp 1677622389
transform -1 0 184 0 1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_310
timestamp 1677622389
transform -1 0 224 0 1 1170
box -8 -3 46 105
use FILL  FILL_8467
timestamp 1677622389
transform 1 0 224 0 1 1170
box -8 -3 16 105
use FILL  FILL_8468
timestamp 1677622389
transform 1 0 232 0 1 1170
box -8 -3 16 105
use FILL  FILL_8469
timestamp 1677622389
transform 1 0 240 0 1 1170
box -8 -3 16 105
use FILL  FILL_8470
timestamp 1677622389
transform 1 0 248 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_534
timestamp 1677622389
transform -1 0 272 0 1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_311
timestamp 1677622389
transform 1 0 272 0 1 1170
box -8 -3 46 105
use FILL  FILL_8471
timestamp 1677622389
transform 1 0 312 0 1 1170
box -8 -3 16 105
use FILL  FILL_8479
timestamp 1677622389
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_8481
timestamp 1677622389
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8483
timestamp 1677622389
transform 1 0 336 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_317
timestamp 1677622389
transform 1 0 344 0 1 1170
box -8 -3 46 105
use FILL  FILL_8485
timestamp 1677622389
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_8486
timestamp 1677622389
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_8487
timestamp 1677622389
transform 1 0 400 0 1 1170
box -8 -3 16 105
use FILL  FILL_8488
timestamp 1677622389
transform 1 0 408 0 1 1170
box -8 -3 16 105
use FILL  FILL_8489
timestamp 1677622389
transform 1 0 416 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_535
timestamp 1677622389
transform -1 0 440 0 1 1170
box -9 -3 26 105
use FILL  FILL_8490
timestamp 1677622389
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8491
timestamp 1677622389
transform 1 0 448 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_312
timestamp 1677622389
transform 1 0 456 0 1 1170
box -8 -3 46 105
use FILL  FILL_8492
timestamp 1677622389
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_8493
timestamp 1677622389
transform 1 0 504 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_536
timestamp 1677622389
transform 1 0 512 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_463
timestamp 1677622389
transform 1 0 528 0 1 1170
box -8 -3 104 105
use FILL  FILL_8494
timestamp 1677622389
transform 1 0 624 0 1 1170
box -8 -3 16 105
use FILL  FILL_8495
timestamp 1677622389
transform 1 0 632 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_318
timestamp 1677622389
transform 1 0 640 0 1 1170
box -8 -3 46 105
use FILL  FILL_8496
timestamp 1677622389
transform 1 0 680 0 1 1170
box -8 -3 16 105
use FILL  FILL_8497
timestamp 1677622389
transform 1 0 688 0 1 1170
box -8 -3 16 105
use FILL  FILL_8498
timestamp 1677622389
transform 1 0 696 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_319
timestamp 1677622389
transform 1 0 704 0 1 1170
box -8 -3 46 105
use FILL  FILL_8499
timestamp 1677622389
transform 1 0 744 0 1 1170
box -8 -3 16 105
use FILL  FILL_8500
timestamp 1677622389
transform 1 0 752 0 1 1170
box -8 -3 16 105
use FILL  FILL_8510
timestamp 1677622389
transform 1 0 760 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6565
timestamp 1677622389
transform 1 0 780 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_538
timestamp 1677622389
transform -1 0 784 0 1 1170
box -9 -3 26 105
use FILL  FILL_8511
timestamp 1677622389
transform 1 0 784 0 1 1170
box -8 -3 16 105
use FILL  FILL_8512
timestamp 1677622389
transform 1 0 792 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_314
timestamp 1677622389
transform -1 0 840 0 1 1170
box -8 -3 46 105
use FILL  FILL_8513
timestamp 1677622389
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_8514
timestamp 1677622389
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8515
timestamp 1677622389
transform 1 0 856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8516
timestamp 1677622389
transform 1 0 864 0 1 1170
box -8 -3 16 105
use FILL  FILL_8519
timestamp 1677622389
transform 1 0 872 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_315
timestamp 1677622389
transform -1 0 920 0 1 1170
box -8 -3 46 105
use FILL  FILL_8520
timestamp 1677622389
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_8526
timestamp 1677622389
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_8527
timestamp 1677622389
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_8528
timestamp 1677622389
transform 1 0 944 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_85
timestamp 1677622389
transform 1 0 952 0 1 1170
box -8 -3 32 105
use FILL  FILL_8529
timestamp 1677622389
transform 1 0 976 0 1 1170
box -8 -3 16 105
use FILL  FILL_8534
timestamp 1677622389
transform 1 0 984 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_87
timestamp 1677622389
transform 1 0 992 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_6566
timestamp 1677622389
transform 1 0 1052 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_468
timestamp 1677622389
transform 1 0 1016 0 1 1170
box -8 -3 104 105
use FILL  FILL_8536
timestamp 1677622389
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8550
timestamp 1677622389
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_8552
timestamp 1677622389
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use FILL  FILL_8553
timestamp 1677622389
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_8554
timestamp 1677622389
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_8555
timestamp 1677622389
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8558
timestamp 1677622389
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8560
timestamp 1677622389
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8562
timestamp 1677622389
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8564
timestamp 1677622389
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8566
timestamp 1677622389
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_316
timestamp 1677622389
transform -1 0 1240 0 1 1170
box -8 -3 46 105
use FILL  FILL_8567
timestamp 1677622389
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_8575
timestamp 1677622389
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_8577
timestamp 1677622389
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_8579
timestamp 1677622389
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_8581
timestamp 1677622389
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_8583
timestamp 1677622389
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_8584
timestamp 1677622389
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8585
timestamp 1677622389
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8586
timestamp 1677622389
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_320
timestamp 1677622389
transform -1 0 1352 0 1 1170
box -8 -3 46 105
use FILL  FILL_8587
timestamp 1677622389
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_8588
timestamp 1677622389
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_8589
timestamp 1677622389
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_8590
timestamp 1677622389
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_8592
timestamp 1677622389
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_470
timestamp 1677622389
transform 1 0 1392 0 1 1170
box -8 -3 104 105
use FILL  FILL_8593
timestamp 1677622389
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_8594
timestamp 1677622389
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_317
timestamp 1677622389
transform 1 0 1504 0 1 1170
box -8 -3 46 105
use FILL  FILL_8595
timestamp 1677622389
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_541
timestamp 1677622389
transform 1 0 1552 0 1 1170
box -9 -3 26 105
use FILL  FILL_8596
timestamp 1677622389
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_471
timestamp 1677622389
transform -1 0 1672 0 1 1170
box -8 -3 104 105
use BUFX2  BUFX2_104
timestamp 1677622389
transform 1 0 1672 0 1 1170
box -5 -3 28 105
use FILL  FILL_8597
timestamp 1677622389
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_8607
timestamp 1677622389
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_8608
timestamp 1677622389
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_321
timestamp 1677622389
transform 1 0 1720 0 1 1170
box -8 -3 46 105
use FILL  FILL_8609
timestamp 1677622389
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_8610
timestamp 1677622389
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8611
timestamp 1677622389
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_474
timestamp 1677622389
transform -1 0 1880 0 1 1170
box -8 -3 104 105
use FILL  FILL_8612
timestamp 1677622389
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_8613
timestamp 1677622389
transform 1 0 1888 0 1 1170
box -8 -3 16 105
use FILL  FILL_8614
timestamp 1677622389
transform 1 0 1896 0 1 1170
box -8 -3 16 105
use FILL  FILL_8615
timestamp 1677622389
transform 1 0 1904 0 1 1170
box -8 -3 16 105
use FILL  FILL_8616
timestamp 1677622389
transform 1 0 1912 0 1 1170
box -8 -3 16 105
use FILL  FILL_8617
timestamp 1677622389
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_8618
timestamp 1677622389
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_319
timestamp 1677622389
transform 1 0 1936 0 1 1170
box -8 -3 46 105
use FILL  FILL_8619
timestamp 1677622389
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_8620
timestamp 1677622389
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_8636
timestamp 1677622389
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_8638
timestamp 1677622389
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_8640
timestamp 1677622389
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use FILL  FILL_8641
timestamp 1677622389
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_545
timestamp 1677622389
transform 1 0 2024 0 1 1170
box -9 -3 26 105
use FILL  FILL_8642
timestamp 1677622389
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8643
timestamp 1677622389
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_8644
timestamp 1677622389
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_8647
timestamp 1677622389
transform 1 0 2064 0 1 1170
box -8 -3 16 105
use FILL  FILL_8648
timestamp 1677622389
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_8649
timestamp 1677622389
transform 1 0 2080 0 1 1170
box -8 -3 16 105
use FILL  FILL_8650
timestamp 1677622389
transform 1 0 2088 0 1 1170
box -8 -3 16 105
use FILL  FILL_8653
timestamp 1677622389
transform 1 0 2096 0 1 1170
box -8 -3 16 105
use FILL  FILL_8655
timestamp 1677622389
transform 1 0 2104 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1677622389
transform -1 0 2144 0 1 1170
box -8 -3 40 105
use FILL  FILL_8656
timestamp 1677622389
transform 1 0 2144 0 1 1170
box -8 -3 16 105
use FILL  FILL_8657
timestamp 1677622389
transform 1 0 2152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8658
timestamp 1677622389
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_547
timestamp 1677622389
transform -1 0 2184 0 1 1170
box -9 -3 26 105
use FILL  FILL_8659
timestamp 1677622389
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8667
timestamp 1677622389
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8669
timestamp 1677622389
transform 1 0 2200 0 1 1170
box -8 -3 16 105
use FILL  FILL_8670
timestamp 1677622389
transform 1 0 2208 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_476
timestamp 1677622389
transform 1 0 2216 0 1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_16
timestamp 1677622389
transform 1 0 2312 0 1 1170
box -8 -3 32 105
use FILL  FILL_8671
timestamp 1677622389
transform 1 0 2336 0 1 1170
box -8 -3 16 105
use FILL  FILL_8672
timestamp 1677622389
transform 1 0 2344 0 1 1170
box -8 -3 16 105
use FILL  FILL_8673
timestamp 1677622389
transform 1 0 2352 0 1 1170
box -8 -3 16 105
use FILL  FILL_8674
timestamp 1677622389
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_8675
timestamp 1677622389
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_149
timestamp 1677622389
transform -1 0 2408 0 1 1170
box -8 -3 34 105
use FILL  FILL_8676
timestamp 1677622389
transform 1 0 2408 0 1 1170
box -8 -3 16 105
use FILL  FILL_8688
timestamp 1677622389
transform 1 0 2416 0 1 1170
box -8 -3 16 105
use FILL  FILL_8689
timestamp 1677622389
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_8690
timestamp 1677622389
transform 1 0 2432 0 1 1170
box -8 -3 16 105
use FILL  FILL_8691
timestamp 1677622389
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8692
timestamp 1677622389
transform 1 0 2448 0 1 1170
box -8 -3 16 105
use FILL  FILL_8693
timestamp 1677622389
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_8694
timestamp 1677622389
transform 1 0 2464 0 1 1170
box -8 -3 16 105
use FILL  FILL_8695
timestamp 1677622389
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_10
timestamp 1677622389
transform 1 0 2480 0 1 1170
box -7 -3 39 105
use FILL  FILL_8696
timestamp 1677622389
transform 1 0 2512 0 1 1170
box -8 -3 16 105
use FILL  FILL_8697
timestamp 1677622389
transform 1 0 2520 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_548
timestamp 1677622389
transform -1 0 2544 0 1 1170
box -9 -3 26 105
use FILL  FILL_8698
timestamp 1677622389
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_8699
timestamp 1677622389
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_8700
timestamp 1677622389
transform 1 0 2560 0 1 1170
box -8 -3 16 105
use FILL  FILL_8701
timestamp 1677622389
transform 1 0 2568 0 1 1170
box -8 -3 16 105
use FILL  FILL_8702
timestamp 1677622389
transform 1 0 2576 0 1 1170
box -8 -3 16 105
use FILL  FILL_8705
timestamp 1677622389
transform 1 0 2584 0 1 1170
box -8 -3 16 105
use FILL  FILL_8707
timestamp 1677622389
transform 1 0 2592 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6567
timestamp 1677622389
transform 1 0 2620 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6568
timestamp 1677622389
transform 1 0 2708 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_1
timestamp 1677622389
transform 1 0 2600 0 1 1170
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_478
timestamp 1677622389
transform -1 0 2752 0 1 1170
box -8 -3 104 105
use FILL  FILL_8708
timestamp 1677622389
transform 1 0 2752 0 1 1170
box -8 -3 16 105
use FAX1  FAX1_10
timestamp 1677622389
transform 1 0 2760 0 1 1170
box -5 -3 126 105
use FILL  FILL_8709
timestamp 1677622389
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_8715
timestamp 1677622389
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FAX1  FAX1_12
timestamp 1677622389
transform -1 0 3016 0 1 1170
box -5 -3 126 105
use NAND2X1  NAND2X1_17
timestamp 1677622389
transform 1 0 3016 0 1 1170
box -8 -3 32 105
use FILL  FILL_8717
timestamp 1677622389
transform 1 0 3040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8719
timestamp 1677622389
transform 1 0 3048 0 1 1170
box -8 -3 16 105
use FILL  FILL_8721
timestamp 1677622389
transform 1 0 3056 0 1 1170
box -8 -3 16 105
use FILL  FILL_8723
timestamp 1677622389
transform 1 0 3064 0 1 1170
box -8 -3 16 105
use FILL  FILL_8725
timestamp 1677622389
transform 1 0 3072 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_67
timestamp 1677622389
transform -1 0 3112 0 1 1170
box -8 -3 40 105
use FILL  FILL_8726
timestamp 1677622389
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8727
timestamp 1677622389
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_8728
timestamp 1677622389
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_8729
timestamp 1677622389
transform 1 0 3136 0 1 1170
box -8 -3 16 105
use FILL  FILL_8733
timestamp 1677622389
transform 1 0 3144 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_151
timestamp 1677622389
transform -1 0 3184 0 1 1170
box -8 -3 34 105
use FILL  FILL_8734
timestamp 1677622389
transform 1 0 3184 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_550
timestamp 1677622389
transform 1 0 3192 0 1 1170
box -9 -3 26 105
use FILL  FILL_8735
timestamp 1677622389
transform 1 0 3208 0 1 1170
box -8 -3 16 105
use FILL  FILL_8741
timestamp 1677622389
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6569
timestamp 1677622389
transform 1 0 3236 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_551
timestamp 1677622389
transform 1 0 3224 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_6570
timestamp 1677622389
transform 1 0 3284 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_323
timestamp 1677622389
transform 1 0 3240 0 1 1170
box -8 -3 46 105
use FILL  FILL_8742
timestamp 1677622389
transform 1 0 3280 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6571
timestamp 1677622389
transform 1 0 3300 0 1 1175
box -3 -3 3 3
use FILL  FILL_8747
timestamp 1677622389
transform 1 0 3288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8749
timestamp 1677622389
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8751
timestamp 1677622389
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_12
timestamp 1677622389
transform -1 0 3344 0 1 1170
box -7 -3 39 105
use FILL  FILL_8752
timestamp 1677622389
transform 1 0 3344 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6572
timestamp 1677622389
transform 1 0 3364 0 1 1175
box -3 -3 3 3
use FAX1  FAX1_14
timestamp 1677622389
transform -1 0 3472 0 1 1170
box -5 -3 126 105
use FILL  FILL_8753
timestamp 1677622389
transform 1 0 3472 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_480
timestamp 1677622389
transform -1 0 3576 0 1 1170
box -8 -3 104 105
use FILL  FILL_8754
timestamp 1677622389
transform 1 0 3576 0 1 1170
box -8 -3 16 105
use FILL  FILL_8764
timestamp 1677622389
transform 1 0 3584 0 1 1170
box -8 -3 16 105
use FILL  FILL_8765
timestamp 1677622389
transform 1 0 3592 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_322
timestamp 1677622389
transform 1 0 3600 0 1 1170
box -8 -3 46 105
use FILL  FILL_8766
timestamp 1677622389
transform 1 0 3640 0 1 1170
box -8 -3 16 105
use FILL  FILL_8770
timestamp 1677622389
transform 1 0 3648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8772
timestamp 1677622389
transform 1 0 3656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8774
timestamp 1677622389
transform 1 0 3664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8776
timestamp 1677622389
transform 1 0 3672 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_481
timestamp 1677622389
transform 1 0 3680 0 1 1170
box -8 -3 104 105
use FILL  FILL_8777
timestamp 1677622389
transform 1 0 3776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8785
timestamp 1677622389
transform 1 0 3784 0 1 1170
box -8 -3 16 105
use FILL  FILL_8787
timestamp 1677622389
transform 1 0 3792 0 1 1170
box -8 -3 16 105
use FILL  FILL_8789
timestamp 1677622389
transform 1 0 3800 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_325
timestamp 1677622389
transform 1 0 3808 0 1 1170
box -8 -3 46 105
use FILL  FILL_8791
timestamp 1677622389
transform 1 0 3848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8798
timestamp 1677622389
transform 1 0 3856 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_19
timestamp 1677622389
transform 1 0 3864 0 1 1170
box -8 -3 32 105
use FILL  FILL_8800
timestamp 1677622389
transform 1 0 3888 0 1 1170
box -8 -3 16 105
use FILL  FILL_8805
timestamp 1677622389
transform 1 0 3896 0 1 1170
box -8 -3 16 105
use FILL  FILL_8806
timestamp 1677622389
transform 1 0 3904 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6573
timestamp 1677622389
transform 1 0 3924 0 1 1175
box -3 -3 3 3
use FILL  FILL_8807
timestamp 1677622389
transform 1 0 3912 0 1 1170
box -8 -3 16 105
use FILL  FILL_8808
timestamp 1677622389
transform 1 0 3920 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6574
timestamp 1677622389
transform 1 0 3956 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_482
timestamp 1677622389
transform 1 0 3928 0 1 1170
box -8 -3 104 105
use FILL  FILL_8809
timestamp 1677622389
transform 1 0 4024 0 1 1170
box -8 -3 16 105
use FILL  FILL_8820
timestamp 1677622389
transform 1 0 4032 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_557
timestamp 1677622389
transform -1 0 4056 0 1 1170
box -9 -3 26 105
use FILL  FILL_8821
timestamp 1677622389
transform 1 0 4056 0 1 1170
box -8 -3 16 105
use FILL  FILL_8822
timestamp 1677622389
transform 1 0 4064 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_483
timestamp 1677622389
transform 1 0 4072 0 1 1170
box -8 -3 104 105
use FILL  FILL_8823
timestamp 1677622389
transform 1 0 4168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8835
timestamp 1677622389
transform 1 0 4176 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6575
timestamp 1677622389
transform 1 0 4196 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_484
timestamp 1677622389
transform 1 0 4184 0 1 1170
box -8 -3 104 105
use FILL  FILL_8837
timestamp 1677622389
transform 1 0 4280 0 1 1170
box -8 -3 16 105
use FILL  FILL_8846
timestamp 1677622389
transform 1 0 4288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8848
timestamp 1677622389
transform 1 0 4296 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_559
timestamp 1677622389
transform -1 0 4320 0 1 1170
box -9 -3 26 105
use FILL  FILL_8849
timestamp 1677622389
transform 1 0 4320 0 1 1170
box -8 -3 16 105
use FILL  FILL_8850
timestamp 1677622389
transform 1 0 4328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8851
timestamp 1677622389
transform 1 0 4336 0 1 1170
box -8 -3 16 105
use FILL  FILL_8852
timestamp 1677622389
transform 1 0 4344 0 1 1170
box -8 -3 16 105
use FILL  FILL_8855
timestamp 1677622389
transform 1 0 4352 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6576
timestamp 1677622389
transform 1 0 4396 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_330
timestamp 1677622389
transform -1 0 4400 0 1 1170
box -8 -3 46 105
use FILL  FILL_8856
timestamp 1677622389
transform 1 0 4400 0 1 1170
box -8 -3 16 105
use FILL  FILL_8857
timestamp 1677622389
transform 1 0 4408 0 1 1170
box -8 -3 16 105
use FILL  FILL_8858
timestamp 1677622389
transform 1 0 4416 0 1 1170
box -8 -3 16 105
use FILL  FILL_8859
timestamp 1677622389
transform 1 0 4424 0 1 1170
box -8 -3 16 105
use FILL  FILL_8865
timestamp 1677622389
transform 1 0 4432 0 1 1170
box -8 -3 16 105
use FILL  FILL_8867
timestamp 1677622389
transform 1 0 4440 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_560
timestamp 1677622389
transform -1 0 4464 0 1 1170
box -9 -3 26 105
use FILL  FILL_8868
timestamp 1677622389
transform 1 0 4464 0 1 1170
box -8 -3 16 105
use FILL  FILL_8873
timestamp 1677622389
transform 1 0 4472 0 1 1170
box -8 -3 16 105
use FILL  FILL_8874
timestamp 1677622389
transform 1 0 4480 0 1 1170
box -8 -3 16 105
use FILL  FILL_8875
timestamp 1677622389
transform 1 0 4488 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_332
timestamp 1677622389
transform 1 0 4496 0 1 1170
box -8 -3 46 105
use FILL  FILL_8876
timestamp 1677622389
transform 1 0 4536 0 1 1170
box -8 -3 16 105
use FILL  FILL_8881
timestamp 1677622389
transform 1 0 4544 0 1 1170
box -8 -3 16 105
use FILL  FILL_8882
timestamp 1677622389
transform 1 0 4552 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_152
timestamp 1677622389
transform -1 0 4592 0 1 1170
box -8 -3 34 105
use FILL  FILL_8883
timestamp 1677622389
transform 1 0 4592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8886
timestamp 1677622389
transform 1 0 4600 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6577
timestamp 1677622389
transform 1 0 4620 0 1 1175
box -3 -3 3 3
use FILL  FILL_8888
timestamp 1677622389
transform 1 0 4608 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6578
timestamp 1677622389
transform 1 0 4660 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_335
timestamp 1677622389
transform 1 0 4616 0 1 1170
box -8 -3 46 105
use FILL  FILL_8890
timestamp 1677622389
transform 1 0 4656 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6579
timestamp 1677622389
transform 1 0 4676 0 1 1175
box -3 -3 3 3
use FILL  FILL_8891
timestamp 1677622389
transform 1 0 4664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8892
timestamp 1677622389
transform 1 0 4672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8896
timestamp 1677622389
transform 1 0 4680 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_485
timestamp 1677622389
transform 1 0 4688 0 1 1170
box -8 -3 104 105
use FILL  FILL_8897
timestamp 1677622389
transform 1 0 4784 0 1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_71
timestamp 1677622389
transform 1 0 4819 0 1 1170
box -10 -3 10 3
use M2_M1  M2_M1_7482
timestamp 1677622389
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7573
timestamp 1677622389
transform 1 0 108 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6699
timestamp 1677622389
transform 1 0 84 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6700
timestamp 1677622389
transform 1 0 108 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7574
timestamp 1677622389
transform 1 0 172 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6580
timestamp 1677622389
transform 1 0 188 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6581
timestamp 1677622389
transform 1 0 212 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7483
timestamp 1677622389
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7575
timestamp 1677622389
transform 1 0 236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7576
timestamp 1677622389
transform 1 0 308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6633
timestamp 1677622389
transform 1 0 444 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7484
timestamp 1677622389
transform 1 0 444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7577
timestamp 1677622389
transform 1 0 364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7578
timestamp 1677622389
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6582
timestamp 1677622389
transform 1 0 484 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6583
timestamp 1677622389
transform 1 0 540 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6634
timestamp 1677622389
transform 1 0 484 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6635
timestamp 1677622389
transform 1 0 564 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6636
timestamp 1677622389
transform 1 0 596 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7485
timestamp 1677622389
transform 1 0 484 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6668
timestamp 1677622389
transform 1 0 532 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7486
timestamp 1677622389
transform 1 0 572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7487
timestamp 1677622389
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6669
timestamp 1677622389
transform 1 0 612 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7579
timestamp 1677622389
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7580
timestamp 1677622389
transform 1 0 564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7581
timestamp 1677622389
transform 1 0 572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7582
timestamp 1677622389
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7583
timestamp 1677622389
transform 1 0 604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7584
timestamp 1677622389
transform 1 0 612 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6701
timestamp 1677622389
transform 1 0 588 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6736
timestamp 1677622389
transform 1 0 580 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6737
timestamp 1677622389
transform 1 0 612 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6637
timestamp 1677622389
transform 1 0 644 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7488
timestamp 1677622389
transform 1 0 636 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6702
timestamp 1677622389
transform 1 0 636 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6584
timestamp 1677622389
transform 1 0 660 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6585
timestamp 1677622389
transform 1 0 684 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6610
timestamp 1677622389
transform 1 0 692 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7489
timestamp 1677622389
transform 1 0 740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7585
timestamp 1677622389
transform 1 0 660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7586
timestamp 1677622389
transform 1 0 716 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6779
timestamp 1677622389
transform 1 0 684 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7587
timestamp 1677622389
transform 1 0 764 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6586
timestamp 1677622389
transform 1 0 804 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6587
timestamp 1677622389
transform 1 0 836 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6670
timestamp 1677622389
transform 1 0 820 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7490
timestamp 1677622389
transform 1 0 852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7588
timestamp 1677622389
transform 1 0 820 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6588
timestamp 1677622389
transform 1 0 868 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6671
timestamp 1677622389
transform 1 0 868 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7589
timestamp 1677622389
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6767
timestamp 1677622389
transform 1 0 868 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6768
timestamp 1677622389
transform 1 0 884 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7491
timestamp 1677622389
transform 1 0 900 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6589
timestamp 1677622389
transform 1 0 908 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7475
timestamp 1677622389
transform 1 0 908 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6780
timestamp 1677622389
transform 1 0 908 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7476
timestamp 1677622389
transform 1 0 948 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7492
timestamp 1677622389
transform 1 0 940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7590
timestamp 1677622389
transform 1 0 1060 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6738
timestamp 1677622389
transform 1 0 1060 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7591
timestamp 1677622389
transform 1 0 1076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7592
timestamp 1677622389
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6703
timestamp 1677622389
transform 1 0 1084 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7493
timestamp 1677622389
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6704
timestamp 1677622389
transform 1 0 1196 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7494
timestamp 1677622389
transform 1 0 1220 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6739
timestamp 1677622389
transform 1 0 1220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6638
timestamp 1677622389
transform 1 0 1236 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6590
timestamp 1677622389
transform 1 0 1292 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6591
timestamp 1677622389
transform 1 0 1356 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6639
timestamp 1677622389
transform 1 0 1340 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7495
timestamp 1677622389
transform 1 0 1292 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6672
timestamp 1677622389
transform 1 0 1340 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7593
timestamp 1677622389
transform 1 0 1340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7594
timestamp 1677622389
transform 1 0 1372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6740
timestamp 1677622389
transform 1 0 1372 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6673
timestamp 1677622389
transform 1 0 1388 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7595
timestamp 1677622389
transform 1 0 1388 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6592
timestamp 1677622389
transform 1 0 1404 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6593
timestamp 1677622389
transform 1 0 1420 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7596
timestamp 1677622389
transform 1 0 1420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7496
timestamp 1677622389
transform 1 0 1436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7497
timestamp 1677622389
transform 1 0 1444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7498
timestamp 1677622389
transform 1 0 1468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7597
timestamp 1677622389
transform 1 0 1452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7598
timestamp 1677622389
transform 1 0 1468 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6741
timestamp 1677622389
transform 1 0 1444 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6742
timestamp 1677622389
transform 1 0 1468 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7599
timestamp 1677622389
transform 1 0 1484 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6769
timestamp 1677622389
transform 1 0 1476 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6594
timestamp 1677622389
transform 1 0 1556 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6595
timestamp 1677622389
transform 1 0 1572 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7499
timestamp 1677622389
transform 1 0 1572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7600
timestamp 1677622389
transform 1 0 1532 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6705
timestamp 1677622389
transform 1 0 1524 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6743
timestamp 1677622389
transform 1 0 1508 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6640
timestamp 1677622389
transform 1 0 1588 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6596
timestamp 1677622389
transform 1 0 1628 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6597
timestamp 1677622389
transform 1 0 1660 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7500
timestamp 1677622389
transform 1 0 1604 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6674
timestamp 1677622389
transform 1 0 1652 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6675
timestamp 1677622389
transform 1 0 1692 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7601
timestamp 1677622389
transform 1 0 1652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7602
timestamp 1677622389
transform 1 0 1684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7603
timestamp 1677622389
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6744
timestamp 1677622389
transform 1 0 1684 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6676
timestamp 1677622389
transform 1 0 1724 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7604
timestamp 1677622389
transform 1 0 1724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7501
timestamp 1677622389
transform 1 0 1748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7502
timestamp 1677622389
transform 1 0 1756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7503
timestamp 1677622389
transform 1 0 1780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7605
timestamp 1677622389
transform 1 0 1764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7606
timestamp 1677622389
transform 1 0 1780 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6706
timestamp 1677622389
transform 1 0 1780 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6745
timestamp 1677622389
transform 1 0 1756 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7504
timestamp 1677622389
transform 1 0 1828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7505
timestamp 1677622389
transform 1 0 1836 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6677
timestamp 1677622389
transform 1 0 1852 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7607
timestamp 1677622389
transform 1 0 1844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7608
timestamp 1677622389
transform 1 0 1852 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6770
timestamp 1677622389
transform 1 0 1852 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6678
timestamp 1677622389
transform 1 0 1948 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7506
timestamp 1677622389
transform 1 0 1972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7609
timestamp 1677622389
transform 1 0 1948 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6707
timestamp 1677622389
transform 1 0 1892 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6641
timestamp 1677622389
transform 1 0 1988 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7507
timestamp 1677622389
transform 1 0 1988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7610
timestamp 1677622389
transform 1 0 2012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7508
timestamp 1677622389
transform 1 0 2044 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6679
timestamp 1677622389
transform 1 0 2060 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7611
timestamp 1677622389
transform 1 0 2036 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7612
timestamp 1677622389
transform 1 0 2052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7613
timestamp 1677622389
transform 1 0 2060 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6708
timestamp 1677622389
transform 1 0 2036 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6746
timestamp 1677622389
transform 1 0 2052 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7509
timestamp 1677622389
transform 1 0 2084 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6709
timestamp 1677622389
transform 1 0 2084 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7614
timestamp 1677622389
transform 1 0 2140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7675
timestamp 1677622389
transform 1 0 2132 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7676
timestamp 1677622389
transform 1 0 2156 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7681
timestamp 1677622389
transform 1 0 2148 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6747
timestamp 1677622389
transform 1 0 2156 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6611
timestamp 1677622389
transform 1 0 2172 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7677
timestamp 1677622389
transform 1 0 2172 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6748
timestamp 1677622389
transform 1 0 2172 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6598
timestamp 1677622389
transform 1 0 2188 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7682
timestamp 1677622389
transform 1 0 2196 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6599
timestamp 1677622389
transform 1 0 2228 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6642
timestamp 1677622389
transform 1 0 2228 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7683
timestamp 1677622389
transform 1 0 2220 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6600
timestamp 1677622389
transform 1 0 2244 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7615
timestamp 1677622389
transform 1 0 2236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7678
timestamp 1677622389
transform 1 0 2276 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6643
timestamp 1677622389
transform 1 0 2364 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7510
timestamp 1677622389
transform 1 0 2364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7616
timestamp 1677622389
transform 1 0 2332 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6710
timestamp 1677622389
transform 1 0 2332 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6644
timestamp 1677622389
transform 1 0 2380 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6711
timestamp 1677622389
transform 1 0 2388 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6612
timestamp 1677622389
transform 1 0 2404 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6645
timestamp 1677622389
transform 1 0 2412 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7511
timestamp 1677622389
transform 1 0 2412 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6771
timestamp 1677622389
transform 1 0 2404 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6601
timestamp 1677622389
transform 1 0 2460 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6613
timestamp 1677622389
transform 1 0 2492 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7477
timestamp 1677622389
transform 1 0 2524 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7617
timestamp 1677622389
transform 1 0 2428 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7618
timestamp 1677622389
transform 1 0 2436 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6712
timestamp 1677622389
transform 1 0 2428 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6646
timestamp 1677622389
transform 1 0 2548 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7512
timestamp 1677622389
transform 1 0 2540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7513
timestamp 1677622389
transform 1 0 2548 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6749
timestamp 1677622389
transform 1 0 2436 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6750
timestamp 1677622389
transform 1 0 2476 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6751
timestamp 1677622389
transform 1 0 2508 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6752
timestamp 1677622389
transform 1 0 2532 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6772
timestamp 1677622389
transform 1 0 2468 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6781
timestamp 1677622389
transform 1 0 2420 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6782
timestamp 1677622389
transform 1 0 2500 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7619
timestamp 1677622389
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7620
timestamp 1677622389
transform 1 0 2572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7621
timestamp 1677622389
transform 1 0 2588 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6602
timestamp 1677622389
transform 1 0 2628 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6603
timestamp 1677622389
transform 1 0 2660 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7514
timestamp 1677622389
transform 1 0 2604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7515
timestamp 1677622389
transform 1 0 2620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7622
timestamp 1677622389
transform 1 0 2612 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6689
timestamp 1677622389
transform 1 0 2620 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7516
timestamp 1677622389
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7623
timestamp 1677622389
transform 1 0 2628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7624
timestamp 1677622389
transform 1 0 2636 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6690
timestamp 1677622389
transform 1 0 2644 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7625
timestamp 1677622389
transform 1 0 2692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6713
timestamp 1677622389
transform 1 0 2636 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6714
timestamp 1677622389
transform 1 0 2692 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6753
timestamp 1677622389
transform 1 0 2620 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6754
timestamp 1677622389
transform 1 0 2652 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6647
timestamp 1677622389
transform 1 0 2732 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7517
timestamp 1677622389
transform 1 0 2732 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7626
timestamp 1677622389
transform 1 0 2732 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6715
timestamp 1677622389
transform 1 0 2732 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6614
timestamp 1677622389
transform 1 0 2852 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6648
timestamp 1677622389
transform 1 0 2780 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7478
timestamp 1677622389
transform 1 0 2852 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6649
timestamp 1677622389
transform 1 0 2860 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7518
timestamp 1677622389
transform 1 0 2860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7519
timestamp 1677622389
transform 1 0 2868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7627
timestamp 1677622389
transform 1 0 2764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7628
timestamp 1677622389
transform 1 0 2876 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6716
timestamp 1677622389
transform 1 0 2876 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6650
timestamp 1677622389
transform 1 0 2892 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7479
timestamp 1677622389
transform 1 0 2996 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7520
timestamp 1677622389
transform 1 0 2892 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6615
timestamp 1677622389
transform 1 0 3012 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7521
timestamp 1677622389
transform 1 0 3004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7522
timestamp 1677622389
transform 1 0 3012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7629
timestamp 1677622389
transform 1 0 2908 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6691
timestamp 1677622389
transform 1 0 2996 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6755
timestamp 1677622389
transform 1 0 2900 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6692
timestamp 1677622389
transform 1 0 3020 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6756
timestamp 1677622389
transform 1 0 3012 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7679
timestamp 1677622389
transform 1 0 3036 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6651
timestamp 1677622389
transform 1 0 3068 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7523
timestamp 1677622389
transform 1 0 3068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7630
timestamp 1677622389
transform 1 0 3084 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6616
timestamp 1677622389
transform 1 0 3108 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7680
timestamp 1677622389
transform 1 0 3100 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7524
timestamp 1677622389
transform 1 0 3108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7631
timestamp 1677622389
transform 1 0 3108 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6757
timestamp 1677622389
transform 1 0 3084 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6758
timestamp 1677622389
transform 1 0 3100 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6773
timestamp 1677622389
transform 1 0 3100 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6693
timestamp 1677622389
transform 1 0 3116 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6617
timestamp 1677622389
transform 1 0 3148 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7480
timestamp 1677622389
transform 1 0 3148 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7525
timestamp 1677622389
transform 1 0 3140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7632
timestamp 1677622389
transform 1 0 3124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7633
timestamp 1677622389
transform 1 0 3132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6717
timestamp 1677622389
transform 1 0 3140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6774
timestamp 1677622389
transform 1 0 3132 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7526
timestamp 1677622389
transform 1 0 3180 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6680
timestamp 1677622389
transform 1 0 3188 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6694
timestamp 1677622389
transform 1 0 3180 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7634
timestamp 1677622389
transform 1 0 3188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7635
timestamp 1677622389
transform 1 0 3196 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6759
timestamp 1677622389
transform 1 0 3196 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6618
timestamp 1677622389
transform 1 0 3260 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7527
timestamp 1677622389
transform 1 0 3236 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6681
timestamp 1677622389
transform 1 0 3244 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7528
timestamp 1677622389
transform 1 0 3260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7636
timestamp 1677622389
transform 1 0 3244 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6718
timestamp 1677622389
transform 1 0 3244 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6619
timestamp 1677622389
transform 1 0 3292 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7529
timestamp 1677622389
transform 1 0 3284 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6760
timestamp 1677622389
transform 1 0 3284 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7637
timestamp 1677622389
transform 1 0 3308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6719
timestamp 1677622389
transform 1 0 3308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6620
timestamp 1677622389
transform 1 0 3332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6652
timestamp 1677622389
transform 1 0 3332 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6653
timestamp 1677622389
transform 1 0 3348 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7530
timestamp 1677622389
transform 1 0 3364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7638
timestamp 1677622389
transform 1 0 3340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7639
timestamp 1677622389
transform 1 0 3356 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6654
timestamp 1677622389
transform 1 0 3396 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7481
timestamp 1677622389
transform 1 0 3404 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6655
timestamp 1677622389
transform 1 0 3452 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7531
timestamp 1677622389
transform 1 0 3396 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7640
timestamp 1677622389
transform 1 0 3388 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6682
timestamp 1677622389
transform 1 0 3500 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7532
timestamp 1677622389
transform 1 0 3508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7641
timestamp 1677622389
transform 1 0 3492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7642
timestamp 1677622389
transform 1 0 3500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6720
timestamp 1677622389
transform 1 0 3500 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7533
timestamp 1677622389
transform 1 0 3524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7534
timestamp 1677622389
transform 1 0 3540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7643
timestamp 1677622389
transform 1 0 3540 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6775
timestamp 1677622389
transform 1 0 3540 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6621
timestamp 1677622389
transform 1 0 3556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6622
timestamp 1677622389
transform 1 0 3588 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6656
timestamp 1677622389
transform 1 0 3580 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7535
timestamp 1677622389
transform 1 0 3580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7536
timestamp 1677622389
transform 1 0 3604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7537
timestamp 1677622389
transform 1 0 3620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7644
timestamp 1677622389
transform 1 0 3588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7645
timestamp 1677622389
transform 1 0 3596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7646
timestamp 1677622389
transform 1 0 3612 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6721
timestamp 1677622389
transform 1 0 3588 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6722
timestamp 1677622389
transform 1 0 3620 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6776
timestamp 1677622389
transform 1 0 3612 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6657
timestamp 1677622389
transform 1 0 3668 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7538
timestamp 1677622389
transform 1 0 3668 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6658
timestamp 1677622389
transform 1 0 3700 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7539
timestamp 1677622389
transform 1 0 3692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7540
timestamp 1677622389
transform 1 0 3708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7647
timestamp 1677622389
transform 1 0 3684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7648
timestamp 1677622389
transform 1 0 3700 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6723
timestamp 1677622389
transform 1 0 3708 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6761
timestamp 1677622389
transform 1 0 3700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6777
timestamp 1677622389
transform 1 0 3684 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6778
timestamp 1677622389
transform 1 0 3708 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6783
timestamp 1677622389
transform 1 0 3684 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6604
timestamp 1677622389
transform 1 0 3724 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7649
timestamp 1677622389
transform 1 0 3732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7541
timestamp 1677622389
transform 1 0 3780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7542
timestamp 1677622389
transform 1 0 3796 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6659
timestamp 1677622389
transform 1 0 3812 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7650
timestamp 1677622389
transform 1 0 3804 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6683
timestamp 1677622389
transform 1 0 3828 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6623
timestamp 1677622389
transform 1 0 3900 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6660
timestamp 1677622389
transform 1 0 3932 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7543
timestamp 1677622389
transform 1 0 3900 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6684
timestamp 1677622389
transform 1 0 3908 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7544
timestamp 1677622389
transform 1 0 3916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7545
timestamp 1677622389
transform 1 0 3932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7651
timestamp 1677622389
transform 1 0 3908 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7652
timestamp 1677622389
transform 1 0 3924 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6695
timestamp 1677622389
transform 1 0 3932 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7653
timestamp 1677622389
transform 1 0 3940 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6724
timestamp 1677622389
transform 1 0 3908 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6685
timestamp 1677622389
transform 1 0 3948 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6725
timestamp 1677622389
transform 1 0 3940 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6686
timestamp 1677622389
transform 1 0 3972 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7654
timestamp 1677622389
transform 1 0 3972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7546
timestamp 1677622389
transform 1 0 4020 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6661
timestamp 1677622389
transform 1 0 4044 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6624
timestamp 1677622389
transform 1 0 4076 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7547
timestamp 1677622389
transform 1 0 4044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7548
timestamp 1677622389
transform 1 0 4060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7549
timestamp 1677622389
transform 1 0 4076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7655
timestamp 1677622389
transform 1 0 4052 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6696
timestamp 1677622389
transform 1 0 4060 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7656
timestamp 1677622389
transform 1 0 4132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6697
timestamp 1677622389
transform 1 0 4140 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7550
timestamp 1677622389
transform 1 0 4164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7551
timestamp 1677622389
transform 1 0 4196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7552
timestamp 1677622389
transform 1 0 4236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7657
timestamp 1677622389
transform 1 0 4228 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6698
timestamp 1677622389
transform 1 0 4236 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7658
timestamp 1677622389
transform 1 0 4244 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6726
timestamp 1677622389
transform 1 0 4228 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7659
timestamp 1677622389
transform 1 0 4260 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6605
timestamp 1677622389
transform 1 0 4284 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6625
timestamp 1677622389
transform 1 0 4284 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7553
timestamp 1677622389
transform 1 0 4284 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6662
timestamp 1677622389
transform 1 0 4300 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7554
timestamp 1677622389
transform 1 0 4300 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6727
timestamp 1677622389
transform 1 0 4300 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6626
timestamp 1677622389
transform 1 0 4332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6663
timestamp 1677622389
transform 1 0 4324 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7555
timestamp 1677622389
transform 1 0 4324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7556
timestamp 1677622389
transform 1 0 4340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7660
timestamp 1677622389
transform 1 0 4316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7661
timestamp 1677622389
transform 1 0 4332 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6728
timestamp 1677622389
transform 1 0 4316 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6762
timestamp 1677622389
transform 1 0 4332 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7662
timestamp 1677622389
transform 1 0 4356 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6729
timestamp 1677622389
transform 1 0 4356 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6606
timestamp 1677622389
transform 1 0 4412 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6627
timestamp 1677622389
transform 1 0 4396 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7557
timestamp 1677622389
transform 1 0 4388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7558
timestamp 1677622389
transform 1 0 4404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7663
timestamp 1677622389
transform 1 0 4396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7664
timestamp 1677622389
transform 1 0 4412 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6763
timestamp 1677622389
transform 1 0 4412 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7665
timestamp 1677622389
transform 1 0 4428 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6664
timestamp 1677622389
transform 1 0 4452 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7559
timestamp 1677622389
transform 1 0 4452 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6687
timestamp 1677622389
transform 1 0 4460 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7560
timestamp 1677622389
transform 1 0 4468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7666
timestamp 1677622389
transform 1 0 4468 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6730
timestamp 1677622389
transform 1 0 4468 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6628
timestamp 1677622389
transform 1 0 4508 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6665
timestamp 1677622389
transform 1 0 4508 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6688
timestamp 1677622389
transform 1 0 4484 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7561
timestamp 1677622389
transform 1 0 4492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7562
timestamp 1677622389
transform 1 0 4508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7667
timestamp 1677622389
transform 1 0 4500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6764
timestamp 1677622389
transform 1 0 4500 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6607
timestamp 1677622389
transform 1 0 4524 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7563
timestamp 1677622389
transform 1 0 4540 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6629
timestamp 1677622389
transform 1 0 4596 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6666
timestamp 1677622389
transform 1 0 4588 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7564
timestamp 1677622389
transform 1 0 4572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7565
timestamp 1677622389
transform 1 0 4588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7668
timestamp 1677622389
transform 1 0 4564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7669
timestamp 1677622389
transform 1 0 4580 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6731
timestamp 1677622389
transform 1 0 4580 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7670
timestamp 1677622389
transform 1 0 4596 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6765
timestamp 1677622389
transform 1 0 4564 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6766
timestamp 1677622389
transform 1 0 4588 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7566
timestamp 1677622389
transform 1 0 4628 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6732
timestamp 1677622389
transform 1 0 4628 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6608
timestamp 1677622389
transform 1 0 4660 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6609
timestamp 1677622389
transform 1 0 4684 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7567
timestamp 1677622389
transform 1 0 4652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7568
timestamp 1677622389
transform 1 0 4668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7569
timestamp 1677622389
transform 1 0 4676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7671
timestamp 1677622389
transform 1 0 4660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7672
timestamp 1677622389
transform 1 0 4676 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6630
timestamp 1677622389
transform 1 0 4708 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6631
timestamp 1677622389
transform 1 0 4732 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6667
timestamp 1677622389
transform 1 0 4724 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7570
timestamp 1677622389
transform 1 0 4700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7571
timestamp 1677622389
transform 1 0 4716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7673
timestamp 1677622389
transform 1 0 4708 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6733
timestamp 1677622389
transform 1 0 4676 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6734
timestamp 1677622389
transform 1 0 4692 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6735
timestamp 1677622389
transform 1 0 4708 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7674
timestamp 1677622389
transform 1 0 4724 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6632
timestamp 1677622389
transform 1 0 4756 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7572
timestamp 1677622389
transform 1 0 4780 0 1 1135
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_72
timestamp 1677622389
transform 1 0 24 0 1 1070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_461
timestamp 1677622389
transform 1 0 72 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8472
timestamp 1677622389
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8473
timestamp 1677622389
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8474
timestamp 1677622389
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_462
timestamp 1677622389
transform 1 0 192 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8475
timestamp 1677622389
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8476
timestamp 1677622389
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8477
timestamp 1677622389
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8478
timestamp 1677622389
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8480
timestamp 1677622389
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8482
timestamp 1677622389
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8484
timestamp 1677622389
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8501
timestamp 1677622389
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8502
timestamp 1677622389
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_464
timestamp 1677622389
transform -1 0 456 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8503
timestamp 1677622389
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8504
timestamp 1677622389
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_465
timestamp 1677622389
transform 1 0 472 0 -1 1170
box -8 -3 104 105
use AOI22X1  AOI22X1_313
timestamp 1677622389
transform 1 0 568 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8505
timestamp 1677622389
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8506
timestamp 1677622389
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_537
timestamp 1677622389
transform -1 0 640 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8507
timestamp 1677622389
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8508
timestamp 1677622389
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_466
timestamp 1677622389
transform -1 0 752 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8509
timestamp 1677622389
transform 1 0 752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8517
timestamp 1677622389
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_467
timestamp 1677622389
transform -1 0 864 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8518
timestamp 1677622389
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8521
timestamp 1677622389
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_539
timestamp 1677622389
transform -1 0 896 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8522
timestamp 1677622389
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8523
timestamp 1677622389
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8524
timestamp 1677622389
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8525
timestamp 1677622389
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_86
timestamp 1677622389
transform 1 0 928 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8530
timestamp 1677622389
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8531
timestamp 1677622389
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8532
timestamp 1677622389
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8533
timestamp 1677622389
transform 1 0 976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8535
timestamp 1677622389
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8537
timestamp 1677622389
transform 1 0 992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8538
timestamp 1677622389
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8539
timestamp 1677622389
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8540
timestamp 1677622389
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8541
timestamp 1677622389
transform 1 0 1024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8542
timestamp 1677622389
transform 1 0 1032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8543
timestamp 1677622389
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8544
timestamp 1677622389
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_88
timestamp 1677622389
transform 1 0 1056 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8545
timestamp 1677622389
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8546
timestamp 1677622389
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8547
timestamp 1677622389
transform 1 0 1096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8548
timestamp 1677622389
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8549
timestamp 1677622389
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8551
timestamp 1677622389
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8556
timestamp 1677622389
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_540
timestamp 1677622389
transform -1 0 1152 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8557
timestamp 1677622389
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8559
timestamp 1677622389
transform 1 0 1160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8561
timestamp 1677622389
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8563
timestamp 1677622389
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8565
timestamp 1677622389
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8568
timestamp 1677622389
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8569
timestamp 1677622389
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8570
timestamp 1677622389
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8571
timestamp 1677622389
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8572
timestamp 1677622389
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8573
timestamp 1677622389
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8574
timestamp 1677622389
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8576
timestamp 1677622389
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8578
timestamp 1677622389
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8580
timestamp 1677622389
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8582
timestamp 1677622389
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_469
timestamp 1677622389
transform 1 0 1280 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8591
timestamp 1677622389
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8598
timestamp 1677622389
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_542
timestamp 1677622389
transform -1 0 1408 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8599
timestamp 1677622389
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8600
timestamp 1677622389
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8601
timestamp 1677622389
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_318
timestamp 1677622389
transform -1 0 1472 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8602
timestamp 1677622389
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8603
timestamp 1677622389
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_472
timestamp 1677622389
transform -1 0 1584 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8604
timestamp 1677622389
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_473
timestamp 1677622389
transform 1 0 1592 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8605
timestamp 1677622389
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8606
timestamp 1677622389
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8621
timestamp 1677622389
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_543
timestamp 1677622389
transform -1 0 1728 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8622
timestamp 1677622389
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8623
timestamp 1677622389
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_320
timestamp 1677622389
transform -1 0 1784 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8624
timestamp 1677622389
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8625
timestamp 1677622389
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8626
timestamp 1677622389
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8627
timestamp 1677622389
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8628
timestamp 1677622389
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8629
timestamp 1677622389
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_544
timestamp 1677622389
transform 1 0 1832 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8630
timestamp 1677622389
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8631
timestamp 1677622389
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8632
timestamp 1677622389
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8633
timestamp 1677622389
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8634
timestamp 1677622389
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_475
timestamp 1677622389
transform -1 0 1984 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8635
timestamp 1677622389
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8637
timestamp 1677622389
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8639
timestamp 1677622389
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8645
timestamp 1677622389
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_321
timestamp 1677622389
transform -1 0 2056 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8646
timestamp 1677622389
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8651
timestamp 1677622389
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_546
timestamp 1677622389
transform -1 0 2088 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8652
timestamp 1677622389
transform 1 0 2088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8654
timestamp 1677622389
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8660
timestamp 1677622389
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8661
timestamp 1677622389
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8662
timestamp 1677622389
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_65
timestamp 1677622389
transform 1 0 2128 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8663
timestamp 1677622389
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8664
timestamp 1677622389
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8665
timestamp 1677622389
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8666
timestamp 1677622389
transform 1 0 2184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8668
timestamp 1677622389
transform 1 0 2192 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_66
timestamp 1677622389
transform 1 0 2200 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8677
timestamp 1677622389
transform 1 0 2232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8678
timestamp 1677622389
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8679
timestamp 1677622389
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8680
timestamp 1677622389
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8681
timestamp 1677622389
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8682
timestamp 1677622389
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_477
timestamp 1677622389
transform -1 0 2376 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8683
timestamp 1677622389
transform 1 0 2376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8684
timestamp 1677622389
transform 1 0 2384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8685
timestamp 1677622389
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8686
timestamp 1677622389
transform 1 0 2400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8687
timestamp 1677622389
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_9
timestamp 1677622389
transform 1 0 2416 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8703
timestamp 1677622389
transform 1 0 2536 0 -1 1170
box -8 -3 16 105
use AND2X2  AND2X2_52
timestamp 1677622389
transform 1 0 2544 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8704
timestamp 1677622389
transform 1 0 2576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8706
timestamp 1677622389
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_322
timestamp 1677622389
transform 1 0 2592 0 -1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_479
timestamp 1677622389
transform -1 0 2728 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8710
timestamp 1677622389
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8711
timestamp 1677622389
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_11
timestamp 1677622389
transform 1 0 2744 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8712
timestamp 1677622389
transform 1 0 2864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8713
timestamp 1677622389
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8714
timestamp 1677622389
transform 1 0 2880 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_13
timestamp 1677622389
transform 1 0 2888 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8716
timestamp 1677622389
transform 1 0 3008 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_18
timestamp 1677622389
transform 1 0 3016 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8718
timestamp 1677622389
transform 1 0 3040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8720
timestamp 1677622389
transform 1 0 3048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8722
timestamp 1677622389
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8724
timestamp 1677622389
transform 1 0 3064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8730
timestamp 1677622389
transform 1 0 3072 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_549
timestamp 1677622389
transform 1 0 3080 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8731
timestamp 1677622389
transform 1 0 3096 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_150
timestamp 1677622389
transform -1 0 3136 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8732
timestamp 1677622389
transform 1 0 3136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8736
timestamp 1677622389
transform 1 0 3144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8737
timestamp 1677622389
transform 1 0 3152 0 -1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_11
timestamp 1677622389
transform -1 0 3192 0 -1 1170
box -7 -3 39 105
use FILL  FILL_8738
timestamp 1677622389
transform 1 0 3192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8739
timestamp 1677622389
transform 1 0 3200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8740
timestamp 1677622389
transform 1 0 3208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8743
timestamp 1677622389
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_324
timestamp 1677622389
transform -1 0 3264 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8744
timestamp 1677622389
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8745
timestamp 1677622389
transform 1 0 3272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8746
timestamp 1677622389
transform 1 0 3280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8748
timestamp 1677622389
transform 1 0 3288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8750
timestamp 1677622389
transform 1 0 3296 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_552
timestamp 1677622389
transform 1 0 3304 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8755
timestamp 1677622389
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8756
timestamp 1677622389
transform 1 0 3328 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_325
timestamp 1677622389
transform 1 0 3336 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8757
timestamp 1677622389
transform 1 0 3376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8758
timestamp 1677622389
transform 1 0 3384 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_15
timestamp 1677622389
transform -1 0 3512 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8759
timestamp 1677622389
transform 1 0 3512 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_553
timestamp 1677622389
transform 1 0 3520 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_554
timestamp 1677622389
transform 1 0 3536 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8760
timestamp 1677622389
transform 1 0 3552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8761
timestamp 1677622389
transform 1 0 3560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8762
timestamp 1677622389
transform 1 0 3568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8763
timestamp 1677622389
transform 1 0 3576 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_323
timestamp 1677622389
transform 1 0 3584 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8767
timestamp 1677622389
transform 1 0 3624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8768
timestamp 1677622389
transform 1 0 3632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8769
timestamp 1677622389
transform 1 0 3640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8771
timestamp 1677622389
transform 1 0 3648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8773
timestamp 1677622389
transform 1 0 3656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8775
timestamp 1677622389
transform 1 0 3664 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_324
timestamp 1677622389
transform 1 0 3672 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8778
timestamp 1677622389
transform 1 0 3712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8779
timestamp 1677622389
transform 1 0 3720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8780
timestamp 1677622389
transform 1 0 3728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8781
timestamp 1677622389
transform 1 0 3736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8782
timestamp 1677622389
transform 1 0 3744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8783
timestamp 1677622389
transform 1 0 3752 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_555
timestamp 1677622389
transform -1 0 3776 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8784
timestamp 1677622389
transform 1 0 3776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8786
timestamp 1677622389
transform 1 0 3784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8788
timestamp 1677622389
transform 1 0 3792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8790
timestamp 1677622389
transform 1 0 3800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8792
timestamp 1677622389
transform 1 0 3808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8793
timestamp 1677622389
transform 1 0 3816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8794
timestamp 1677622389
transform 1 0 3824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8795
timestamp 1677622389
transform 1 0 3832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8796
timestamp 1677622389
transform 1 0 3840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8797
timestamp 1677622389
transform 1 0 3848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8799
timestamp 1677622389
transform 1 0 3856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8801
timestamp 1677622389
transform 1 0 3864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8802
timestamp 1677622389
transform 1 0 3872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8803
timestamp 1677622389
transform 1 0 3880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8804
timestamp 1677622389
transform 1 0 3888 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_326
timestamp 1677622389
transform 1 0 3896 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8810
timestamp 1677622389
transform 1 0 3936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8811
timestamp 1677622389
transform 1 0 3944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8812
timestamp 1677622389
transform 1 0 3952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8813
timestamp 1677622389
transform 1 0 3960 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_556
timestamp 1677622389
transform -1 0 3984 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8814
timestamp 1677622389
transform 1 0 3984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8815
timestamp 1677622389
transform 1 0 3992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8816
timestamp 1677622389
transform 1 0 4000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8817
timestamp 1677622389
transform 1 0 4008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8818
timestamp 1677622389
transform 1 0 4016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8819
timestamp 1677622389
transform 1 0 4024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8824
timestamp 1677622389
transform 1 0 4032 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_327
timestamp 1677622389
transform -1 0 4080 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8825
timestamp 1677622389
transform 1 0 4080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8826
timestamp 1677622389
transform 1 0 4088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8827
timestamp 1677622389
transform 1 0 4096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8828
timestamp 1677622389
transform 1 0 4104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8829
timestamp 1677622389
transform 1 0 4112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8830
timestamp 1677622389
transform 1 0 4120 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_558
timestamp 1677622389
transform -1 0 4144 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8831
timestamp 1677622389
transform 1 0 4144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8832
timestamp 1677622389
transform 1 0 4152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8833
timestamp 1677622389
transform 1 0 4160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8834
timestamp 1677622389
transform 1 0 4168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8836
timestamp 1677622389
transform 1 0 4176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8838
timestamp 1677622389
transform 1 0 4184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8839
timestamp 1677622389
transform 1 0 4192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8840
timestamp 1677622389
transform 1 0 4200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8841
timestamp 1677622389
transform 1 0 4208 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6784
timestamp 1677622389
transform 1 0 4236 0 1 1075
box -3 -3 3 3
use OAI22X1  OAI22X1_328
timestamp 1677622389
transform 1 0 4216 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8842
timestamp 1677622389
transform 1 0 4256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8843
timestamp 1677622389
transform 1 0 4264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8844
timestamp 1677622389
transform 1 0 4272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8845
timestamp 1677622389
transform 1 0 4280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8847
timestamp 1677622389
transform 1 0 4288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8853
timestamp 1677622389
transform 1 0 4296 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_329
timestamp 1677622389
transform 1 0 4304 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8854
timestamp 1677622389
transform 1 0 4344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8860
timestamp 1677622389
transform 1 0 4352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8861
timestamp 1677622389
transform 1 0 4360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8862
timestamp 1677622389
transform 1 0 4368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8863
timestamp 1677622389
transform 1 0 4376 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6785
timestamp 1677622389
transform 1 0 4428 0 1 1075
box -3 -3 3 3
use OAI22X1  OAI22X1_331
timestamp 1677622389
transform 1 0 4384 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8864
timestamp 1677622389
transform 1 0 4424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8866
timestamp 1677622389
transform 1 0 4432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8869
timestamp 1677622389
transform 1 0 4440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8870
timestamp 1677622389
transform 1 0 4448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8871
timestamp 1677622389
transform 1 0 4456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8872
timestamp 1677622389
transform 1 0 4464 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_333
timestamp 1677622389
transform 1 0 4472 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8877
timestamp 1677622389
transform 1 0 4512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8878
timestamp 1677622389
transform 1 0 4520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8879
timestamp 1677622389
transform 1 0 4528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8880
timestamp 1677622389
transform 1 0 4536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8884
timestamp 1677622389
transform 1 0 4544 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_334
timestamp 1677622389
transform -1 0 4592 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8885
timestamp 1677622389
transform 1 0 4592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8887
timestamp 1677622389
transform 1 0 4600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8889
timestamp 1677622389
transform 1 0 4608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8893
timestamp 1677622389
transform 1 0 4616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8894
timestamp 1677622389
transform 1 0 4624 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_336
timestamp 1677622389
transform 1 0 4632 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8895
timestamp 1677622389
transform 1 0 4672 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_337
timestamp 1677622389
transform 1 0 4680 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8898
timestamp 1677622389
transform 1 0 4720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8899
timestamp 1677622389
transform 1 0 4728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8900
timestamp 1677622389
transform 1 0 4736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8901
timestamp 1677622389
transform 1 0 4744 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_561
timestamp 1677622389
transform -1 0 4768 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8902
timestamp 1677622389
transform 1 0 4768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8903
timestamp 1677622389
transform 1 0 4776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8904
timestamp 1677622389
transform 1 0 4784 0 -1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_73
timestamp 1677622389
transform 1 0 4843 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_6813
timestamp 1677622389
transform 1 0 92 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6842
timestamp 1677622389
transform 1 0 76 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7699
timestamp 1677622389
transform 1 0 84 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7700
timestamp 1677622389
transform 1 0 92 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7701
timestamp 1677622389
transform 1 0 108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7806
timestamp 1677622389
transform 1 0 76 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7807
timestamp 1677622389
transform 1 0 100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7808
timestamp 1677622389
transform 1 0 132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6914
timestamp 1677622389
transform 1 0 132 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6814
timestamp 1677622389
transform 1 0 156 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7702
timestamp 1677622389
transform 1 0 148 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6895
timestamp 1677622389
transform 1 0 148 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7703
timestamp 1677622389
transform 1 0 156 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6815
timestamp 1677622389
transform 1 0 180 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6843
timestamp 1677622389
transform 1 0 180 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6873
timestamp 1677622389
transform 1 0 172 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7704
timestamp 1677622389
transform 1 0 180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7809
timestamp 1677622389
transform 1 0 172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7810
timestamp 1677622389
transform 1 0 188 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6915
timestamp 1677622389
transform 1 0 188 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6844
timestamp 1677622389
transform 1 0 228 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7705
timestamp 1677622389
transform 1 0 228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7706
timestamp 1677622389
transform 1 0 236 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6845
timestamp 1677622389
transform 1 0 252 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7707
timestamp 1677622389
transform 1 0 252 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6792
timestamp 1677622389
transform 1 0 284 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6846
timestamp 1677622389
transform 1 0 292 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7708
timestamp 1677622389
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7709
timestamp 1677622389
transform 1 0 300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7710
timestamp 1677622389
transform 1 0 316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7811
timestamp 1677622389
transform 1 0 284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7812
timestamp 1677622389
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7813
timestamp 1677622389
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6847
timestamp 1677622389
transform 1 0 332 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6896
timestamp 1677622389
transform 1 0 340 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7711
timestamp 1677622389
transform 1 0 356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7712
timestamp 1677622389
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6874
timestamp 1677622389
transform 1 0 380 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7814
timestamp 1677622389
transform 1 0 364 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6897
timestamp 1677622389
transform 1 0 372 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7815
timestamp 1677622389
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6916
timestamp 1677622389
transform 1 0 364 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6940
timestamp 1677622389
transform 1 0 356 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6875
timestamp 1677622389
transform 1 0 404 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7713
timestamp 1677622389
transform 1 0 444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7714
timestamp 1677622389
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7816
timestamp 1677622389
transform 1 0 404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6793
timestamp 1677622389
transform 1 0 572 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6876
timestamp 1677622389
transform 1 0 516 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7715
timestamp 1677622389
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7716
timestamp 1677622389
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7817
timestamp 1677622389
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7717
timestamp 1677622389
transform 1 0 612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7818
timestamp 1677622389
transform 1 0 628 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6941
timestamp 1677622389
transform 1 0 628 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7718
timestamp 1677622389
transform 1 0 652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7819
timestamp 1677622389
transform 1 0 644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7719
timestamp 1677622389
transform 1 0 692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7820
timestamp 1677622389
transform 1 0 684 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6786
timestamp 1677622389
transform 1 0 812 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6848
timestamp 1677622389
transform 1 0 804 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7720
timestamp 1677622389
transform 1 0 748 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6877
timestamp 1677622389
transform 1 0 756 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7721
timestamp 1677622389
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7821
timestamp 1677622389
transform 1 0 828 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6942
timestamp 1677622389
transform 1 0 780 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6943
timestamp 1677622389
transform 1 0 796 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6849
timestamp 1677622389
transform 1 0 844 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7722
timestamp 1677622389
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7723
timestamp 1677622389
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6850
timestamp 1677622389
transform 1 0 884 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7822
timestamp 1677622389
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6794
timestamp 1677622389
transform 1 0 924 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6851
timestamp 1677622389
transform 1 0 908 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6852
timestamp 1677622389
transform 1 0 924 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6878
timestamp 1677622389
transform 1 0 900 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7724
timestamp 1677622389
transform 1 0 908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7725
timestamp 1677622389
transform 1 0 924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7823
timestamp 1677622389
transform 1 0 900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7824
timestamp 1677622389
transform 1 0 916 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6917
timestamp 1677622389
transform 1 0 924 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7908
timestamp 1677622389
transform 1 0 932 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_6898
timestamp 1677622389
transform 1 0 948 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7825
timestamp 1677622389
transform 1 0 988 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7909
timestamp 1677622389
transform 1 0 1012 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_6944
timestamp 1677622389
transform 1 0 1012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6787
timestamp 1677622389
transform 1 0 1060 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6795
timestamp 1677622389
transform 1 0 1076 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6853
timestamp 1677622389
transform 1 0 1076 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6945
timestamp 1677622389
transform 1 0 1076 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6854
timestamp 1677622389
transform 1 0 1124 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7726
timestamp 1677622389
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7826
timestamp 1677622389
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7827
timestamp 1677622389
transform 1 0 1156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7727
timestamp 1677622389
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6918
timestamp 1677622389
transform 1 0 1196 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7728
timestamp 1677622389
transform 1 0 1212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7729
timestamp 1677622389
transform 1 0 1236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7828
timestamp 1677622389
transform 1 0 1220 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6919
timestamp 1677622389
transform 1 0 1228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6879
timestamp 1677622389
transform 1 0 1252 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7829
timestamp 1677622389
transform 1 0 1252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7730
timestamp 1677622389
transform 1 0 1332 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6816
timestamp 1677622389
transform 1 0 1420 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7731
timestamp 1677622389
transform 1 0 1420 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6880
timestamp 1677622389
transform 1 0 1428 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7732
timestamp 1677622389
transform 1 0 1436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7830
timestamp 1677622389
transform 1 0 1420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7831
timestamp 1677622389
transform 1 0 1428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7832
timestamp 1677622389
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6946
timestamp 1677622389
transform 1 0 1444 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6817
timestamp 1677622389
transform 1 0 1476 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7733
timestamp 1677622389
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7833
timestamp 1677622389
transform 1 0 1492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7734
timestamp 1677622389
transform 1 0 1508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7735
timestamp 1677622389
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7834
timestamp 1677622389
transform 1 0 1572 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6920
timestamp 1677622389
transform 1 0 1572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6818
timestamp 1677622389
transform 1 0 1596 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7736
timestamp 1677622389
transform 1 0 1588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7737
timestamp 1677622389
transform 1 0 1596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6796
timestamp 1677622389
transform 1 0 1628 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6819
timestamp 1677622389
transform 1 0 1652 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7738
timestamp 1677622389
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6881
timestamp 1677622389
transform 1 0 1644 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7835
timestamp 1677622389
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7836
timestamp 1677622389
transform 1 0 1628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7837
timestamp 1677622389
transform 1 0 1644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7838
timestamp 1677622389
transform 1 0 1652 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6820
timestamp 1677622389
transform 1 0 1676 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7739
timestamp 1677622389
transform 1 0 1668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7740
timestamp 1677622389
transform 1 0 1676 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6921
timestamp 1677622389
transform 1 0 1692 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6821
timestamp 1677622389
transform 1 0 1724 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6855
timestamp 1677622389
transform 1 0 1748 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7741
timestamp 1677622389
transform 1 0 1732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7742
timestamp 1677622389
transform 1 0 1756 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6882
timestamp 1677622389
transform 1 0 1764 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7839
timestamp 1677622389
transform 1 0 1732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6899
timestamp 1677622389
transform 1 0 1740 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7840
timestamp 1677622389
transform 1 0 1748 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6947
timestamp 1677622389
transform 1 0 1748 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6948
timestamp 1677622389
transform 1 0 1772 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7743
timestamp 1677622389
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7841
timestamp 1677622389
transform 1 0 1788 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6822
timestamp 1677622389
transform 1 0 1804 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7744
timestamp 1677622389
transform 1 0 1804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7745
timestamp 1677622389
transform 1 0 1836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7746
timestamp 1677622389
transform 1 0 1852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7747
timestamp 1677622389
transform 1 0 1860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7842
timestamp 1677622389
transform 1 0 1844 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6900
timestamp 1677622389
transform 1 0 1860 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6922
timestamp 1677622389
transform 1 0 1860 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6856
timestamp 1677622389
transform 1 0 1940 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7748
timestamp 1677622389
transform 1 0 1940 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7843
timestamp 1677622389
transform 1 0 1964 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6923
timestamp 1677622389
transform 1 0 1884 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6857
timestamp 1677622389
transform 1 0 1980 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7749
timestamp 1677622389
transform 1 0 1980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7750
timestamp 1677622389
transform 1 0 2012 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6803
timestamp 1677622389
transform 1 0 2052 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6883
timestamp 1677622389
transform 1 0 2028 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6823
timestamp 1677622389
transform 1 0 2060 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7751
timestamp 1677622389
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7752
timestamp 1677622389
transform 1 0 2052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7753
timestamp 1677622389
transform 1 0 2060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7844
timestamp 1677622389
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7845
timestamp 1677622389
transform 1 0 2028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7846
timestamp 1677622389
transform 1 0 2044 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6949
timestamp 1677622389
transform 1 0 2052 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7847
timestamp 1677622389
transform 1 0 2068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7848
timestamp 1677622389
transform 1 0 2092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7754
timestamp 1677622389
transform 1 0 2116 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6858
timestamp 1677622389
transform 1 0 2132 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6804
timestamp 1677622389
transform 1 0 2148 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7755
timestamp 1677622389
transform 1 0 2140 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6859
timestamp 1677622389
transform 1 0 2196 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7756
timestamp 1677622389
transform 1 0 2196 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6884
timestamp 1677622389
transform 1 0 2220 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7849
timestamp 1677622389
transform 1 0 2220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7850
timestamp 1677622389
transform 1 0 2252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7851
timestamp 1677622389
transform 1 0 2260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7852
timestamp 1677622389
transform 1 0 2276 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6824
timestamp 1677622389
transform 1 0 2316 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7685
timestamp 1677622389
transform 1 0 2316 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7757
timestamp 1677622389
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7853
timestamp 1677622389
transform 1 0 2316 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6825
timestamp 1677622389
transform 1 0 2356 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6860
timestamp 1677622389
transform 1 0 2348 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7686
timestamp 1677622389
transform 1 0 2356 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7758
timestamp 1677622389
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6861
timestamp 1677622389
transform 1 0 2404 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6885
timestamp 1677622389
transform 1 0 2380 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7759
timestamp 1677622389
transform 1 0 2404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7854
timestamp 1677622389
transform 1 0 2364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7804
timestamp 1677622389
transform 1 0 2380 0 1 1007
box -2 -2 2 2
use M2_M1  M2_M1_7855
timestamp 1677622389
transform 1 0 2388 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6826
timestamp 1677622389
transform 1 0 2452 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7856
timestamp 1677622389
transform 1 0 2452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7857
timestamp 1677622389
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7760
timestamp 1677622389
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6901
timestamp 1677622389
transform 1 0 2508 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7761
timestamp 1677622389
transform 1 0 2524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7762
timestamp 1677622389
transform 1 0 2548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7858
timestamp 1677622389
transform 1 0 2516 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6950
timestamp 1677622389
transform 1 0 2516 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6886
timestamp 1677622389
transform 1 0 2604 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6902
timestamp 1677622389
transform 1 0 2596 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7859
timestamp 1677622389
transform 1 0 2604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7860
timestamp 1677622389
transform 1 0 2612 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6951
timestamp 1677622389
transform 1 0 2588 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7763
timestamp 1677622389
transform 1 0 2636 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6903
timestamp 1677622389
transform 1 0 2636 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7861
timestamp 1677622389
transform 1 0 2644 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6827
timestamp 1677622389
transform 1 0 2684 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6862
timestamp 1677622389
transform 1 0 2676 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6863
timestamp 1677622389
transform 1 0 2692 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7764
timestamp 1677622389
transform 1 0 2676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7765
timestamp 1677622389
transform 1 0 2684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7766
timestamp 1677622389
transform 1 0 2692 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6904
timestamp 1677622389
transform 1 0 2676 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7862
timestamp 1677622389
transform 1 0 2692 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6788
timestamp 1677622389
transform 1 0 2764 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6828
timestamp 1677622389
transform 1 0 2772 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7767
timestamp 1677622389
transform 1 0 2772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7863
timestamp 1677622389
transform 1 0 2796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7768
timestamp 1677622389
transform 1 0 2820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7864
timestamp 1677622389
transform 1 0 2812 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6952
timestamp 1677622389
transform 1 0 2812 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6789
timestamp 1677622389
transform 1 0 2940 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6829
timestamp 1677622389
transform 1 0 2868 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6830
timestamp 1677622389
transform 1 0 2916 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7769
timestamp 1677622389
transform 1 0 2844 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6887
timestamp 1677622389
transform 1 0 2876 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7865
timestamp 1677622389
transform 1 0 2940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7866
timestamp 1677622389
transform 1 0 2948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7910
timestamp 1677622389
transform 1 0 2932 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_6797
timestamp 1677622389
transform 1 0 3044 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6831
timestamp 1677622389
transform 1 0 3044 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7687
timestamp 1677622389
transform 1 0 3036 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7867
timestamp 1677622389
transform 1 0 3028 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6924
timestamp 1677622389
transform 1 0 3028 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7770
timestamp 1677622389
transform 1 0 3044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7688
timestamp 1677622389
transform 1 0 3060 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6925
timestamp 1677622389
transform 1 0 3052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6798
timestamp 1677622389
transform 1 0 3076 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6805
timestamp 1677622389
transform 1 0 3084 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7684
timestamp 1677622389
transform 1 0 3100 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_7689
timestamp 1677622389
transform 1 0 3084 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6832
timestamp 1677622389
transform 1 0 3116 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7690
timestamp 1677622389
transform 1 0 3108 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7691
timestamp 1677622389
transform 1 0 3116 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7868
timestamp 1677622389
transform 1 0 3156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7771
timestamp 1677622389
transform 1 0 3180 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6864
timestamp 1677622389
transform 1 0 3196 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7869
timestamp 1677622389
transform 1 0 3196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7870
timestamp 1677622389
transform 1 0 3220 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6926
timestamp 1677622389
transform 1 0 3220 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7871
timestamp 1677622389
transform 1 0 3236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7772
timestamp 1677622389
transform 1 0 3252 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6865
timestamp 1677622389
transform 1 0 3284 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7773
timestamp 1677622389
transform 1 0 3284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7872
timestamp 1677622389
transform 1 0 3292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7873
timestamp 1677622389
transform 1 0 3300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6927
timestamp 1677622389
transform 1 0 3300 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6806
timestamp 1677622389
transform 1 0 3356 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7774
timestamp 1677622389
transform 1 0 3404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7775
timestamp 1677622389
transform 1 0 3412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7874
timestamp 1677622389
transform 1 0 3396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6905
timestamp 1677622389
transform 1 0 3404 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7875
timestamp 1677622389
transform 1 0 3508 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6928
timestamp 1677622389
transform 1 0 3476 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7911
timestamp 1677622389
transform 1 0 3500 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7776
timestamp 1677622389
transform 1 0 3524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7777
timestamp 1677622389
transform 1 0 3540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7876
timestamp 1677622389
transform 1 0 3548 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6929
timestamp 1677622389
transform 1 0 3532 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6930
timestamp 1677622389
transform 1 0 3548 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7778
timestamp 1677622389
transform 1 0 3596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6906
timestamp 1677622389
transform 1 0 3620 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6953
timestamp 1677622389
transform 1 0 3644 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6807
timestamp 1677622389
transform 1 0 3684 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6866
timestamp 1677622389
transform 1 0 3668 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7779
timestamp 1677622389
transform 1 0 3668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7780
timestamp 1677622389
transform 1 0 3684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7877
timestamp 1677622389
transform 1 0 3660 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7878
timestamp 1677622389
transform 1 0 3676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6931
timestamp 1677622389
transform 1 0 3660 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7781
timestamp 1677622389
transform 1 0 3708 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6932
timestamp 1677622389
transform 1 0 3716 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6888
timestamp 1677622389
transform 1 0 3732 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7879
timestamp 1677622389
transform 1 0 3732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7880
timestamp 1677622389
transform 1 0 3740 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6933
timestamp 1677622389
transform 1 0 3740 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6799
timestamp 1677622389
transform 1 0 3812 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6833
timestamp 1677622389
transform 1 0 3796 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7782
timestamp 1677622389
transform 1 0 3796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7783
timestamp 1677622389
transform 1 0 3812 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6889
timestamp 1677622389
transform 1 0 3820 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7784
timestamp 1677622389
transform 1 0 3828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7881
timestamp 1677622389
transform 1 0 3804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7882
timestamp 1677622389
transform 1 0 3820 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7692
timestamp 1677622389
transform 1 0 3836 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6890
timestamp 1677622389
transform 1 0 3900 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6800
timestamp 1677622389
transform 1 0 3916 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6834
timestamp 1677622389
transform 1 0 3932 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7785
timestamp 1677622389
transform 1 0 3916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7786
timestamp 1677622389
transform 1 0 3932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7883
timestamp 1677622389
transform 1 0 3900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7884
timestamp 1677622389
transform 1 0 3908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7885
timestamp 1677622389
transform 1 0 3924 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7886
timestamp 1677622389
transform 1 0 3964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7887
timestamp 1677622389
transform 1 0 3972 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6934
timestamp 1677622389
transform 1 0 3964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6808
timestamp 1677622389
transform 1 0 3996 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6867
timestamp 1677622389
transform 1 0 4012 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7787
timestamp 1677622389
transform 1 0 3996 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7788
timestamp 1677622389
transform 1 0 4012 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6835
timestamp 1677622389
transform 1 0 4028 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7789
timestamp 1677622389
transform 1 0 4028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7888
timestamp 1677622389
transform 1 0 4004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7889
timestamp 1677622389
transform 1 0 4020 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6935
timestamp 1677622389
transform 1 0 4020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6790
timestamp 1677622389
transform 1 0 4092 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6801
timestamp 1677622389
transform 1 0 4084 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7790
timestamp 1677622389
transform 1 0 4092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7890
timestamp 1677622389
transform 1 0 4068 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6936
timestamp 1677622389
transform 1 0 4060 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6907
timestamp 1677622389
transform 1 0 4076 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7891
timestamp 1677622389
transform 1 0 4084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7892
timestamp 1677622389
transform 1 0 4132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6809
timestamp 1677622389
transform 1 0 4156 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6810
timestamp 1677622389
transform 1 0 4172 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6868
timestamp 1677622389
transform 1 0 4172 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7791
timestamp 1677622389
transform 1 0 4156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7792
timestamp 1677622389
transform 1 0 4172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7893
timestamp 1677622389
transform 1 0 4164 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6908
timestamp 1677622389
transform 1 0 4172 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7894
timestamp 1677622389
transform 1 0 4180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6802
timestamp 1677622389
transform 1 0 4212 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6811
timestamp 1677622389
transform 1 0 4252 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6836
timestamp 1677622389
transform 1 0 4260 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6869
timestamp 1677622389
transform 1 0 4236 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6870
timestamp 1677622389
transform 1 0 4260 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7793
timestamp 1677622389
transform 1 0 4228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7794
timestamp 1677622389
transform 1 0 4236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7795
timestamp 1677622389
transform 1 0 4252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7895
timestamp 1677622389
transform 1 0 4244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7896
timestamp 1677622389
transform 1 0 4260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7897
timestamp 1677622389
transform 1 0 4268 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6937
timestamp 1677622389
transform 1 0 4268 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7693
timestamp 1677622389
transform 1 0 4308 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6791
timestamp 1677622389
transform 1 0 4332 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6871
timestamp 1677622389
transform 1 0 4340 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6837
timestamp 1677622389
transform 1 0 4372 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7694
timestamp 1677622389
transform 1 0 4372 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6909
timestamp 1677622389
transform 1 0 4372 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7796
timestamp 1677622389
transform 1 0 4404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7898
timestamp 1677622389
transform 1 0 4404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6838
timestamp 1677622389
transform 1 0 4412 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7695
timestamp 1677622389
transform 1 0 4412 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6891
timestamp 1677622389
transform 1 0 4412 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7899
timestamp 1677622389
transform 1 0 4412 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6910
timestamp 1677622389
transform 1 0 4420 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7696
timestamp 1677622389
transform 1 0 4444 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7900
timestamp 1677622389
transform 1 0 4444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7901
timestamp 1677622389
transform 1 0 4452 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6954
timestamp 1677622389
transform 1 0 4452 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7697
timestamp 1677622389
transform 1 0 4476 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6812
timestamp 1677622389
transform 1 0 4500 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7797
timestamp 1677622389
transform 1 0 4516 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6872
timestamp 1677622389
transform 1 0 4548 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7798
timestamp 1677622389
transform 1 0 4548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7902
timestamp 1677622389
transform 1 0 4548 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6938
timestamp 1677622389
transform 1 0 4540 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7799
timestamp 1677622389
transform 1 0 4572 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6892
timestamp 1677622389
transform 1 0 4580 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7800
timestamp 1677622389
transform 1 0 4588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7903
timestamp 1677622389
transform 1 0 4564 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6911
timestamp 1677622389
transform 1 0 4572 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7904
timestamp 1677622389
transform 1 0 4580 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6939
timestamp 1677622389
transform 1 0 4564 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6839
timestamp 1677622389
transform 1 0 4612 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7698
timestamp 1677622389
transform 1 0 4612 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6893
timestamp 1677622389
transform 1 0 4620 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7905
timestamp 1677622389
transform 1 0 4620 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6912
timestamp 1677622389
transform 1 0 4628 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7801
timestamp 1677622389
transform 1 0 4652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7906
timestamp 1677622389
transform 1 0 4636 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6894
timestamp 1677622389
transform 1 0 4668 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7907
timestamp 1677622389
transform 1 0 4676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6840
timestamp 1677622389
transform 1 0 4700 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6841
timestamp 1677622389
transform 1 0 4732 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7802
timestamp 1677622389
transform 1 0 4732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7803
timestamp 1677622389
transform 1 0 4788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7805
timestamp 1677622389
transform 1 0 4708 0 1 1007
box -2 -2 2 2
use M3_M2  M3_M2_6913
timestamp 1677622389
transform 1 0 4780 0 1 1005
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_74
timestamp 1677622389
transform 1 0 48 0 1 970
box -10 -3 10 3
use INVX2  INVX2_562
timestamp 1677622389
transform 1 0 72 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_326
timestamp 1677622389
transform -1 0 128 0 1 970
box -8 -3 46 105
use FILL  FILL_8905
timestamp 1677622389
transform 1 0 128 0 1 970
box -8 -3 16 105
use FILL  FILL_8912
timestamp 1677622389
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_8914
timestamp 1677622389
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_8916
timestamp 1677622389
transform 1 0 152 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_327
timestamp 1677622389
transform -1 0 200 0 1 970
box -8 -3 46 105
use FILL  FILL_8917
timestamp 1677622389
transform 1 0 200 0 1 970
box -8 -3 16 105
use FILL  FILL_8918
timestamp 1677622389
transform 1 0 208 0 1 970
box -8 -3 16 105
use FILL  FILL_8919
timestamp 1677622389
transform 1 0 216 0 1 970
box -8 -3 16 105
use FILL  FILL_8920
timestamp 1677622389
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_8921
timestamp 1677622389
transform 1 0 232 0 1 970
box -8 -3 16 105
use INVX2  INVX2_564
timestamp 1677622389
transform -1 0 256 0 1 970
box -9 -3 26 105
use FILL  FILL_8922
timestamp 1677622389
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_8923
timestamp 1677622389
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_8924
timestamp 1677622389
transform 1 0 272 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_328
timestamp 1677622389
transform 1 0 280 0 1 970
box -8 -3 46 105
use FILL  FILL_8925
timestamp 1677622389
transform 1 0 320 0 1 970
box -8 -3 16 105
use FILL  FILL_8926
timestamp 1677622389
transform 1 0 328 0 1 970
box -8 -3 16 105
use FILL  FILL_8927
timestamp 1677622389
transform 1 0 336 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_338
timestamp 1677622389
transform 1 0 344 0 1 970
box -8 -3 46 105
use FILL  FILL_8928
timestamp 1677622389
transform 1 0 384 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_486
timestamp 1677622389
transform 1 0 392 0 1 970
box -8 -3 104 105
use FILL  FILL_8929
timestamp 1677622389
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_8930
timestamp 1677622389
transform 1 0 496 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_488
timestamp 1677622389
transform 1 0 504 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_6955
timestamp 1677622389
transform 1 0 612 0 1 975
box -3 -3 3 3
use FILL  FILL_8940
timestamp 1677622389
transform 1 0 600 0 1 970
box -8 -3 16 105
use BUFX2  BUFX2_105
timestamp 1677622389
transform 1 0 608 0 1 970
box -5 -3 28 105
use M3_M2  M3_M2_6956
timestamp 1677622389
transform 1 0 644 0 1 975
box -3 -3 3 3
use FILL  FILL_8941
timestamp 1677622389
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_8952
timestamp 1677622389
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_8954
timestamp 1677622389
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_8956
timestamp 1677622389
transform 1 0 656 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6957
timestamp 1677622389
transform 1 0 692 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_340
timestamp 1677622389
transform 1 0 664 0 1 970
box -8 -3 46 105
use FILL  FILL_8957
timestamp 1677622389
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_8958
timestamp 1677622389
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_8959
timestamp 1677622389
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_8960
timestamp 1677622389
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_8961
timestamp 1677622389
transform 1 0 736 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6958
timestamp 1677622389
transform 1 0 804 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_489
timestamp 1677622389
transform -1 0 840 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_6959
timestamp 1677622389
transform 1 0 852 0 1 975
box -3 -3 3 3
use FILL  FILL_8962
timestamp 1677622389
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_8963
timestamp 1677622389
transform 1 0 848 0 1 970
box -8 -3 16 105
use INVX2  INVX2_570
timestamp 1677622389
transform -1 0 872 0 1 970
box -9 -3 26 105
use FILL  FILL_8964
timestamp 1677622389
transform 1 0 872 0 1 970
box -8 -3 16 105
use FILL  FILL_8971
timestamp 1677622389
transform 1 0 880 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_333
timestamp 1677622389
transform -1 0 928 0 1 970
box -8 -3 46 105
use FILL  FILL_8972
timestamp 1677622389
transform 1 0 928 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6960
timestamp 1677622389
transform 1 0 948 0 1 975
box -3 -3 3 3
use FILL  FILL_8980
timestamp 1677622389
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_8981
timestamp 1677622389
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_8982
timestamp 1677622389
transform 1 0 952 0 1 970
box -8 -3 16 105
use FILL  FILL_8983
timestamp 1677622389
transform 1 0 960 0 1 970
box -8 -3 16 105
use FILL  FILL_8984
timestamp 1677622389
transform 1 0 968 0 1 970
box -8 -3 16 105
use FILL  FILL_8985
timestamp 1677622389
transform 1 0 976 0 1 970
box -8 -3 16 105
use FILL  FILL_8986
timestamp 1677622389
transform 1 0 984 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_89
timestamp 1677622389
transform 1 0 992 0 1 970
box -8 -3 32 105
use FILL  FILL_8987
timestamp 1677622389
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_8988
timestamp 1677622389
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_8989
timestamp 1677622389
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_8991
timestamp 1677622389
transform 1 0 1040 0 1 970
box -8 -3 16 105
use FILL  FILL_8993
timestamp 1677622389
transform 1 0 1048 0 1 970
box -8 -3 16 105
use FILL  FILL_8994
timestamp 1677622389
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_8995
timestamp 1677622389
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_8996
timestamp 1677622389
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_8999
timestamp 1677622389
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_9001
timestamp 1677622389
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_9003
timestamp 1677622389
transform 1 0 1096 0 1 970
box -8 -3 16 105
use FILL  FILL_9005
timestamp 1677622389
transform 1 0 1104 0 1 970
box -8 -3 16 105
use FILL  FILL_9007
timestamp 1677622389
transform 1 0 1112 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6961
timestamp 1677622389
transform 1 0 1140 0 1 975
box -3 -3 3 3
use NOR2X1  NOR2X1_90
timestamp 1677622389
transform 1 0 1120 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_6962
timestamp 1677622389
transform 1 0 1156 0 1 975
box -3 -3 3 3
use FILL  FILL_9009
timestamp 1677622389
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_9010
timestamp 1677622389
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_9011
timestamp 1677622389
transform 1 0 1160 0 1 970
box -8 -3 16 105
use FILL  FILL_9013
timestamp 1677622389
transform 1 0 1168 0 1 970
box -8 -3 16 105
use FILL  FILL_9015
timestamp 1677622389
transform 1 0 1176 0 1 970
box -8 -3 16 105
use FILL  FILL_9017
timestamp 1677622389
transform 1 0 1184 0 1 970
box -8 -3 16 105
use FILL  FILL_9019
timestamp 1677622389
transform 1 0 1192 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_342
timestamp 1677622389
transform -1 0 1240 0 1 970
box -8 -3 46 105
use FILL  FILL_9020
timestamp 1677622389
transform 1 0 1240 0 1 970
box -8 -3 16 105
use FILL  FILL_9021
timestamp 1677622389
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_9025
timestamp 1677622389
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_9027
timestamp 1677622389
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_9028
timestamp 1677622389
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_9029
timestamp 1677622389
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_9030
timestamp 1677622389
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_9031
timestamp 1677622389
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_9032
timestamp 1677622389
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_9033
timestamp 1677622389
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_9034
timestamp 1677622389
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_9035
timestamp 1677622389
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_9036
timestamp 1677622389
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_9037
timestamp 1677622389
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_9038
timestamp 1677622389
transform 1 0 1352 0 1 970
box -8 -3 16 105
use INVX2  INVX2_572
timestamp 1677622389
transform -1 0 1376 0 1 970
box -9 -3 26 105
use FILL  FILL_9039
timestamp 1677622389
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_9040
timestamp 1677622389
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_9041
timestamp 1677622389
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_9042
timestamp 1677622389
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_9043
timestamp 1677622389
transform 1 0 1408 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_335
timestamp 1677622389
transform -1 0 1456 0 1 970
box -8 -3 46 105
use FILL  FILL_9044
timestamp 1677622389
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_9053
timestamp 1677622389
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_9054
timestamp 1677622389
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_9055
timestamp 1677622389
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_9056
timestamp 1677622389
transform 1 0 1488 0 1 970
box -8 -3 16 105
use FILL  FILL_9057
timestamp 1677622389
transform 1 0 1496 0 1 970
box -8 -3 16 105
use FILL  FILL_9058
timestamp 1677622389
transform 1 0 1504 0 1 970
box -8 -3 16 105
use INVX2  INVX2_573
timestamp 1677622389
transform 1 0 1512 0 1 970
box -9 -3 26 105
use FILL  FILL_9059
timestamp 1677622389
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_9064
timestamp 1677622389
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_9066
timestamp 1677622389
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_9068
timestamp 1677622389
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_9069
timestamp 1677622389
transform 1 0 1560 0 1 970
box -8 -3 16 105
use INVX2  INVX2_574
timestamp 1677622389
transform 1 0 1568 0 1 970
box -9 -3 26 105
use FILL  FILL_9070
timestamp 1677622389
transform 1 0 1584 0 1 970
box -8 -3 16 105
use FILL  FILL_9071
timestamp 1677622389
transform 1 0 1592 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6963
timestamp 1677622389
transform 1 0 1612 0 1 975
box -3 -3 3 3
use FILL  FILL_9072
timestamp 1677622389
transform 1 0 1600 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_345
timestamp 1677622389
transform 1 0 1608 0 1 970
box -8 -3 46 105
use BUFX2  BUFX2_106
timestamp 1677622389
transform -1 0 1672 0 1 970
box -5 -3 28 105
use FILL  FILL_9073
timestamp 1677622389
transform 1 0 1672 0 1 970
box -8 -3 16 105
use FILL  FILL_9074
timestamp 1677622389
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_9075
timestamp 1677622389
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_9076
timestamp 1677622389
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_9077
timestamp 1677622389
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_9078
timestamp 1677622389
transform 1 0 1712 0 1 970
box -8 -3 16 105
use FILL  FILL_9083
timestamp 1677622389
transform 1 0 1720 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_346
timestamp 1677622389
transform 1 0 1728 0 1 970
box -8 -3 46 105
use FILL  FILL_9085
timestamp 1677622389
transform 1 0 1768 0 1 970
box -8 -3 16 105
use FILL  FILL_9086
timestamp 1677622389
transform 1 0 1776 0 1 970
box -8 -3 16 105
use FILL  FILL_9087
timestamp 1677622389
transform 1 0 1784 0 1 970
box -8 -3 16 105
use FILL  FILL_9088
timestamp 1677622389
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_9089
timestamp 1677622389
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_9090
timestamp 1677622389
transform 1 0 1808 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_338
timestamp 1677622389
transform -1 0 1856 0 1 970
box -8 -3 46 105
use FILL  FILL_9091
timestamp 1677622389
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_9092
timestamp 1677622389
transform 1 0 1864 0 1 970
box -8 -3 16 105
use FILL  FILL_9093
timestamp 1677622389
transform 1 0 1872 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_494
timestamp 1677622389
transform -1 0 1976 0 1 970
box -8 -3 104 105
use FILL  FILL_9094
timestamp 1677622389
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_9095
timestamp 1677622389
transform 1 0 1984 0 1 970
box -8 -3 16 105
use INVX2  INVX2_575
timestamp 1677622389
transform -1 0 2008 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_6964
timestamp 1677622389
transform 1 0 2020 0 1 975
box -3 -3 3 3
use FILL  FILL_9096
timestamp 1677622389
transform 1 0 2008 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6965
timestamp 1677622389
transform 1 0 2044 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_339
timestamp 1677622389
transform -1 0 2056 0 1 970
box -8 -3 46 105
use FILL  FILL_9097
timestamp 1677622389
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_9098
timestamp 1677622389
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_9099
timestamp 1677622389
transform 1 0 2072 0 1 970
box -8 -3 16 105
use INVX2  INVX2_576
timestamp 1677622389
transform -1 0 2096 0 1 970
box -9 -3 26 105
use FILL  FILL_9100
timestamp 1677622389
transform 1 0 2096 0 1 970
box -8 -3 16 105
use FILL  FILL_9101
timestamp 1677622389
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_9102
timestamp 1677622389
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_9103
timestamp 1677622389
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_9104
timestamp 1677622389
transform 1 0 2128 0 1 970
box -8 -3 16 105
use FILL  FILL_9114
timestamp 1677622389
transform 1 0 2136 0 1 970
box -8 -3 16 105
use FILL  FILL_9116
timestamp 1677622389
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_9118
timestamp 1677622389
transform 1 0 2152 0 1 970
box -8 -3 16 105
use FILL  FILL_9120
timestamp 1677622389
transform 1 0 2160 0 1 970
box -8 -3 16 105
use INVX2  INVX2_579
timestamp 1677622389
transform -1 0 2184 0 1 970
box -9 -3 26 105
use FILL  FILL_9121
timestamp 1677622389
transform 1 0 2184 0 1 970
box -8 -3 16 105
use FILL  FILL_9124
timestamp 1677622389
transform 1 0 2192 0 1 970
box -8 -3 16 105
use FILL  FILL_9126
timestamp 1677622389
transform 1 0 2200 0 1 970
box -8 -3 16 105
use FILL  FILL_9127
timestamp 1677622389
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_9128
timestamp 1677622389
transform 1 0 2216 0 1 970
box -8 -3 16 105
use INVX2  INVX2_581
timestamp 1677622389
transform -1 0 2240 0 1 970
box -9 -3 26 105
use FILL  FILL_9129
timestamp 1677622389
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_9130
timestamp 1677622389
transform 1 0 2248 0 1 970
box -8 -3 16 105
use INVX2  INVX2_582
timestamp 1677622389
transform 1 0 2256 0 1 970
box -9 -3 26 105
use FILL  FILL_9131
timestamp 1677622389
transform 1 0 2272 0 1 970
box -8 -3 16 105
use FILL  FILL_9132
timestamp 1677622389
transform 1 0 2280 0 1 970
box -8 -3 16 105
use FILL  FILL_9133
timestamp 1677622389
transform 1 0 2288 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_20
timestamp 1677622389
transform 1 0 2296 0 1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_153
timestamp 1677622389
transform -1 0 2352 0 1 970
box -8 -3 34 105
use FILL  FILL_9134
timestamp 1677622389
transform 1 0 2352 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_21
timestamp 1677622389
transform -1 0 2384 0 1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_154
timestamp 1677622389
transform -1 0 2416 0 1 970
box -8 -3 34 105
use FILL  FILL_9135
timestamp 1677622389
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_9149
timestamp 1677622389
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_9151
timestamp 1677622389
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_9153
timestamp 1677622389
transform 1 0 2440 0 1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_13
timestamp 1677622389
transform -1 0 2480 0 1 970
box -7 -3 39 105
use FILL  FILL_9154
timestamp 1677622389
transform 1 0 2480 0 1 970
box -8 -3 16 105
use FILL  FILL_9155
timestamp 1677622389
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_9159
timestamp 1677622389
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_9161
timestamp 1677622389
transform 1 0 2504 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_53
timestamp 1677622389
transform 1 0 2512 0 1 970
box -8 -3 40 105
use XOR2X1  XOR2X1_2
timestamp 1677622389
transform 1 0 2544 0 1 970
box -8 -3 64 105
use FILL  FILL_9163
timestamp 1677622389
transform 1 0 2600 0 1 970
box -8 -3 16 105
use FILL  FILL_9167
timestamp 1677622389
transform 1 0 2608 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_342
timestamp 1677622389
transform 1 0 2616 0 1 970
box -8 -3 46 105
use FILL  FILL_9169
timestamp 1677622389
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_9170
timestamp 1677622389
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_9171
timestamp 1677622389
transform 1 0 2672 0 1 970
box -8 -3 16 105
use INVX2  INVX2_584
timestamp 1677622389
transform -1 0 2696 0 1 970
box -9 -3 26 105
use FILL  FILL_9172
timestamp 1677622389
transform 1 0 2696 0 1 970
box -8 -3 16 105
use FILL  FILL_9173
timestamp 1677622389
transform 1 0 2704 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6966
timestamp 1677622389
transform 1 0 2796 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_498
timestamp 1677622389
transform -1 0 2808 0 1 970
box -8 -3 104 105
use FILL  FILL_9174
timestamp 1677622389
transform 1 0 2808 0 1 970
box -8 -3 16 105
use FILL  FILL_9175
timestamp 1677622389
transform 1 0 2816 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6967
timestamp 1677622389
transform 1 0 2852 0 1 975
box -3 -3 3 3
use FAX1  FAX1_16
timestamp 1677622389
transform 1 0 2824 0 1 970
box -5 -3 126 105
use FILL  FILL_9176
timestamp 1677622389
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_9177
timestamp 1677622389
transform 1 0 2952 0 1 970
box -8 -3 16 105
use FILL  FILL_9178
timestamp 1677622389
transform 1 0 2960 0 1 970
box -8 -3 16 105
use FILL  FILL_9179
timestamp 1677622389
transform 1 0 2968 0 1 970
box -8 -3 16 105
use FILL  FILL_9180
timestamp 1677622389
transform 1 0 2976 0 1 970
box -8 -3 16 105
use FILL  FILL_9181
timestamp 1677622389
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_9182
timestamp 1677622389
transform 1 0 2992 0 1 970
box -8 -3 16 105
use FILL  FILL_9187
timestamp 1677622389
transform 1 0 3000 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_23
timestamp 1677622389
transform 1 0 3008 0 1 970
box -8 -3 32 105
use FILL  FILL_9189
timestamp 1677622389
transform 1 0 3032 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_24
timestamp 1677622389
transform 1 0 3040 0 1 970
box -8 -3 32 105
use FILL  FILL_9190
timestamp 1677622389
transform 1 0 3064 0 1 970
box -8 -3 16 105
use FILL  FILL_9196
timestamp 1677622389
transform 1 0 3072 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1677622389
transform 1 0 3080 0 1 970
box -8 -3 40 105
use FILL  FILL_9198
timestamp 1677622389
transform 1 0 3112 0 1 970
box -8 -3 16 105
use FILL  FILL_9200
timestamp 1677622389
transform 1 0 3120 0 1 970
box -8 -3 16 105
use FILL  FILL_9202
timestamp 1677622389
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_9204
timestamp 1677622389
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_9206
timestamp 1677622389
transform 1 0 3144 0 1 970
box -8 -3 16 105
use FILL  FILL_9207
timestamp 1677622389
transform 1 0 3152 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_155
timestamp 1677622389
transform -1 0 3192 0 1 970
box -8 -3 34 105
use FILL  FILL_9208
timestamp 1677622389
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_9212
timestamp 1677622389
transform 1 0 3200 0 1 970
box -8 -3 16 105
use INVX2  INVX2_585
timestamp 1677622389
transform -1 0 3224 0 1 970
box -9 -3 26 105
use FILL  FILL_9213
timestamp 1677622389
transform 1 0 3224 0 1 970
box -8 -3 16 105
use FILL  FILL_9218
timestamp 1677622389
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_9220
timestamp 1677622389
transform 1 0 3240 0 1 970
box -8 -3 16 105
use FILL  FILL_9222
timestamp 1677622389
transform 1 0 3248 0 1 970
box -8 -3 16 105
use FILL  FILL_9224
timestamp 1677622389
transform 1 0 3256 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_344
timestamp 1677622389
transform -1 0 3304 0 1 970
box -8 -3 46 105
use FILL  FILL_9225
timestamp 1677622389
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_9226
timestamp 1677622389
transform 1 0 3312 0 1 970
box -8 -3 16 105
use FILL  FILL_9230
timestamp 1677622389
transform 1 0 3320 0 1 970
box -8 -3 16 105
use FILL  FILL_9232
timestamp 1677622389
transform 1 0 3328 0 1 970
box -8 -3 16 105
use FILL  FILL_9234
timestamp 1677622389
transform 1 0 3336 0 1 970
box -8 -3 16 105
use FILL  FILL_9236
timestamp 1677622389
transform 1 0 3344 0 1 970
box -8 -3 16 105
use FILL  FILL_9237
timestamp 1677622389
transform 1 0 3352 0 1 970
box -8 -3 16 105
use FILL  FILL_9238
timestamp 1677622389
transform 1 0 3360 0 1 970
box -8 -3 16 105
use FILL  FILL_9239
timestamp 1677622389
transform 1 0 3368 0 1 970
box -8 -3 16 105
use FILL  FILL_9240
timestamp 1677622389
transform 1 0 3376 0 1 970
box -8 -3 16 105
use FILL  FILL_9241
timestamp 1677622389
transform 1 0 3384 0 1 970
box -8 -3 16 105
use FAX1  FAX1_18
timestamp 1677622389
transform 1 0 3392 0 1 970
box -5 -3 126 105
use FILL  FILL_9243
timestamp 1677622389
transform 1 0 3512 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_54
timestamp 1677622389
transform -1 0 3552 0 1 970
box -8 -3 40 105
use FILL  FILL_9244
timestamp 1677622389
transform 1 0 3552 0 1 970
box -8 -3 16 105
use FILL  FILL_9258
timestamp 1677622389
transform 1 0 3560 0 1 970
box -8 -3 16 105
use FILL  FILL_9260
timestamp 1677622389
transform 1 0 3568 0 1 970
box -8 -3 16 105
use FILL  FILL_9261
timestamp 1677622389
transform 1 0 3576 0 1 970
box -8 -3 16 105
use FILL  FILL_9262
timestamp 1677622389
transform 1 0 3584 0 1 970
box -8 -3 16 105
use FILL  FILL_9263
timestamp 1677622389
transform 1 0 3592 0 1 970
box -8 -3 16 105
use FILL  FILL_9264
timestamp 1677622389
transform 1 0 3600 0 1 970
box -8 -3 16 105
use FILL  FILL_9265
timestamp 1677622389
transform 1 0 3608 0 1 970
box -8 -3 16 105
use FILL  FILL_9266
timestamp 1677622389
transform 1 0 3616 0 1 970
box -8 -3 16 105
use FILL  FILL_9267
timestamp 1677622389
transform 1 0 3624 0 1 970
box -8 -3 16 105
use FILL  FILL_9268
timestamp 1677622389
transform 1 0 3632 0 1 970
box -8 -3 16 105
use FILL  FILL_9271
timestamp 1677622389
transform 1 0 3640 0 1 970
box -8 -3 16 105
use FILL  FILL_9272
timestamp 1677622389
transform 1 0 3648 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_347
timestamp 1677622389
transform 1 0 3656 0 1 970
box -8 -3 46 105
use FILL  FILL_9273
timestamp 1677622389
transform 1 0 3696 0 1 970
box -8 -3 16 105
use FILL  FILL_9278
timestamp 1677622389
transform 1 0 3704 0 1 970
box -8 -3 16 105
use FILL  FILL_9280
timestamp 1677622389
transform 1 0 3712 0 1 970
box -8 -3 16 105
use FILL  FILL_9281
timestamp 1677622389
transform 1 0 3720 0 1 970
box -8 -3 16 105
use FILL  FILL_9282
timestamp 1677622389
transform 1 0 3728 0 1 970
box -8 -3 16 105
use FILL  FILL_9283
timestamp 1677622389
transform 1 0 3736 0 1 970
box -8 -3 16 105
use FILL  FILL_9284
timestamp 1677622389
transform 1 0 3744 0 1 970
box -8 -3 16 105
use FILL  FILL_9287
timestamp 1677622389
transform 1 0 3752 0 1 970
box -8 -3 16 105
use FILL  FILL_9289
timestamp 1677622389
transform 1 0 3760 0 1 970
box -8 -3 16 105
use FILL  FILL_9291
timestamp 1677622389
transform 1 0 3768 0 1 970
box -8 -3 16 105
use FILL  FILL_9293
timestamp 1677622389
transform 1 0 3776 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_348
timestamp 1677622389
transform 1 0 3784 0 1 970
box -8 -3 46 105
use FILL  FILL_9295
timestamp 1677622389
transform 1 0 3824 0 1 970
box -8 -3 16 105
use FILL  FILL_9298
timestamp 1677622389
transform 1 0 3832 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6968
timestamp 1677622389
transform 1 0 3860 0 1 975
box -3 -3 3 3
use NAND2X1  NAND2X1_28
timestamp 1677622389
transform -1 0 3864 0 1 970
box -8 -3 32 105
use FILL  FILL_9299
timestamp 1677622389
transform 1 0 3864 0 1 970
box -8 -3 16 105
use FILL  FILL_9300
timestamp 1677622389
transform 1 0 3872 0 1 970
box -8 -3 16 105
use FILL  FILL_9301
timestamp 1677622389
transform 1 0 3880 0 1 970
box -8 -3 16 105
use FILL  FILL_9306
timestamp 1677622389
transform 1 0 3888 0 1 970
box -8 -3 16 105
use FILL  FILL_9308
timestamp 1677622389
transform 1 0 3896 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_349
timestamp 1677622389
transform -1 0 3944 0 1 970
box -8 -3 46 105
use FILL  FILL_9309
timestamp 1677622389
transform 1 0 3944 0 1 970
box -8 -3 16 105
use FILL  FILL_9310
timestamp 1677622389
transform 1 0 3952 0 1 970
box -8 -3 16 105
use FILL  FILL_9311
timestamp 1677622389
transform 1 0 3960 0 1 970
box -8 -3 16 105
use FILL  FILL_9317
timestamp 1677622389
transform 1 0 3968 0 1 970
box -8 -3 16 105
use FILL  FILL_9319
timestamp 1677622389
transform 1 0 3976 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_350
timestamp 1677622389
transform -1 0 4024 0 1 970
box -8 -3 46 105
use FILL  FILL_9320
timestamp 1677622389
transform 1 0 4024 0 1 970
box -8 -3 16 105
use FILL  FILL_9325
timestamp 1677622389
transform 1 0 4032 0 1 970
box -8 -3 16 105
use FILL  FILL_9327
timestamp 1677622389
transform 1 0 4040 0 1 970
box -8 -3 16 105
use FILL  FILL_9329
timestamp 1677622389
transform 1 0 4048 0 1 970
box -8 -3 16 105
use FILL  FILL_9331
timestamp 1677622389
transform 1 0 4056 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_351
timestamp 1677622389
transform 1 0 4064 0 1 970
box -8 -3 46 105
use FILL  FILL_9332
timestamp 1677622389
transform 1 0 4104 0 1 970
box -8 -3 16 105
use FILL  FILL_9336
timestamp 1677622389
transform 1 0 4112 0 1 970
box -8 -3 16 105
use FILL  FILL_9338
timestamp 1677622389
transform 1 0 4120 0 1 970
box -8 -3 16 105
use FILL  FILL_9340
timestamp 1677622389
transform 1 0 4128 0 1 970
box -8 -3 16 105
use FILL  FILL_9341
timestamp 1677622389
transform 1 0 4136 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_352
timestamp 1677622389
transform -1 0 4184 0 1 970
box -8 -3 46 105
use FILL  FILL_9342
timestamp 1677622389
transform 1 0 4184 0 1 970
box -8 -3 16 105
use FILL  FILL_9344
timestamp 1677622389
transform 1 0 4192 0 1 970
box -8 -3 16 105
use FILL  FILL_9346
timestamp 1677622389
transform 1 0 4200 0 1 970
box -8 -3 16 105
use FILL  FILL_9348
timestamp 1677622389
transform 1 0 4208 0 1 970
box -8 -3 16 105
use FILL  FILL_9349
timestamp 1677622389
transform 1 0 4216 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_353
timestamp 1677622389
transform 1 0 4224 0 1 970
box -8 -3 46 105
use FILL  FILL_9350
timestamp 1677622389
transform 1 0 4264 0 1 970
box -8 -3 16 105
use FILL  FILL_9355
timestamp 1677622389
transform 1 0 4272 0 1 970
box -8 -3 16 105
use FILL  FILL_9357
timestamp 1677622389
transform 1 0 4280 0 1 970
box -8 -3 16 105
use FILL  FILL_9359
timestamp 1677622389
transform 1 0 4288 0 1 970
box -8 -3 16 105
use FILL  FILL_9361
timestamp 1677622389
transform 1 0 4296 0 1 970
box -8 -3 16 105
use FILL  FILL_9362
timestamp 1677622389
transform 1 0 4304 0 1 970
box -8 -3 16 105
use FILL  FILL_9363
timestamp 1677622389
transform 1 0 4312 0 1 970
box -8 -3 16 105
use FILL  FILL_9364
timestamp 1677622389
transform 1 0 4320 0 1 970
box -8 -3 16 105
use FILL  FILL_9365
timestamp 1677622389
transform 1 0 4328 0 1 970
box -8 -3 16 105
use FILL  FILL_9366
timestamp 1677622389
transform 1 0 4336 0 1 970
box -8 -3 16 105
use FILL  FILL_9369
timestamp 1677622389
transform 1 0 4344 0 1 970
box -8 -3 16 105
use FILL  FILL_9371
timestamp 1677622389
transform 1 0 4352 0 1 970
box -8 -3 16 105
use FILL  FILL_9373
timestamp 1677622389
transform 1 0 4360 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_164
timestamp 1677622389
transform -1 0 4400 0 1 970
box -8 -3 34 105
use FILL  FILL_9374
timestamp 1677622389
transform 1 0 4400 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_165
timestamp 1677622389
transform -1 0 4440 0 1 970
box -8 -3 34 105
use FILL  FILL_9381
timestamp 1677622389
transform 1 0 4440 0 1 970
box -8 -3 16 105
use FILL  FILL_9383
timestamp 1677622389
transform 1 0 4448 0 1 970
box -8 -3 16 105
use FILL  FILL_9385
timestamp 1677622389
transform 1 0 4456 0 1 970
box -8 -3 16 105
use FILL  FILL_9387
timestamp 1677622389
transform 1 0 4464 0 1 970
box -8 -3 16 105
use FILL  FILL_9388
timestamp 1677622389
transform 1 0 4472 0 1 970
box -8 -3 16 105
use FILL  FILL_9389
timestamp 1677622389
transform 1 0 4480 0 1 970
box -8 -3 16 105
use FILL  FILL_9390
timestamp 1677622389
transform 1 0 4488 0 1 970
box -8 -3 16 105
use FILL  FILL_9391
timestamp 1677622389
transform 1 0 4496 0 1 970
box -8 -3 16 105
use FILL  FILL_9392
timestamp 1677622389
transform 1 0 4504 0 1 970
box -8 -3 16 105
use FILL  FILL_9395
timestamp 1677622389
transform 1 0 4512 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_168
timestamp 1677622389
transform -1 0 4552 0 1 970
box -8 -3 34 105
use FILL  FILL_9396
timestamp 1677622389
transform 1 0 4552 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_354
timestamp 1677622389
transform 1 0 4560 0 1 970
box -8 -3 46 105
use FILL  FILL_9403
timestamp 1677622389
transform 1 0 4600 0 1 970
box -8 -3 16 105
use FILL  FILL_9410
timestamp 1677622389
transform 1 0 4608 0 1 970
box -8 -3 16 105
use FILL  FILL_9412
timestamp 1677622389
transform 1 0 4616 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_6969
timestamp 1677622389
transform 1 0 4636 0 1 975
box -3 -3 3 3
use FILL  FILL_9414
timestamp 1677622389
transform 1 0 4624 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_169
timestamp 1677622389
transform -1 0 4664 0 1 970
box -8 -3 34 105
use FILL  FILL_9415
timestamp 1677622389
transform 1 0 4664 0 1 970
box -8 -3 16 105
use FILL  FILL_9422
timestamp 1677622389
transform 1 0 4672 0 1 970
box -8 -3 16 105
use FILL  FILL_9424
timestamp 1677622389
transform 1 0 4680 0 1 970
box -8 -3 16 105
use FILL  FILL_9425
timestamp 1677622389
transform 1 0 4688 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_501
timestamp 1677622389
transform 1 0 4696 0 1 970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_75
timestamp 1677622389
transform 1 0 4819 0 1 970
box -10 -3 10 3
use M2_M1  M2_M1_7914
timestamp 1677622389
transform 1 0 108 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7071
timestamp 1677622389
transform 1 0 100 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8013
timestamp 1677622389
transform 1 0 116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7915
timestamp 1677622389
transform 1 0 132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7916
timestamp 1677622389
transform 1 0 148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8014
timestamp 1677622389
transform 1 0 156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7917
timestamp 1677622389
transform 1 0 188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8015
timestamp 1677622389
transform 1 0 172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8016
timestamp 1677622389
transform 1 0 236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8017
timestamp 1677622389
transform 1 0 268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8018
timestamp 1677622389
transform 1 0 276 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7072
timestamp 1677622389
transform 1 0 164 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7073
timestamp 1677622389
transform 1 0 236 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7074
timestamp 1677622389
transform 1 0 276 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7110
timestamp 1677622389
transform 1 0 188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7111
timestamp 1677622389
transform 1 0 220 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7112
timestamp 1677622389
transform 1 0 268 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7918
timestamp 1677622389
transform 1 0 308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7919
timestamp 1677622389
transform 1 0 316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7920
timestamp 1677622389
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8019
timestamp 1677622389
transform 1 0 300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7921
timestamp 1677622389
transform 1 0 348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8020
timestamp 1677622389
transform 1 0 324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8021
timestamp 1677622389
transform 1 0 340 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7075
timestamp 1677622389
transform 1 0 340 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7113
timestamp 1677622389
transform 1 0 316 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7922
timestamp 1677622389
transform 1 0 372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7923
timestamp 1677622389
transform 1 0 388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8022
timestamp 1677622389
transform 1 0 356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8023
timestamp 1677622389
transform 1 0 380 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7114
timestamp 1677622389
transform 1 0 348 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7040
timestamp 1677622389
transform 1 0 388 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8024
timestamp 1677622389
transform 1 0 396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7924
timestamp 1677622389
transform 1 0 436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8025
timestamp 1677622389
transform 1 0 444 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7001
timestamp 1677622389
transform 1 0 484 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7925
timestamp 1677622389
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7926
timestamp 1677622389
transform 1 0 468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7927
timestamp 1677622389
transform 1 0 484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8026
timestamp 1677622389
transform 1 0 460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7041
timestamp 1677622389
transform 1 0 468 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8027
timestamp 1677622389
transform 1 0 476 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7076
timestamp 1677622389
transform 1 0 460 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8028
timestamp 1677622389
transform 1 0 516 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7077
timestamp 1677622389
transform 1 0 516 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7042
timestamp 1677622389
transform 1 0 540 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7928
timestamp 1677622389
transform 1 0 572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7929
timestamp 1677622389
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7930
timestamp 1677622389
transform 1 0 596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8029
timestamp 1677622389
transform 1 0 548 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7043
timestamp 1677622389
transform 1 0 556 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8030
timestamp 1677622389
transform 1 0 572 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7044
timestamp 1677622389
transform 1 0 580 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8031
timestamp 1677622389
transform 1 0 588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8032
timestamp 1677622389
transform 1 0 604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7078
timestamp 1677622389
transform 1 0 564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7142
timestamp 1677622389
transform 1 0 572 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7079
timestamp 1677622389
transform 1 0 604 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_6980
timestamp 1677622389
transform 1 0 668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6981
timestamp 1677622389
transform 1 0 740 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7931
timestamp 1677622389
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8033
timestamp 1677622389
transform 1 0 716 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7143
timestamp 1677622389
transform 1 0 684 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7002
timestamp 1677622389
transform 1 0 756 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7932
timestamp 1677622389
transform 1 0 756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7933
timestamp 1677622389
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8034
timestamp 1677622389
transform 1 0 780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8035
timestamp 1677622389
transform 1 0 788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8036
timestamp 1677622389
transform 1 0 804 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6982
timestamp 1677622389
transform 1 0 836 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7003
timestamp 1677622389
transform 1 0 820 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7004
timestamp 1677622389
transform 1 0 852 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7934
timestamp 1677622389
transform 1 0 820 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7023
timestamp 1677622389
transform 1 0 828 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7935
timestamp 1677622389
transform 1 0 836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7936
timestamp 1677622389
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8037
timestamp 1677622389
transform 1 0 820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8038
timestamp 1677622389
transform 1 0 828 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7045
timestamp 1677622389
transform 1 0 836 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8039
timestamp 1677622389
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8040
timestamp 1677622389
transform 1 0 860 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7115
timestamp 1677622389
transform 1 0 820 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7937
timestamp 1677622389
transform 1 0 884 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7046
timestamp 1677622389
transform 1 0 916 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7938
timestamp 1677622389
transform 1 0 948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8041
timestamp 1677622389
transform 1 0 996 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7047
timestamp 1677622389
transform 1 0 1020 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8042
timestamp 1677622389
transform 1 0 1028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8043
timestamp 1677622389
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7080
timestamp 1677622389
transform 1 0 996 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7081
timestamp 1677622389
transform 1 0 1036 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8044
timestamp 1677622389
transform 1 0 1076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7939
timestamp 1677622389
transform 1 0 1124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7940
timestamp 1677622389
transform 1 0 1132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7941
timestamp 1677622389
transform 1 0 1148 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7161
timestamp 1677622389
transform 1 0 1116 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8045
timestamp 1677622389
transform 1 0 1140 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7048
timestamp 1677622389
transform 1 0 1148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7144
timestamp 1677622389
transform 1 0 1132 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8046
timestamp 1677622389
transform 1 0 1164 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7116
timestamp 1677622389
transform 1 0 1164 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7942
timestamp 1677622389
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7943
timestamp 1677622389
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8047
timestamp 1677622389
transform 1 0 1220 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7049
timestamp 1677622389
transform 1 0 1228 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8048
timestamp 1677622389
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7082
timestamp 1677622389
transform 1 0 1220 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7117
timestamp 1677622389
transform 1 0 1220 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8049
timestamp 1677622389
transform 1 0 1252 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7145
timestamp 1677622389
transform 1 0 1244 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7005
timestamp 1677622389
transform 1 0 1268 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7944
timestamp 1677622389
transform 1 0 1268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7945
timestamp 1677622389
transform 1 0 1356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8050
timestamp 1677622389
transform 1 0 1332 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7083
timestamp 1677622389
transform 1 0 1276 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7118
timestamp 1677622389
transform 1 0 1356 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7946
timestamp 1677622389
transform 1 0 1372 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7006
timestamp 1677622389
transform 1 0 1428 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7947
timestamp 1677622389
transform 1 0 1404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7948
timestamp 1677622389
transform 1 0 1420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7949
timestamp 1677622389
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8051
timestamp 1677622389
transform 1 0 1396 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7162
timestamp 1677622389
transform 1 0 1404 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7950
timestamp 1677622389
transform 1 0 1484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7951
timestamp 1677622389
transform 1 0 1500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7952
timestamp 1677622389
transform 1 0 1508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8052
timestamp 1677622389
transform 1 0 1468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8053
timestamp 1677622389
transform 1 0 1476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8054
timestamp 1677622389
transform 1 0 1492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7084
timestamp 1677622389
transform 1 0 1468 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7050
timestamp 1677622389
transform 1 0 1500 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7119
timestamp 1677622389
transform 1 0 1476 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8055
timestamp 1677622389
transform 1 0 1524 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7007
timestamp 1677622389
transform 1 0 1564 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7008
timestamp 1677622389
transform 1 0 1604 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7009
timestamp 1677622389
transform 1 0 1644 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7953
timestamp 1677622389
transform 1 0 1564 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7024
timestamp 1677622389
transform 1 0 1652 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8056
timestamp 1677622389
transform 1 0 1588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8057
timestamp 1677622389
transform 1 0 1644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8058
timestamp 1677622389
transform 1 0 1652 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7085
timestamp 1677622389
transform 1 0 1644 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7120
timestamp 1677622389
transform 1 0 1668 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7010
timestamp 1677622389
transform 1 0 1700 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7954
timestamp 1677622389
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7955
timestamp 1677622389
transform 1 0 1700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8059
timestamp 1677622389
transform 1 0 1692 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7146
timestamp 1677622389
transform 1 0 1684 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8060
timestamp 1677622389
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7051
timestamp 1677622389
transform 1 0 1732 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_6983
timestamp 1677622389
transform 1 0 1868 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6984
timestamp 1677622389
transform 1 0 1884 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7011
timestamp 1677622389
transform 1 0 1788 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7012
timestamp 1677622389
transform 1 0 1804 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7956
timestamp 1677622389
transform 1 0 1764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7957
timestamp 1677622389
transform 1 0 1772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7958
timestamp 1677622389
transform 1 0 1788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8061
timestamp 1677622389
transform 1 0 1756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8062
timestamp 1677622389
transform 1 0 1764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8063
timestamp 1677622389
transform 1 0 1780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7086
timestamp 1677622389
transform 1 0 1756 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7052
timestamp 1677622389
transform 1 0 1788 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7959
timestamp 1677622389
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8064
timestamp 1677622389
transform 1 0 1796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8065
timestamp 1677622389
transform 1 0 1804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8066
timestamp 1677622389
transform 1 0 1836 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7147
timestamp 1677622389
transform 1 0 1772 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7087
timestamp 1677622389
transform 1 0 1836 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7088
timestamp 1677622389
transform 1 0 1884 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7148
timestamp 1677622389
transform 1 0 1844 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7163
timestamp 1677622389
transform 1 0 1828 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7960
timestamp 1677622389
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7961
timestamp 1677622389
transform 1 0 1956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7962
timestamp 1677622389
transform 1 0 2044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7963
timestamp 1677622389
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7053
timestamp 1677622389
transform 1 0 1932 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8067
timestamp 1677622389
transform 1 0 1940 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7054
timestamp 1677622389
transform 1 0 1956 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7025
timestamp 1677622389
transform 1 0 2076 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8068
timestamp 1677622389
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8069
timestamp 1677622389
transform 1 0 2036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8070
timestamp 1677622389
transform 1 0 2044 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8071
timestamp 1677622389
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8072
timestamp 1677622389
transform 1 0 2076 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7089
timestamp 1677622389
transform 1 0 1924 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7090
timestamp 1677622389
transform 1 0 1940 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7091
timestamp 1677622389
transform 1 0 1980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7092
timestamp 1677622389
transform 1 0 2028 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7093
timestamp 1677622389
transform 1 0 2044 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7121
timestamp 1677622389
transform 1 0 2004 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8123
timestamp 1677622389
transform 1 0 2084 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7122
timestamp 1677622389
transform 1 0 2084 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8073
timestamp 1677622389
transform 1 0 2116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8144
timestamp 1677622389
transform 1 0 2108 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_7964
timestamp 1677622389
transform 1 0 2132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8074
timestamp 1677622389
transform 1 0 2156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8075
timestamp 1677622389
transform 1 0 2164 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7013
timestamp 1677622389
transform 1 0 2188 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7026
timestamp 1677622389
transform 1 0 2196 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8076
timestamp 1677622389
transform 1 0 2196 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6970
timestamp 1677622389
transform 1 0 2252 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6971
timestamp 1677622389
transform 1 0 2292 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6985
timestamp 1677622389
transform 1 0 2212 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6986
timestamp 1677622389
transform 1 0 2236 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7014
timestamp 1677622389
transform 1 0 2212 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7015
timestamp 1677622389
transform 1 0 2260 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7965
timestamp 1677622389
transform 1 0 2212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7027
timestamp 1677622389
transform 1 0 2276 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8077
timestamp 1677622389
transform 1 0 2260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8078
timestamp 1677622389
transform 1 0 2292 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7016
timestamp 1677622389
transform 1 0 2308 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7017
timestamp 1677622389
transform 1 0 2324 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7966
timestamp 1677622389
transform 1 0 2316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8079
timestamp 1677622389
transform 1 0 2308 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7055
timestamp 1677622389
transform 1 0 2316 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8124
timestamp 1677622389
transform 1 0 2332 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7018
timestamp 1677622389
transform 1 0 2348 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7028
timestamp 1677622389
transform 1 0 2348 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6987
timestamp 1677622389
transform 1 0 2364 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8125
timestamp 1677622389
transform 1 0 2356 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7123
timestamp 1677622389
transform 1 0 2356 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8080
timestamp 1677622389
transform 1 0 2452 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6988
timestamp 1677622389
transform 1 0 2484 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7967
timestamp 1677622389
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8081
timestamp 1677622389
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6972
timestamp 1677622389
transform 1 0 2516 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7968
timestamp 1677622389
transform 1 0 2532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7969
timestamp 1677622389
transform 1 0 2540 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7056
timestamp 1677622389
transform 1 0 2540 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7094
timestamp 1677622389
transform 1 0 2532 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7970
timestamp 1677622389
transform 1 0 2588 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7057
timestamp 1677622389
transform 1 0 2588 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7149
timestamp 1677622389
transform 1 0 2556 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7971
timestamp 1677622389
transform 1 0 2612 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7150
timestamp 1677622389
transform 1 0 2612 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7972
timestamp 1677622389
transform 1 0 2644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8082
timestamp 1677622389
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7058
timestamp 1677622389
transform 1 0 2644 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_6973
timestamp 1677622389
transform 1 0 2716 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6974
timestamp 1677622389
transform 1 0 2740 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6989
timestamp 1677622389
transform 1 0 2716 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7973
timestamp 1677622389
transform 1 0 2740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8083
timestamp 1677622389
transform 1 0 2652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8084
timestamp 1677622389
transform 1 0 2660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8085
timestamp 1677622389
transform 1 0 2716 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7095
timestamp 1677622389
transform 1 0 2636 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7096
timestamp 1677622389
transform 1 0 2652 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7124
timestamp 1677622389
transform 1 0 2660 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8086
timestamp 1677622389
transform 1 0 2756 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7097
timestamp 1677622389
transform 1 0 2756 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_6975
timestamp 1677622389
transform 1 0 2796 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6976
timestamp 1677622389
transform 1 0 2844 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6977
timestamp 1677622389
transform 1 0 2868 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_6990
timestamp 1677622389
transform 1 0 2820 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7029
timestamp 1677622389
transform 1 0 2828 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7974
timestamp 1677622389
transform 1 0 2852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8087
timestamp 1677622389
transform 1 0 2828 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7098
timestamp 1677622389
transform 1 0 2820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_6991
timestamp 1677622389
transform 1 0 2884 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7912
timestamp 1677622389
transform 1 0 2884 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7975
timestamp 1677622389
transform 1 0 2876 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7030
timestamp 1677622389
transform 1 0 2980 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6992
timestamp 1677622389
transform 1 0 2996 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7976
timestamp 1677622389
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7977
timestamp 1677622389
transform 1 0 2996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8088
timestamp 1677622389
transform 1 0 2972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8089
timestamp 1677622389
transform 1 0 2980 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7099
timestamp 1677622389
transform 1 0 2980 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8126
timestamp 1677622389
transform 1 0 3052 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8127
timestamp 1677622389
transform 1 0 3084 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7125
timestamp 1677622389
transform 1 0 3084 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7059
timestamp 1677622389
transform 1 0 3108 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8090
timestamp 1677622389
transform 1 0 3116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8145
timestamp 1677622389
transform 1 0 3100 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_8128
timestamp 1677622389
transform 1 0 3140 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7151
timestamp 1677622389
transform 1 0 3140 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7913
timestamp 1677622389
transform 1 0 3156 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7060
timestamp 1677622389
transform 1 0 3148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7152
timestamp 1677622389
transform 1 0 3156 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7978
timestamp 1677622389
transform 1 0 3180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8091
timestamp 1677622389
transform 1 0 3180 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7031
timestamp 1677622389
transform 1 0 3220 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7979
timestamp 1677622389
transform 1 0 3236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8092
timestamp 1677622389
transform 1 0 3220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8093
timestamp 1677622389
transform 1 0 3228 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6993
timestamp 1677622389
transform 1 0 3252 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7100
timestamp 1677622389
transform 1 0 3252 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7019
timestamp 1677622389
transform 1 0 3276 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7980
timestamp 1677622389
transform 1 0 3300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7981
timestamp 1677622389
transform 1 0 3308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8094
timestamp 1677622389
transform 1 0 3276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8095
timestamp 1677622389
transform 1 0 3292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8096
timestamp 1677622389
transform 1 0 3316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8097
timestamp 1677622389
transform 1 0 3324 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7164
timestamp 1677622389
transform 1 0 3316 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7982
timestamp 1677622389
transform 1 0 3340 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7153
timestamp 1677622389
transform 1 0 3332 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7983
timestamp 1677622389
transform 1 0 3356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7984
timestamp 1677622389
transform 1 0 3372 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7061
timestamp 1677622389
transform 1 0 3348 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8098
timestamp 1677622389
transform 1 0 3364 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7062
timestamp 1677622389
transform 1 0 3372 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7101
timestamp 1677622389
transform 1 0 3356 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7126
timestamp 1677622389
transform 1 0 3364 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7154
timestamp 1677622389
transform 1 0 3356 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7155
timestamp 1677622389
transform 1 0 3372 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_6978
timestamp 1677622389
transform 1 0 3396 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7156
timestamp 1677622389
transform 1 0 3412 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7032
timestamp 1677622389
transform 1 0 3460 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6994
timestamp 1677622389
transform 1 0 3476 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7020
timestamp 1677622389
transform 1 0 3484 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7985
timestamp 1677622389
transform 1 0 3476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7986
timestamp 1677622389
transform 1 0 3484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8099
timestamp 1677622389
transform 1 0 3460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8100
timestamp 1677622389
transform 1 0 3468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7102
timestamp 1677622389
transform 1 0 3468 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7165
timestamp 1677622389
transform 1 0 3476 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_6995
timestamp 1677622389
transform 1 0 3492 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8101
timestamp 1677622389
transform 1 0 3492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7033
timestamp 1677622389
transform 1 0 3500 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6996
timestamp 1677622389
transform 1 0 3540 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7987
timestamp 1677622389
transform 1 0 3508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7988
timestamp 1677622389
transform 1 0 3524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8102
timestamp 1677622389
transform 1 0 3532 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7103
timestamp 1677622389
transform 1 0 3524 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8103
timestamp 1677622389
transform 1 0 3572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8129
timestamp 1677622389
transform 1 0 3564 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7989
timestamp 1677622389
transform 1 0 3580 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7127
timestamp 1677622389
transform 1 0 3572 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7157
timestamp 1677622389
transform 1 0 3564 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7034
timestamp 1677622389
transform 1 0 3588 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7990
timestamp 1677622389
transform 1 0 3604 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7035
timestamp 1677622389
transform 1 0 3612 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8104
timestamp 1677622389
transform 1 0 3596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8105
timestamp 1677622389
transform 1 0 3620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7104
timestamp 1677622389
transform 1 0 3604 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8130
timestamp 1677622389
transform 1 0 3612 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7128
timestamp 1677622389
transform 1 0 3612 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7991
timestamp 1677622389
transform 1 0 3644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8131
timestamp 1677622389
transform 1 0 3636 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7158
timestamp 1677622389
transform 1 0 3636 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7992
timestamp 1677622389
transform 1 0 3652 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7036
timestamp 1677622389
transform 1 0 3660 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8106
timestamp 1677622389
transform 1 0 3668 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7105
timestamp 1677622389
transform 1 0 3668 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_6997
timestamp 1677622389
transform 1 0 3692 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7037
timestamp 1677622389
transform 1 0 3684 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7993
timestamp 1677622389
transform 1 0 3692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8132
timestamp 1677622389
transform 1 0 3684 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8107
timestamp 1677622389
transform 1 0 3700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_6998
timestamp 1677622389
transform 1 0 3764 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7021
timestamp 1677622389
transform 1 0 3756 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7994
timestamp 1677622389
transform 1 0 3756 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7159
timestamp 1677622389
transform 1 0 3748 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7995
timestamp 1677622389
transform 1 0 3780 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_6979
timestamp 1677622389
transform 1 0 3812 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8108
timestamp 1677622389
transform 1 0 3796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8109
timestamp 1677622389
transform 1 0 3812 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7129
timestamp 1677622389
transform 1 0 3788 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7160
timestamp 1677622389
transform 1 0 3788 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7130
timestamp 1677622389
transform 1 0 3812 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7996
timestamp 1677622389
transform 1 0 3836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7997
timestamp 1677622389
transform 1 0 3860 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7063
timestamp 1677622389
transform 1 0 3860 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8133
timestamp 1677622389
transform 1 0 3852 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7131
timestamp 1677622389
transform 1 0 3852 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7064
timestamp 1677622389
transform 1 0 3892 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8134
timestamp 1677622389
transform 1 0 3892 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7132
timestamp 1677622389
transform 1 0 3884 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7998
timestamp 1677622389
transform 1 0 3924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8110
timestamp 1677622389
transform 1 0 3916 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7106
timestamp 1677622389
transform 1 0 3932 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7065
timestamp 1677622389
transform 1 0 3956 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8135
timestamp 1677622389
transform 1 0 3956 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7133
timestamp 1677622389
transform 1 0 3940 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8111
timestamp 1677622389
transform 1 0 3972 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7066
timestamp 1677622389
transform 1 0 4028 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8136
timestamp 1677622389
transform 1 0 4028 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7999
timestamp 1677622389
transform 1 0 4060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8000
timestamp 1677622389
transform 1 0 4068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8001
timestamp 1677622389
transform 1 0 4092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8112
timestamp 1677622389
transform 1 0 4084 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7134
timestamp 1677622389
transform 1 0 4068 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8113
timestamp 1677622389
transform 1 0 4100 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7166
timestamp 1677622389
transform 1 0 4100 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_6999
timestamp 1677622389
transform 1 0 4132 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8002
timestamp 1677622389
transform 1 0 4132 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7135
timestamp 1677622389
transform 1 0 4124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7067
timestamp 1677622389
transform 1 0 4148 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8114
timestamp 1677622389
transform 1 0 4172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8137
timestamp 1677622389
transform 1 0 4156 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7000
timestamp 1677622389
transform 1 0 4188 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8003
timestamp 1677622389
transform 1 0 4188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8115
timestamp 1677622389
transform 1 0 4204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8004
timestamp 1677622389
transform 1 0 4244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8005
timestamp 1677622389
transform 1 0 4252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8116
timestamp 1677622389
transform 1 0 4236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8138
timestamp 1677622389
transform 1 0 4220 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7136
timestamp 1677622389
transform 1 0 4220 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7068
timestamp 1677622389
transform 1 0 4252 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8006
timestamp 1677622389
transform 1 0 4332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8007
timestamp 1677622389
transform 1 0 4340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8117
timestamp 1677622389
transform 1 0 4324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8139
timestamp 1677622389
transform 1 0 4308 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7107
timestamp 1677622389
transform 1 0 4340 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8140
timestamp 1677622389
transform 1 0 4356 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7137
timestamp 1677622389
transform 1 0 4356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7069
timestamp 1677622389
transform 1 0 4396 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8141
timestamp 1677622389
transform 1 0 4412 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7138
timestamp 1677622389
transform 1 0 4412 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8008
timestamp 1677622389
transform 1 0 4436 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7070
timestamp 1677622389
transform 1 0 4436 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7022
timestamp 1677622389
transform 1 0 4452 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8009
timestamp 1677622389
transform 1 0 4452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8142
timestamp 1677622389
transform 1 0 4452 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7139
timestamp 1677622389
transform 1 0 4452 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7038
timestamp 1677622389
transform 1 0 4468 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8118
timestamp 1677622389
transform 1 0 4468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7039
timestamp 1677622389
transform 1 0 4492 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8143
timestamp 1677622389
transform 1 0 4476 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8010
timestamp 1677622389
transform 1 0 4516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8119
timestamp 1677622389
transform 1 0 4556 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7108
timestamp 1677622389
transform 1 0 4668 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8012
timestamp 1677622389
transform 1 0 4692 0 1 933
box -2 -2 2 2
use M2_M1  M2_M1_8011
timestamp 1677622389
transform 1 0 4788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8120
timestamp 1677622389
transform 1 0 4716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8121
timestamp 1677622389
transform 1 0 4772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8122
timestamp 1677622389
transform 1 0 4780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7109
timestamp 1677622389
transform 1 0 4716 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7140
timestamp 1677622389
transform 1 0 4716 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7141
timestamp 1677622389
transform 1 0 4740 0 1 905
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_76
timestamp 1677622389
transform 1 0 24 0 1 870
box -10 -3 10 3
use FILL  FILL_8906
timestamp 1677622389
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_8907
timestamp 1677622389
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_8908
timestamp 1677622389
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_8909
timestamp 1677622389
transform 1 0 96 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_563
timestamp 1677622389
transform 1 0 104 0 -1 970
box -9 -3 26 105
use FILL  FILL_8910
timestamp 1677622389
transform 1 0 120 0 -1 970
box -8 -3 16 105
use FILL  FILL_8911
timestamp 1677622389
transform 1 0 128 0 -1 970
box -8 -3 16 105
use FILL  FILL_8913
timestamp 1677622389
transform 1 0 136 0 -1 970
box -8 -3 16 105
use FILL  FILL_8915
timestamp 1677622389
transform 1 0 144 0 -1 970
box -8 -3 16 105
use FILL  FILL_8931
timestamp 1677622389
transform 1 0 152 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_565
timestamp 1677622389
transform 1 0 160 0 -1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_487
timestamp 1677622389
transform 1 0 176 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_566
timestamp 1677622389
transform -1 0 288 0 -1 970
box -9 -3 26 105
use FILL  FILL_8932
timestamp 1677622389
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_8933
timestamp 1677622389
transform 1 0 296 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_329
timestamp 1677622389
transform -1 0 344 0 -1 970
box -8 -3 46 105
use FILL  FILL_8934
timestamp 1677622389
transform 1 0 344 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_339
timestamp 1677622389
transform 1 0 352 0 -1 970
box -8 -3 46 105
use FILL  FILL_8935
timestamp 1677622389
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_8936
timestamp 1677622389
transform 1 0 400 0 -1 970
box -8 -3 16 105
use FILL  FILL_8937
timestamp 1677622389
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_8938
timestamp 1677622389
transform 1 0 416 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_567
timestamp 1677622389
transform -1 0 440 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_568
timestamp 1677622389
transform -1 0 456 0 -1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_330
timestamp 1677622389
transform 1 0 456 0 -1 970
box -8 -3 46 105
use FILL  FILL_8939
timestamp 1677622389
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_8942
timestamp 1677622389
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_8943
timestamp 1677622389
transform 1 0 512 0 -1 970
box -8 -3 16 105
use FILL  FILL_8944
timestamp 1677622389
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_8945
timestamp 1677622389
transform 1 0 528 0 -1 970
box -8 -3 16 105
use FILL  FILL_8946
timestamp 1677622389
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_8947
timestamp 1677622389
transform 1 0 544 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_569
timestamp 1677622389
transform -1 0 568 0 -1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_331
timestamp 1677622389
transform 1 0 568 0 -1 970
box -8 -3 46 105
use FILL  FILL_8948
timestamp 1677622389
transform 1 0 608 0 -1 970
box -8 -3 16 105
use FILL  FILL_8949
timestamp 1677622389
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_8950
timestamp 1677622389
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_8951
timestamp 1677622389
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_8953
timestamp 1677622389
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_8955
timestamp 1677622389
transform 1 0 648 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_490
timestamp 1677622389
transform 1 0 656 0 -1 970
box -8 -3 104 105
use FILL  FILL_8965
timestamp 1677622389
transform 1 0 752 0 -1 970
box -8 -3 16 105
use FILL  FILL_8966
timestamp 1677622389
transform 1 0 760 0 -1 970
box -8 -3 16 105
use FILL  FILL_8967
timestamp 1677622389
transform 1 0 768 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_341
timestamp 1677622389
transform 1 0 776 0 -1 970
box -8 -3 46 105
use FILL  FILL_8968
timestamp 1677622389
transform 1 0 816 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_332
timestamp 1677622389
transform 1 0 824 0 -1 970
box -8 -3 46 105
use FILL  FILL_8969
timestamp 1677622389
transform 1 0 864 0 -1 970
box -8 -3 16 105
use FILL  FILL_8970
timestamp 1677622389
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_8973
timestamp 1677622389
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_8974
timestamp 1677622389
transform 1 0 888 0 -1 970
box -8 -3 16 105
use FILL  FILL_8975
timestamp 1677622389
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_8976
timestamp 1677622389
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_8977
timestamp 1677622389
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_8978
timestamp 1677622389
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_8979
timestamp 1677622389
transform 1 0 928 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_491
timestamp 1677622389
transform 1 0 936 0 -1 970
box -8 -3 104 105
use FILL  FILL_8990
timestamp 1677622389
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_8992
timestamp 1677622389
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use FILL  FILL_8997
timestamp 1677622389
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_571
timestamp 1677622389
transform -1 0 1072 0 -1 970
box -9 -3 26 105
use FILL  FILL_8998
timestamp 1677622389
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_9000
timestamp 1677622389
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_9002
timestamp 1677622389
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_9004
timestamp 1677622389
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_9006
timestamp 1677622389
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_9008
timestamp 1677622389
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7167
timestamp 1677622389
transform 1 0 1132 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_334
timestamp 1677622389
transform 1 0 1120 0 -1 970
box -8 -3 46 105
use FILL  FILL_9012
timestamp 1677622389
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7168
timestamp 1677622389
transform 1 0 1180 0 1 875
box -3 -3 3 3
use FILL  FILL_9014
timestamp 1677622389
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_9016
timestamp 1677622389
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_9018
timestamp 1677622389
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9022
timestamp 1677622389
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9023
timestamp 1677622389
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7169
timestamp 1677622389
transform 1 0 1228 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7170
timestamp 1677622389
transform 1 0 1252 0 1 875
box -3 -3 3 3
use OAI22X1  OAI22X1_343
timestamp 1677622389
transform -1 0 1248 0 -1 970
box -8 -3 46 105
use FILL  FILL_9024
timestamp 1677622389
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_9026
timestamp 1677622389
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9045
timestamp 1677622389
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_492
timestamp 1677622389
transform -1 0 1368 0 -1 970
box -8 -3 104 105
use FILL  FILL_9046
timestamp 1677622389
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_9047
timestamp 1677622389
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7171
timestamp 1677622389
transform 1 0 1396 0 1 875
box -3 -3 3 3
use OAI22X1  OAI22X1_344
timestamp 1677622389
transform -1 0 1424 0 -1 970
box -8 -3 46 105
use FILL  FILL_9048
timestamp 1677622389
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use FILL  FILL_9049
timestamp 1677622389
transform 1 0 1432 0 -1 970
box -8 -3 16 105
use FILL  FILL_9050
timestamp 1677622389
transform 1 0 1440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9051
timestamp 1677622389
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9052
timestamp 1677622389
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_9060
timestamp 1677622389
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_336
timestamp 1677622389
transform -1 0 1512 0 -1 970
box -8 -3 46 105
use FILL  FILL_9061
timestamp 1677622389
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9062
timestamp 1677622389
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9063
timestamp 1677622389
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9065
timestamp 1677622389
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_9067
timestamp 1677622389
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_493
timestamp 1677622389
transform 1 0 1552 0 -1 970
box -8 -3 104 105
use FILL  FILL_9079
timestamp 1677622389
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use FILL  FILL_9080
timestamp 1677622389
transform 1 0 1656 0 -1 970
box -8 -3 16 105
use FILL  FILL_9081
timestamp 1677622389
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7172
timestamp 1677622389
transform 1 0 1700 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_337
timestamp 1677622389
transform 1 0 1672 0 -1 970
box -8 -3 46 105
use FILL  FILL_9082
timestamp 1677622389
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_9084
timestamp 1677622389
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_9105
timestamp 1677622389
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_577
timestamp 1677622389
transform -1 0 1752 0 -1 970
box -9 -3 26 105
use FILL  FILL_9106
timestamp 1677622389
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_340
timestamp 1677622389
transform 1 0 1760 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_495
timestamp 1677622389
transform -1 0 1896 0 -1 970
box -8 -3 104 105
use FILL  FILL_9107
timestamp 1677622389
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_9108
timestamp 1677622389
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use FILL  FILL_9109
timestamp 1677622389
transform 1 0 1912 0 -1 970
box -8 -3 16 105
use FILL  FILL_9110
timestamp 1677622389
transform 1 0 1920 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_578
timestamp 1677622389
transform 1 0 1928 0 -1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_496
timestamp 1677622389
transform 1 0 1944 0 -1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_341
timestamp 1677622389
transform -1 0 2080 0 -1 970
box -8 -3 46 105
use FILL  FILL_9111
timestamp 1677622389
transform 1 0 2080 0 -1 970
box -8 -3 16 105
use FILL  FILL_9112
timestamp 1677622389
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_68
timestamp 1677622389
transform -1 0 2128 0 -1 970
box -8 -3 40 105
use FILL  FILL_9113
timestamp 1677622389
transform 1 0 2128 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7173
timestamp 1677622389
transform 1 0 2148 0 1 875
box -3 -3 3 3
use FILL  FILL_9115
timestamp 1677622389
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_9117
timestamp 1677622389
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_9119
timestamp 1677622389
transform 1 0 2152 0 -1 970
box -8 -3 16 105
use FILL  FILL_9122
timestamp 1677622389
transform 1 0 2160 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_580
timestamp 1677622389
transform 1 0 2168 0 -1 970
box -9 -3 26 105
use FILL  FILL_9123
timestamp 1677622389
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9125
timestamp 1677622389
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7174
timestamp 1677622389
transform 1 0 2220 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_497
timestamp 1677622389
transform 1 0 2200 0 -1 970
box -8 -3 104 105
use FILL  FILL_9136
timestamp 1677622389
transform 1 0 2296 0 -1 970
box -8 -3 16 105
use FILL  FILL_9137
timestamp 1677622389
transform 1 0 2304 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_22
timestamp 1677622389
transform 1 0 2312 0 -1 970
box -8 -3 32 105
use FILL  FILL_9138
timestamp 1677622389
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use FILL  FILL_9139
timestamp 1677622389
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use FILL  FILL_9140
timestamp 1677622389
transform 1 0 2352 0 -1 970
box -8 -3 16 105
use FILL  FILL_9141
timestamp 1677622389
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_9142
timestamp 1677622389
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_9143
timestamp 1677622389
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_9144
timestamp 1677622389
transform 1 0 2384 0 -1 970
box -8 -3 16 105
use FILL  FILL_9145
timestamp 1677622389
transform 1 0 2392 0 -1 970
box -8 -3 16 105
use FILL  FILL_9146
timestamp 1677622389
transform 1 0 2400 0 -1 970
box -8 -3 16 105
use FILL  FILL_9147
timestamp 1677622389
transform 1 0 2408 0 -1 970
box -8 -3 16 105
use FILL  FILL_9148
timestamp 1677622389
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use FILL  FILL_9150
timestamp 1677622389
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_9152
timestamp 1677622389
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_9156
timestamp 1677622389
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9157
timestamp 1677622389
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_14
timestamp 1677622389
transform 1 0 2456 0 -1 970
box -7 -3 39 105
use FILL  FILL_9158
timestamp 1677622389
transform 1 0 2488 0 -1 970
box -8 -3 16 105
use FILL  FILL_9160
timestamp 1677622389
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use FILL  FILL_9162
timestamp 1677622389
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_9164
timestamp 1677622389
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_583
timestamp 1677622389
transform -1 0 2536 0 -1 970
box -9 -3 26 105
use XOR2X1  XOR2X1_3
timestamp 1677622389
transform 1 0 2536 0 -1 970
box -8 -3 64 105
use FILL  FILL_9165
timestamp 1677622389
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_9166
timestamp 1677622389
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_9168
timestamp 1677622389
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_343
timestamp 1677622389
transform 1 0 2616 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_499
timestamp 1677622389
transform -1 0 2752 0 -1 970
box -8 -3 104 105
use FILL  FILL_9183
timestamp 1677622389
transform 1 0 2752 0 -1 970
box -8 -3 16 105
use FILL  FILL_9184
timestamp 1677622389
transform 1 0 2760 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_500
timestamp 1677622389
transform -1 0 2864 0 -1 970
box -8 -3 104 105
use FILL  FILL_9185
timestamp 1677622389
transform 1 0 2864 0 -1 970
box -8 -3 16 105
use FAX1  FAX1_17
timestamp 1677622389
transform -1 0 2992 0 -1 970
box -5 -3 126 105
use FILL  FILL_9186
timestamp 1677622389
transform 1 0 2992 0 -1 970
box -8 -3 16 105
use FILL  FILL_9188
timestamp 1677622389
transform 1 0 3000 0 -1 970
box -8 -3 16 105
use FILL  FILL_9191
timestamp 1677622389
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_25
timestamp 1677622389
transform 1 0 3016 0 -1 970
box -8 -3 32 105
use FILL  FILL_9192
timestamp 1677622389
transform 1 0 3040 0 -1 970
box -8 -3 16 105
use FILL  FILL_9193
timestamp 1677622389
transform 1 0 3048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9194
timestamp 1677622389
transform 1 0 3056 0 -1 970
box -8 -3 16 105
use FILL  FILL_9195
timestamp 1677622389
transform 1 0 3064 0 -1 970
box -8 -3 16 105
use FILL  FILL_9197
timestamp 1677622389
transform 1 0 3072 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1677622389
transform 1 0 3080 0 -1 970
box -8 -3 40 105
use FILL  FILL_9199
timestamp 1677622389
transform 1 0 3112 0 -1 970
box -8 -3 16 105
use FILL  FILL_9201
timestamp 1677622389
transform 1 0 3120 0 -1 970
box -8 -3 16 105
use FILL  FILL_9203
timestamp 1677622389
transform 1 0 3128 0 -1 970
box -8 -3 16 105
use FILL  FILL_9205
timestamp 1677622389
transform 1 0 3136 0 -1 970
box -8 -3 16 105
use FILL  FILL_9209
timestamp 1677622389
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_15
timestamp 1677622389
transform -1 0 3184 0 -1 970
box -7 -3 39 105
use FILL  FILL_9210
timestamp 1677622389
transform 1 0 3184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9211
timestamp 1677622389
transform 1 0 3192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9214
timestamp 1677622389
transform 1 0 3200 0 -1 970
box -8 -3 16 105
use FILL  FILL_9215
timestamp 1677622389
transform 1 0 3208 0 -1 970
box -8 -3 16 105
use FILL  FILL_9216
timestamp 1677622389
transform 1 0 3216 0 -1 970
box -8 -3 16 105
use FILL  FILL_9217
timestamp 1677622389
transform 1 0 3224 0 -1 970
box -8 -3 16 105
use FILL  FILL_9219
timestamp 1677622389
transform 1 0 3232 0 -1 970
box -8 -3 16 105
use FILL  FILL_9221
timestamp 1677622389
transform 1 0 3240 0 -1 970
box -8 -3 16 105
use FILL  FILL_9223
timestamp 1677622389
transform 1 0 3248 0 -1 970
box -8 -3 16 105
use FILL  FILL_9227
timestamp 1677622389
transform 1 0 3256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9228
timestamp 1677622389
transform 1 0 3264 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_345
timestamp 1677622389
transform -1 0 3312 0 -1 970
box -8 -3 46 105
use FILL  FILL_9229
timestamp 1677622389
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use FILL  FILL_9231
timestamp 1677622389
transform 1 0 3320 0 -1 970
box -8 -3 16 105
use FILL  FILL_9233
timestamp 1677622389
transform 1 0 3328 0 -1 970
box -8 -3 16 105
use FILL  FILL_9235
timestamp 1677622389
transform 1 0 3336 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_346
timestamp 1677622389
transform 1 0 3344 0 -1 970
box -8 -3 46 105
use FILL  FILL_9242
timestamp 1677622389
transform 1 0 3384 0 -1 970
box -8 -3 16 105
use FILL  FILL_9245
timestamp 1677622389
transform 1 0 3392 0 -1 970
box -8 -3 16 105
use FILL  FILL_9246
timestamp 1677622389
transform 1 0 3400 0 -1 970
box -8 -3 16 105
use FILL  FILL_9247
timestamp 1677622389
transform 1 0 3408 0 -1 970
box -8 -3 16 105
use FILL  FILL_9248
timestamp 1677622389
transform 1 0 3416 0 -1 970
box -8 -3 16 105
use FILL  FILL_9249
timestamp 1677622389
transform 1 0 3424 0 -1 970
box -8 -3 16 105
use FILL  FILL_9250
timestamp 1677622389
transform 1 0 3432 0 -1 970
box -8 -3 16 105
use FILL  FILL_9251
timestamp 1677622389
transform 1 0 3440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9252
timestamp 1677622389
transform 1 0 3448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9253
timestamp 1677622389
transform 1 0 3456 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_586
timestamp 1677622389
transform -1 0 3480 0 -1 970
box -9 -3 26 105
use FILL  FILL_9254
timestamp 1677622389
transform 1 0 3480 0 -1 970
box -8 -3 16 105
use FILL  FILL_9255
timestamp 1677622389
transform 1 0 3488 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7175
timestamp 1677622389
transform 1 0 3508 0 1 875
box -3 -3 3 3
use FILL  FILL_9256
timestamp 1677622389
transform 1 0 3496 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_587
timestamp 1677622389
transform 1 0 3504 0 -1 970
box -9 -3 26 105
use AND2X2  AND2X2_55
timestamp 1677622389
transform 1 0 3520 0 -1 970
box -8 -3 40 105
use FILL  FILL_9257
timestamp 1677622389
transform 1 0 3552 0 -1 970
box -8 -3 16 105
use FILL  FILL_9259
timestamp 1677622389
transform 1 0 3560 0 -1 970
box -8 -3 16 105
use FILL  FILL_9269
timestamp 1677622389
transform 1 0 3568 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_156
timestamp 1677622389
transform -1 0 3608 0 -1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_26
timestamp 1677622389
transform -1 0 3632 0 -1 970
box -8 -3 32 105
use FILL  FILL_9270
timestamp 1677622389
transform 1 0 3632 0 -1 970
box -8 -3 16 105
use FILL  FILL_9274
timestamp 1677622389
transform 1 0 3640 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_157
timestamp 1677622389
transform -1 0 3680 0 -1 970
box -8 -3 34 105
use FILL  FILL_9275
timestamp 1677622389
transform 1 0 3680 0 -1 970
box -8 -3 16 105
use FILL  FILL_9276
timestamp 1677622389
transform 1 0 3688 0 -1 970
box -8 -3 16 105
use FILL  FILL_9277
timestamp 1677622389
transform 1 0 3696 0 -1 970
box -8 -3 16 105
use FILL  FILL_9279
timestamp 1677622389
transform 1 0 3704 0 -1 970
box -8 -3 16 105
use FILL  FILL_9285
timestamp 1677622389
transform 1 0 3712 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_27
timestamp 1677622389
transform -1 0 3744 0 -1 970
box -8 -3 32 105
use FILL  FILL_9286
timestamp 1677622389
transform 1 0 3744 0 -1 970
box -8 -3 16 105
use FILL  FILL_9288
timestamp 1677622389
transform 1 0 3752 0 -1 970
box -8 -3 16 105
use FILL  FILL_9290
timestamp 1677622389
transform 1 0 3760 0 -1 970
box -8 -3 16 105
use FILL  FILL_9292
timestamp 1677622389
transform 1 0 3768 0 -1 970
box -8 -3 16 105
use FILL  FILL_9294
timestamp 1677622389
transform 1 0 3776 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_158
timestamp 1677622389
transform 1 0 3784 0 -1 970
box -8 -3 34 105
use FILL  FILL_9296
timestamp 1677622389
transform 1 0 3816 0 -1 970
box -8 -3 16 105
use FILL  FILL_9297
timestamp 1677622389
transform 1 0 3824 0 -1 970
box -8 -3 16 105
use FILL  FILL_9302
timestamp 1677622389
transform 1 0 3832 0 -1 970
box -8 -3 16 105
use FILL  FILL_9303
timestamp 1677622389
transform 1 0 3840 0 -1 970
box -8 -3 16 105
use FILL  FILL_9304
timestamp 1677622389
transform 1 0 3848 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_29
timestamp 1677622389
transform 1 0 3856 0 -1 970
box -8 -3 32 105
use FILL  FILL_9305
timestamp 1677622389
transform 1 0 3880 0 -1 970
box -8 -3 16 105
use FILL  FILL_9307
timestamp 1677622389
transform 1 0 3888 0 -1 970
box -8 -3 16 105
use FILL  FILL_9312
timestamp 1677622389
transform 1 0 3896 0 -1 970
box -8 -3 16 105
use FILL  FILL_9313
timestamp 1677622389
transform 1 0 3904 0 -1 970
box -8 -3 16 105
use FILL  FILL_9314
timestamp 1677622389
transform 1 0 3912 0 -1 970
box -8 -3 16 105
use FILL  FILL_9315
timestamp 1677622389
transform 1 0 3920 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_159
timestamp 1677622389
transform 1 0 3928 0 -1 970
box -8 -3 34 105
use FILL  FILL_9316
timestamp 1677622389
transform 1 0 3960 0 -1 970
box -8 -3 16 105
use FILL  FILL_9318
timestamp 1677622389
transform 1 0 3968 0 -1 970
box -8 -3 16 105
use FILL  FILL_9321
timestamp 1677622389
transform 1 0 3976 0 -1 970
box -8 -3 16 105
use FILL  FILL_9322
timestamp 1677622389
transform 1 0 3984 0 -1 970
box -8 -3 16 105
use FILL  FILL_9323
timestamp 1677622389
transform 1 0 3992 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_30
timestamp 1677622389
transform -1 0 4024 0 -1 970
box -8 -3 32 105
use FILL  FILL_9324
timestamp 1677622389
transform 1 0 4024 0 -1 970
box -8 -3 16 105
use FILL  FILL_9326
timestamp 1677622389
transform 1 0 4032 0 -1 970
box -8 -3 16 105
use FILL  FILL_9328
timestamp 1677622389
transform 1 0 4040 0 -1 970
box -8 -3 16 105
use FILL  FILL_9330
timestamp 1677622389
transform 1 0 4048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9333
timestamp 1677622389
transform 1 0 4056 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_160
timestamp 1677622389
transform -1 0 4096 0 -1 970
box -8 -3 34 105
use FILL  FILL_9334
timestamp 1677622389
transform 1 0 4096 0 -1 970
box -8 -3 16 105
use FILL  FILL_9335
timestamp 1677622389
transform 1 0 4104 0 -1 970
box -8 -3 16 105
use FILL  FILL_9337
timestamp 1677622389
transform 1 0 4112 0 -1 970
box -8 -3 16 105
use FILL  FILL_9339
timestamp 1677622389
transform 1 0 4120 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1677622389
transform 1 0 4128 0 -1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_161
timestamp 1677622389
transform -1 0 4184 0 -1 970
box -8 -3 34 105
use M3_M2  M3_M2_7176
timestamp 1677622389
transform 1 0 4196 0 1 875
box -3 -3 3 3
use FILL  FILL_9343
timestamp 1677622389
transform 1 0 4184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9345
timestamp 1677622389
transform 1 0 4192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9347
timestamp 1677622389
transform 1 0 4200 0 -1 970
box -8 -3 16 105
use FILL  FILL_9351
timestamp 1677622389
transform 1 0 4208 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_162
timestamp 1677622389
transform -1 0 4248 0 -1 970
box -8 -3 34 105
use FILL  FILL_9352
timestamp 1677622389
transform 1 0 4248 0 -1 970
box -8 -3 16 105
use FILL  FILL_9353
timestamp 1677622389
transform 1 0 4256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9354
timestamp 1677622389
transform 1 0 4264 0 -1 970
box -8 -3 16 105
use FILL  FILL_9356
timestamp 1677622389
transform 1 0 4272 0 -1 970
box -8 -3 16 105
use FILL  FILL_9358
timestamp 1677622389
transform 1 0 4280 0 -1 970
box -8 -3 16 105
use FILL  FILL_9360
timestamp 1677622389
transform 1 0 4288 0 -1 970
box -8 -3 16 105
use FILL  FILL_9367
timestamp 1677622389
transform 1 0 4296 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_163
timestamp 1677622389
transform -1 0 4336 0 -1 970
box -8 -3 34 105
use FILL  FILL_9368
timestamp 1677622389
transform 1 0 4336 0 -1 970
box -8 -3 16 105
use FILL  FILL_9370
timestamp 1677622389
transform 1 0 4344 0 -1 970
box -8 -3 16 105
use FILL  FILL_9372
timestamp 1677622389
transform 1 0 4352 0 -1 970
box -8 -3 16 105
use FILL  FILL_9375
timestamp 1677622389
transform 1 0 4360 0 -1 970
box -8 -3 16 105
use FILL  FILL_9376
timestamp 1677622389
transform 1 0 4368 0 -1 970
box -8 -3 16 105
use FILL  FILL_9377
timestamp 1677622389
transform 1 0 4376 0 -1 970
box -8 -3 16 105
use FILL  FILL_9378
timestamp 1677622389
transform 1 0 4384 0 -1 970
box -8 -3 16 105
use FILL  FILL_9379
timestamp 1677622389
transform 1 0 4392 0 -1 970
box -8 -3 16 105
use FILL  FILL_9380
timestamp 1677622389
transform 1 0 4400 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_166
timestamp 1677622389
transform -1 0 4440 0 -1 970
box -8 -3 34 105
use FILL  FILL_9382
timestamp 1677622389
transform 1 0 4440 0 -1 970
box -8 -3 16 105
use FILL  FILL_9384
timestamp 1677622389
transform 1 0 4448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9386
timestamp 1677622389
transform 1 0 4456 0 -1 970
box -8 -3 16 105
use FILL  FILL_9393
timestamp 1677622389
transform 1 0 4464 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_167
timestamp 1677622389
transform -1 0 4504 0 -1 970
box -8 -3 34 105
use FILL  FILL_9394
timestamp 1677622389
transform 1 0 4504 0 -1 970
box -8 -3 16 105
use FILL  FILL_9397
timestamp 1677622389
transform 1 0 4512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9398
timestamp 1677622389
transform 1 0 4520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9399
timestamp 1677622389
transform 1 0 4528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9400
timestamp 1677622389
transform 1 0 4536 0 -1 970
box -8 -3 16 105
use FILL  FILL_9401
timestamp 1677622389
transform 1 0 4544 0 -1 970
box -8 -3 16 105
use FILL  FILL_9402
timestamp 1677622389
transform 1 0 4552 0 -1 970
box -8 -3 16 105
use FILL  FILL_9404
timestamp 1677622389
transform 1 0 4560 0 -1 970
box -8 -3 16 105
use FILL  FILL_9405
timestamp 1677622389
transform 1 0 4568 0 -1 970
box -8 -3 16 105
use FILL  FILL_9406
timestamp 1677622389
transform 1 0 4576 0 -1 970
box -8 -3 16 105
use FILL  FILL_9407
timestamp 1677622389
transform 1 0 4584 0 -1 970
box -8 -3 16 105
use FILL  FILL_9408
timestamp 1677622389
transform 1 0 4592 0 -1 970
box -8 -3 16 105
use FILL  FILL_9409
timestamp 1677622389
transform 1 0 4600 0 -1 970
box -8 -3 16 105
use FILL  FILL_9411
timestamp 1677622389
transform 1 0 4608 0 -1 970
box -8 -3 16 105
use FILL  FILL_9413
timestamp 1677622389
transform 1 0 4616 0 -1 970
box -8 -3 16 105
use FILL  FILL_9416
timestamp 1677622389
transform 1 0 4624 0 -1 970
box -8 -3 16 105
use FILL  FILL_9417
timestamp 1677622389
transform 1 0 4632 0 -1 970
box -8 -3 16 105
use FILL  FILL_9418
timestamp 1677622389
transform 1 0 4640 0 -1 970
box -8 -3 16 105
use FILL  FILL_9419
timestamp 1677622389
transform 1 0 4648 0 -1 970
box -8 -3 16 105
use FILL  FILL_9420
timestamp 1677622389
transform 1 0 4656 0 -1 970
box -8 -3 16 105
use FILL  FILL_9421
timestamp 1677622389
transform 1 0 4664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9423
timestamp 1677622389
transform 1 0 4672 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_502
timestamp 1677622389
transform 1 0 4680 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_588
timestamp 1677622389
transform -1 0 4792 0 -1 970
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_77
timestamp 1677622389
transform 1 0 4843 0 1 870
box -10 -3 10 3
use M2_M1  M2_M1_8157
timestamp 1677622389
transform 1 0 116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8158
timestamp 1677622389
transform 1 0 164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8273
timestamp 1677622389
transform 1 0 84 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7193
timestamp 1677622389
transform 1 0 212 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7209
timestamp 1677622389
transform 1 0 300 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7236
timestamp 1677622389
transform 1 0 204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7237
timestamp 1677622389
transform 1 0 244 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8159
timestamp 1677622389
transform 1 0 204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8160
timestamp 1677622389
transform 1 0 244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8274
timestamp 1677622389
transform 1 0 196 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7319
timestamp 1677622389
transform 1 0 196 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8275
timestamp 1677622389
transform 1 0 220 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7320
timestamp 1677622389
transform 1 0 252 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7350
timestamp 1677622389
transform 1 0 220 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7351
timestamp 1677622389
transform 1 0 260 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7238
timestamp 1677622389
transform 1 0 308 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8161
timestamp 1677622389
transform 1 0 316 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7194
timestamp 1677622389
transform 1 0 340 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7210
timestamp 1677622389
transform 1 0 332 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8162
timestamp 1677622389
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8276
timestamp 1677622389
transform 1 0 340 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7195
timestamp 1677622389
transform 1 0 436 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7196
timestamp 1677622389
transform 1 0 476 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7211
timestamp 1677622389
transform 1 0 484 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7239
timestamp 1677622389
transform 1 0 460 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8163
timestamp 1677622389
transform 1 0 460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8164
timestamp 1677622389
transform 1 0 476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8277
timestamp 1677622389
transform 1 0 468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8278
timestamp 1677622389
transform 1 0 484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8279
timestamp 1677622389
transform 1 0 492 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7352
timestamp 1677622389
transform 1 0 468 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7197
timestamp 1677622389
transform 1 0 532 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8165
timestamp 1677622389
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8166
timestamp 1677622389
transform 1 0 548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8167
timestamp 1677622389
transform 1 0 564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8280
timestamp 1677622389
transform 1 0 540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8281
timestamp 1677622389
transform 1 0 564 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7321
timestamp 1677622389
transform 1 0 564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7274
timestamp 1677622389
transform 1 0 596 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8282
timestamp 1677622389
transform 1 0 596 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7212
timestamp 1677622389
transform 1 0 612 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7240
timestamp 1677622389
transform 1 0 636 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8168
timestamp 1677622389
transform 1 0 612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8169
timestamp 1677622389
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8170
timestamp 1677622389
transform 1 0 644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8283
timestamp 1677622389
transform 1 0 620 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7296
timestamp 1677622389
transform 1 0 628 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8284
timestamp 1677622389
transform 1 0 636 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7353
timestamp 1677622389
transform 1 0 636 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7177
timestamp 1677622389
transform 1 0 700 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7213
timestamp 1677622389
transform 1 0 700 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7241
timestamp 1677622389
transform 1 0 676 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8171
timestamp 1677622389
transform 1 0 676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8172
timestamp 1677622389
transform 1 0 700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8285
timestamp 1677622389
transform 1 0 676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8286
timestamp 1677622389
transform 1 0 692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7322
timestamp 1677622389
transform 1 0 676 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8173
timestamp 1677622389
transform 1 0 716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8287
timestamp 1677622389
transform 1 0 716 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7323
timestamp 1677622389
transform 1 0 716 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7242
timestamp 1677622389
transform 1 0 740 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7214
timestamp 1677622389
transform 1 0 772 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7275
timestamp 1677622389
transform 1 0 748 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8174
timestamp 1677622389
transform 1 0 756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8175
timestamp 1677622389
transform 1 0 772 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7198
timestamp 1677622389
transform 1 0 828 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7215
timestamp 1677622389
transform 1 0 804 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7243
timestamp 1677622389
transform 1 0 812 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8176
timestamp 1677622389
transform 1 0 796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8177
timestamp 1677622389
transform 1 0 812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8178
timestamp 1677622389
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8288
timestamp 1677622389
transform 1 0 740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8289
timestamp 1677622389
transform 1 0 748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8290
timestamp 1677622389
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8291
timestamp 1677622389
transform 1 0 780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8292
timestamp 1677622389
transform 1 0 788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8293
timestamp 1677622389
transform 1 0 820 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7324
timestamp 1677622389
transform 1 0 788 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7354
timestamp 1677622389
transform 1 0 764 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8179
timestamp 1677622389
transform 1 0 844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8294
timestamp 1677622389
transform 1 0 836 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7244
timestamp 1677622389
transform 1 0 868 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7245
timestamp 1677622389
transform 1 0 916 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8180
timestamp 1677622389
transform 1 0 868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8181
timestamp 1677622389
transform 1 0 884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8182
timestamp 1677622389
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8295
timestamp 1677622389
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8296
timestamp 1677622389
transform 1 0 980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8382
timestamp 1677622389
transform 1 0 980 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7355
timestamp 1677622389
transform 1 0 980 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7297
timestamp 1677622389
transform 1 0 1004 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8383
timestamp 1677622389
transform 1 0 1004 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_8183
timestamp 1677622389
transform 1 0 1044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8297
timestamp 1677622389
transform 1 0 1052 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7325
timestamp 1677622389
transform 1 0 1044 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7356
timestamp 1677622389
transform 1 0 1052 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8384
timestamp 1677622389
transform 1 0 1076 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_8184
timestamp 1677622389
transform 1 0 1092 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7357
timestamp 1677622389
transform 1 0 1084 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7276
timestamp 1677622389
transform 1 0 1100 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8185
timestamp 1677622389
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8298
timestamp 1677622389
transform 1 0 1108 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7298
timestamp 1677622389
transform 1 0 1116 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7182
timestamp 1677622389
transform 1 0 1164 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7199
timestamp 1677622389
transform 1 0 1220 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7216
timestamp 1677622389
transform 1 0 1180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7246
timestamp 1677622389
transform 1 0 1236 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7183
timestamp 1677622389
transform 1 0 1260 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7217
timestamp 1677622389
transform 1 0 1260 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8186
timestamp 1677622389
transform 1 0 1180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8187
timestamp 1677622389
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8188
timestamp 1677622389
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8189
timestamp 1677622389
transform 1 0 1236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8190
timestamp 1677622389
transform 1 0 1252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8191
timestamp 1677622389
transform 1 0 1260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8299
timestamp 1677622389
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7299
timestamp 1677622389
transform 1 0 1196 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8300
timestamp 1677622389
transform 1 0 1220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8301
timestamp 1677622389
transform 1 0 1244 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7358
timestamp 1677622389
transform 1 0 1244 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7218
timestamp 1677622389
transform 1 0 1276 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7247
timestamp 1677622389
transform 1 0 1284 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8192
timestamp 1677622389
transform 1 0 1292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8302
timestamp 1677622389
transform 1 0 1284 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7326
timestamp 1677622389
transform 1 0 1284 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8303
timestamp 1677622389
transform 1 0 1300 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7359
timestamp 1677622389
transform 1 0 1300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7200
timestamp 1677622389
transform 1 0 1356 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8193
timestamp 1677622389
transform 1 0 1340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8194
timestamp 1677622389
transform 1 0 1356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8195
timestamp 1677622389
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8304
timestamp 1677622389
transform 1 0 1348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8305
timestamp 1677622389
transform 1 0 1356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7184
timestamp 1677622389
transform 1 0 1420 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7201
timestamp 1677622389
transform 1 0 1444 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7248
timestamp 1677622389
transform 1 0 1452 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7185
timestamp 1677622389
transform 1 0 1500 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7202
timestamp 1677622389
transform 1 0 1524 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7249
timestamp 1677622389
transform 1 0 1532 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8196
timestamp 1677622389
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8197
timestamp 1677622389
transform 1 0 1452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8198
timestamp 1677622389
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8199
timestamp 1677622389
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8200
timestamp 1677622389
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8201
timestamp 1677622389
transform 1 0 1532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8306
timestamp 1677622389
transform 1 0 1476 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7327
timestamp 1677622389
transform 1 0 1476 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8307
timestamp 1677622389
transform 1 0 1500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8308
timestamp 1677622389
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8309
timestamp 1677622389
transform 1 0 1524 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7328
timestamp 1677622389
transform 1 0 1500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7360
timestamp 1677622389
transform 1 0 1508 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7361
timestamp 1677622389
transform 1 0 1524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7219
timestamp 1677622389
transform 1 0 1604 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8202
timestamp 1677622389
transform 1 0 1588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8203
timestamp 1677622389
transform 1 0 1604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8310
timestamp 1677622389
transform 1 0 1580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8311
timestamp 1677622389
transform 1 0 1596 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7220
timestamp 1677622389
transform 1 0 1636 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7250
timestamp 1677622389
transform 1 0 1644 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8312
timestamp 1677622389
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8313
timestamp 1677622389
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7251
timestamp 1677622389
transform 1 0 1668 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8204
timestamp 1677622389
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8205
timestamp 1677622389
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7277
timestamp 1677622389
transform 1 0 1692 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8206
timestamp 1677622389
transform 1 0 1700 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7278
timestamp 1677622389
transform 1 0 1708 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8207
timestamp 1677622389
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8314
timestamp 1677622389
transform 1 0 1676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8315
timestamp 1677622389
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7362
timestamp 1677622389
transform 1 0 1676 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7221
timestamp 1677622389
transform 1 0 1724 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8316
timestamp 1677622389
transform 1 0 1732 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7329
timestamp 1677622389
transform 1 0 1732 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8317
timestamp 1677622389
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7203
timestamp 1677622389
transform 1 0 1788 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7222
timestamp 1677622389
transform 1 0 1780 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7252
timestamp 1677622389
transform 1 0 1788 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8208
timestamp 1677622389
transform 1 0 1780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8318
timestamp 1677622389
transform 1 0 1788 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7186
timestamp 1677622389
transform 1 0 1812 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7187
timestamp 1677622389
transform 1 0 1836 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7204
timestamp 1677622389
transform 1 0 1804 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7223
timestamp 1677622389
transform 1 0 1876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7253
timestamp 1677622389
transform 1 0 1820 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7254
timestamp 1677622389
transform 1 0 1836 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7224
timestamp 1677622389
transform 1 0 1948 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7255
timestamp 1677622389
transform 1 0 1940 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8209
timestamp 1677622389
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8210
timestamp 1677622389
transform 1 0 1820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8211
timestamp 1677622389
transform 1 0 1836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8212
timestamp 1677622389
transform 1 0 1844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8213
timestamp 1677622389
transform 1 0 1876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8214
timestamp 1677622389
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8215
timestamp 1677622389
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8216
timestamp 1677622389
transform 1 0 1972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8319
timestamp 1677622389
transform 1 0 1804 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8320
timestamp 1677622389
transform 1 0 1828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8321
timestamp 1677622389
transform 1 0 1836 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7330
timestamp 1677622389
transform 1 0 1804 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7300
timestamp 1677622389
transform 1 0 1844 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8322
timestamp 1677622389
transform 1 0 1924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8323
timestamp 1677622389
transform 1 0 1940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8324
timestamp 1677622389
transform 1 0 1948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8325
timestamp 1677622389
transform 1 0 1964 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7331
timestamp 1677622389
transform 1 0 1900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7363
timestamp 1677622389
transform 1 0 1964 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8217
timestamp 1677622389
transform 1 0 2028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8326
timestamp 1677622389
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7225
timestamp 1677622389
transform 1 0 2068 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7256
timestamp 1677622389
transform 1 0 2076 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8218
timestamp 1677622389
transform 1 0 2068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8327
timestamp 1677622389
transform 1 0 2060 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7332
timestamp 1677622389
transform 1 0 2060 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7301
timestamp 1677622389
transform 1 0 2084 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7226
timestamp 1677622389
transform 1 0 2108 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8148
timestamp 1677622389
transform 1 0 2108 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8146
timestamp 1677622389
transform 1 0 2140 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_7257
timestamp 1677622389
transform 1 0 2140 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8147
timestamp 1677622389
transform 1 0 2156 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_8149
timestamp 1677622389
transform 1 0 2148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8219
timestamp 1677622389
transform 1 0 2132 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7279
timestamp 1677622389
transform 1 0 2148 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7364
timestamp 1677622389
transform 1 0 2148 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7178
timestamp 1677622389
transform 1 0 2188 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_8150
timestamp 1677622389
transform 1 0 2164 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7258
timestamp 1677622389
transform 1 0 2172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7227
timestamp 1677622389
transform 1 0 2196 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8151
timestamp 1677622389
transform 1 0 2188 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7280
timestamp 1677622389
transform 1 0 2164 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8220
timestamp 1677622389
transform 1 0 2172 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7302
timestamp 1677622389
transform 1 0 2164 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8221
timestamp 1677622389
transform 1 0 2196 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7281
timestamp 1677622389
transform 1 0 2228 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7365
timestamp 1677622389
transform 1 0 2228 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7179
timestamp 1677622389
transform 1 0 2252 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7205
timestamp 1677622389
transform 1 0 2244 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8328
timestamp 1677622389
transform 1 0 2244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8329
timestamp 1677622389
transform 1 0 2252 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7366
timestamp 1677622389
transform 1 0 2244 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7188
timestamp 1677622389
transform 1 0 2268 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7282
timestamp 1677622389
transform 1 0 2276 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8222
timestamp 1677622389
transform 1 0 2284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8330
timestamp 1677622389
transform 1 0 2292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7189
timestamp 1677622389
transform 1 0 2340 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7206
timestamp 1677622389
transform 1 0 2316 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8152
timestamp 1677622389
transform 1 0 2308 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8223
timestamp 1677622389
transform 1 0 2324 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7283
timestamp 1677622389
transform 1 0 2332 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8224
timestamp 1677622389
transform 1 0 2340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8225
timestamp 1677622389
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8226
timestamp 1677622389
transform 1 0 2356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8227
timestamp 1677622389
transform 1 0 2460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8331
timestamp 1677622389
transform 1 0 2332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7303
timestamp 1677622389
transform 1 0 2340 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7284
timestamp 1677622389
transform 1 0 2468 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8228
timestamp 1677622389
transform 1 0 2484 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7285
timestamp 1677622389
transform 1 0 2492 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8332
timestamp 1677622389
transform 1 0 2452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8333
timestamp 1677622389
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7304
timestamp 1677622389
transform 1 0 2484 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8385
timestamp 1677622389
transform 1 0 2444 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7333
timestamp 1677622389
transform 1 0 2452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7334
timestamp 1677622389
transform 1 0 2476 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7367
timestamp 1677622389
transform 1 0 2468 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7228
timestamp 1677622389
transform 1 0 2532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7259
timestamp 1677622389
transform 1 0 2540 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8229
timestamp 1677622389
transform 1 0 2532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8334
timestamp 1677622389
transform 1 0 2540 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7260
timestamp 1677622389
transform 1 0 2564 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8230
timestamp 1677622389
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8335
timestamp 1677622389
transform 1 0 2556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8336
timestamp 1677622389
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7261
timestamp 1677622389
transform 1 0 2676 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8231
timestamp 1677622389
transform 1 0 2676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8337
timestamp 1677622389
transform 1 0 2700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8338
timestamp 1677622389
transform 1 0 2716 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7368
timestamp 1677622389
transform 1 0 2716 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7229
timestamp 1677622389
transform 1 0 2732 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8232
timestamp 1677622389
transform 1 0 2732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8233
timestamp 1677622389
transform 1 0 2748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8386
timestamp 1677622389
transform 1 0 2836 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7369
timestamp 1677622389
transform 1 0 2836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7230
timestamp 1677622389
transform 1 0 2852 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8234
timestamp 1677622389
transform 1 0 2852 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7262
timestamp 1677622389
transform 1 0 2876 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8235
timestamp 1677622389
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8339
timestamp 1677622389
transform 1 0 2868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8340
timestamp 1677622389
transform 1 0 2876 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8341
timestamp 1677622389
transform 1 0 2988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8342
timestamp 1677622389
transform 1 0 2996 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7335
timestamp 1677622389
transform 1 0 2956 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8387
timestamp 1677622389
transform 1 0 2980 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7370
timestamp 1677622389
transform 1 0 2996 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7336
timestamp 1677622389
transform 1 0 3012 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8153
timestamp 1677622389
transform 1 0 3036 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7286
timestamp 1677622389
transform 1 0 3060 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7263
timestamp 1677622389
transform 1 0 3084 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7264
timestamp 1677622389
transform 1 0 3116 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8236
timestamp 1677622389
transform 1 0 3084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8343
timestamp 1677622389
transform 1 0 3068 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7287
timestamp 1677622389
transform 1 0 3092 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8237
timestamp 1677622389
transform 1 0 3100 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7288
timestamp 1677622389
transform 1 0 3108 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8238
timestamp 1677622389
transform 1 0 3124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8344
timestamp 1677622389
transform 1 0 3092 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7305
timestamp 1677622389
transform 1 0 3100 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7289
timestamp 1677622389
transform 1 0 3132 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8345
timestamp 1677622389
transform 1 0 3116 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7337
timestamp 1677622389
transform 1 0 3084 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8388
timestamp 1677622389
transform 1 0 3100 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7371
timestamp 1677622389
transform 1 0 3068 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7372
timestamp 1677622389
transform 1 0 3100 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7306
timestamp 1677622389
transform 1 0 3124 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7290
timestamp 1677622389
transform 1 0 3180 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8239
timestamp 1677622389
transform 1 0 3188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8346
timestamp 1677622389
transform 1 0 3180 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7373
timestamp 1677622389
transform 1 0 3180 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7231
timestamp 1677622389
transform 1 0 3228 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7265
timestamp 1677622389
transform 1 0 3212 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8240
timestamp 1677622389
transform 1 0 3212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8241
timestamp 1677622389
transform 1 0 3228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8242
timestamp 1677622389
transform 1 0 3244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8347
timestamp 1677622389
transform 1 0 3220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8390
timestamp 1677622389
transform 1 0 3260 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_8243
timestamp 1677622389
transform 1 0 3300 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7338
timestamp 1677622389
transform 1 0 3292 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8391
timestamp 1677622389
transform 1 0 3292 0 1 785
box -2 -2 2 2
use M3_M2  M3_M2_7266
timestamp 1677622389
transform 1 0 3316 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8348
timestamp 1677622389
transform 1 0 3308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8244
timestamp 1677622389
transform 1 0 3324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8245
timestamp 1677622389
transform 1 0 3340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8349
timestamp 1677622389
transform 1 0 3332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8350
timestamp 1677622389
transform 1 0 3348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7339
timestamp 1677622389
transform 1 0 3332 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8246
timestamp 1677622389
transform 1 0 3364 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7232
timestamp 1677622389
transform 1 0 3484 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8247
timestamp 1677622389
transform 1 0 3468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8248
timestamp 1677622389
transform 1 0 3476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8351
timestamp 1677622389
transform 1 0 3372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8352
timestamp 1677622389
transform 1 0 3484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8353
timestamp 1677622389
transform 1 0 3492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8389
timestamp 1677622389
transform 1 0 3380 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7340
timestamp 1677622389
transform 1 0 3492 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7374
timestamp 1677622389
transform 1 0 3484 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8249
timestamp 1677622389
transform 1 0 3532 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7267
timestamp 1677622389
transform 1 0 3564 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7180
timestamp 1677622389
transform 1 0 3588 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7207
timestamp 1677622389
transform 1 0 3604 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8250
timestamp 1677622389
transform 1 0 3604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8354
timestamp 1677622389
transform 1 0 3612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7190
timestamp 1677622389
transform 1 0 3636 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8355
timestamp 1677622389
transform 1 0 3628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7268
timestamp 1677622389
transform 1 0 3644 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8251
timestamp 1677622389
transform 1 0 3644 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7208
timestamp 1677622389
transform 1 0 3660 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7269
timestamp 1677622389
transform 1 0 3676 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8252
timestamp 1677622389
transform 1 0 3660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8253
timestamp 1677622389
transform 1 0 3676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8356
timestamp 1677622389
transform 1 0 3668 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7307
timestamp 1677622389
transform 1 0 3676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7308
timestamp 1677622389
transform 1 0 3692 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8357
timestamp 1677622389
transform 1 0 3708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8254
timestamp 1677622389
transform 1 0 3732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8255
timestamp 1677622389
transform 1 0 3748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8358
timestamp 1677622389
transform 1 0 3740 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7309
timestamp 1677622389
transform 1 0 3748 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8256
timestamp 1677622389
transform 1 0 3764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8359
timestamp 1677622389
transform 1 0 3756 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7341
timestamp 1677622389
transform 1 0 3740 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7375
timestamp 1677622389
transform 1 0 3740 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7376
timestamp 1677622389
transform 1 0 3780 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7310
timestamp 1677622389
transform 1 0 3804 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8360
timestamp 1677622389
transform 1 0 3852 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7342
timestamp 1677622389
transform 1 0 3852 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8154
timestamp 1677622389
transform 1 0 3884 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8257
timestamp 1677622389
transform 1 0 3900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8361
timestamp 1677622389
transform 1 0 3892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8362
timestamp 1677622389
transform 1 0 3932 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7181
timestamp 1677622389
transform 1 0 3972 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7191
timestamp 1677622389
transform 1 0 4004 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8155
timestamp 1677622389
transform 1 0 4004 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7233
timestamp 1677622389
transform 1 0 4028 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8258
timestamp 1677622389
transform 1 0 4020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8259
timestamp 1677622389
transform 1 0 4028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8363
timestamp 1677622389
transform 1 0 4028 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8156
timestamp 1677622389
transform 1 0 4076 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7192
timestamp 1677622389
transform 1 0 4156 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8260
timestamp 1677622389
transform 1 0 4164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8261
timestamp 1677622389
transform 1 0 4188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8364
timestamp 1677622389
transform 1 0 4148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8365
timestamp 1677622389
transform 1 0 4156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8366
timestamp 1677622389
transform 1 0 4180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8367
timestamp 1677622389
transform 1 0 4196 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7343
timestamp 1677622389
transform 1 0 4180 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7377
timestamp 1677622389
transform 1 0 4188 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7344
timestamp 1677622389
transform 1 0 4204 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7378
timestamp 1677622389
transform 1 0 4204 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7291
timestamp 1677622389
transform 1 0 4220 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8262
timestamp 1677622389
transform 1 0 4236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8263
timestamp 1677622389
transform 1 0 4300 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7292
timestamp 1677622389
transform 1 0 4308 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8368
timestamp 1677622389
transform 1 0 4276 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8369
timestamp 1677622389
transform 1 0 4292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7311
timestamp 1677622389
transform 1 0 4300 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8370
timestamp 1677622389
transform 1 0 4308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8371
timestamp 1677622389
transform 1 0 4316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7345
timestamp 1677622389
transform 1 0 4292 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7379
timestamp 1677622389
transform 1 0 4276 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7312
timestamp 1677622389
transform 1 0 4324 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7380
timestamp 1677622389
transform 1 0 4316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7346
timestamp 1677622389
transform 1 0 4332 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8264
timestamp 1677622389
transform 1 0 4348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8265
timestamp 1677622389
transform 1 0 4372 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7293
timestamp 1677622389
transform 1 0 4380 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7313
timestamp 1677622389
transform 1 0 4356 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8372
timestamp 1677622389
transform 1 0 4364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8373
timestamp 1677622389
transform 1 0 4380 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7314
timestamp 1677622389
transform 1 0 4404 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8374
timestamp 1677622389
transform 1 0 4444 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7234
timestamp 1677622389
transform 1 0 4500 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7270
timestamp 1677622389
transform 1 0 4484 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8266
timestamp 1677622389
transform 1 0 4484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8267
timestamp 1677622389
transform 1 0 4500 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7315
timestamp 1677622389
transform 1 0 4484 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8375
timestamp 1677622389
transform 1 0 4492 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7316
timestamp 1677622389
transform 1 0 4500 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8376
timestamp 1677622389
transform 1 0 4508 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7271
timestamp 1677622389
transform 1 0 4532 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8268
timestamp 1677622389
transform 1 0 4532 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7235
timestamp 1677622389
transform 1 0 4572 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7294
timestamp 1677622389
transform 1 0 4548 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8269
timestamp 1677622389
transform 1 0 4572 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7295
timestamp 1677622389
transform 1 0 4580 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8377
timestamp 1677622389
transform 1 0 4548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8378
timestamp 1677622389
transform 1 0 4564 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7347
timestamp 1677622389
transform 1 0 4548 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7272
timestamp 1677622389
transform 1 0 4628 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7273
timestamp 1677622389
transform 1 0 4652 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8379
timestamp 1677622389
transform 1 0 4620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8270
timestamp 1677622389
transform 1 0 4636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8271
timestamp 1677622389
transform 1 0 4652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8380
timestamp 1677622389
transform 1 0 4644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7317
timestamp 1677622389
transform 1 0 4652 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8381
timestamp 1677622389
transform 1 0 4660 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7348
timestamp 1677622389
transform 1 0 4660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7318
timestamp 1677622389
transform 1 0 4676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7349
timestamp 1677622389
transform 1 0 4676 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8272
timestamp 1677622389
transform 1 0 4772 0 1 815
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_78
timestamp 1677622389
transform 1 0 48 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_7381
timestamp 1677622389
transform 1 0 148 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_503
timestamp 1677622389
transform 1 0 72 0 1 770
box -8 -3 104 105
use FILL  FILL_9426
timestamp 1677622389
transform 1 0 168 0 1 770
box -8 -3 16 105
use FILL  FILL_9427
timestamp 1677622389
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_9428
timestamp 1677622389
transform 1 0 184 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7382
timestamp 1677622389
transform 1 0 220 0 1 775
box -3 -3 3 3
use INVX2  INVX2_589
timestamp 1677622389
transform 1 0 192 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_504
timestamp 1677622389
transform 1 0 208 0 1 770
box -8 -3 104 105
use FILL  FILL_9429
timestamp 1677622389
transform 1 0 304 0 1 770
box -8 -3 16 105
use FILL  FILL_9430
timestamp 1677622389
transform 1 0 312 0 1 770
box -8 -3 16 105
use FILL  FILL_9431
timestamp 1677622389
transform 1 0 320 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7383
timestamp 1677622389
transform 1 0 412 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_505
timestamp 1677622389
transform 1 0 328 0 1 770
box -8 -3 104 105
use FILL  FILL_9432
timestamp 1677622389
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_9442
timestamp 1677622389
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_9443
timestamp 1677622389
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_9444
timestamp 1677622389
transform 1 0 448 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_350
timestamp 1677622389
transform -1 0 496 0 1 770
box -8 -3 46 105
use FILL  FILL_9445
timestamp 1677622389
transform 1 0 496 0 1 770
box -8 -3 16 105
use FILL  FILL_9446
timestamp 1677622389
transform 1 0 504 0 1 770
box -8 -3 16 105
use FILL  FILL_9447
timestamp 1677622389
transform 1 0 512 0 1 770
box -8 -3 16 105
use FILL  FILL_9448
timestamp 1677622389
transform 1 0 520 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7384
timestamp 1677622389
transform 1 0 540 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_351
timestamp 1677622389
transform 1 0 528 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_7385
timestamp 1677622389
transform 1 0 580 0 1 775
box -3 -3 3 3
use FILL  FILL_9449
timestamp 1677622389
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_9450
timestamp 1677622389
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_9451
timestamp 1677622389
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_9452
timestamp 1677622389
transform 1 0 592 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_356
timestamp 1677622389
transform -1 0 640 0 1 770
box -8 -3 46 105
use BUFX2  BUFX2_107
timestamp 1677622389
transform 1 0 640 0 1 770
box -5 -3 28 105
use FILL  FILL_9453
timestamp 1677622389
transform 1 0 664 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7386
timestamp 1677622389
transform 1 0 692 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_357
timestamp 1677622389
transform 1 0 672 0 1 770
box -8 -3 46 105
use FILL  FILL_9454
timestamp 1677622389
transform 1 0 712 0 1 770
box -8 -3 16 105
use INVX2  INVX2_592
timestamp 1677622389
transform -1 0 736 0 1 770
box -9 -3 26 105
use FILL  FILL_9455
timestamp 1677622389
transform 1 0 736 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_358
timestamp 1677622389
transform 1 0 744 0 1 770
box -8 -3 46 105
use FILL  FILL_9456
timestamp 1677622389
transform 1 0 784 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_352
timestamp 1677622389
transform -1 0 832 0 1 770
box -8 -3 46 105
use FILL  FILL_9457
timestamp 1677622389
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_9458
timestamp 1677622389
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_9459
timestamp 1677622389
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_9475
timestamp 1677622389
transform 1 0 856 0 1 770
box -8 -3 16 105
use INVX2  INVX2_596
timestamp 1677622389
transform 1 0 864 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_509
timestamp 1677622389
transform -1 0 976 0 1 770
box -8 -3 104 105
use FILL  FILL_9477
timestamp 1677622389
transform 1 0 976 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_91
timestamp 1677622389
transform 1 0 984 0 1 770
box -8 -3 32 105
use FILL  FILL_9478
timestamp 1677622389
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_9484
timestamp 1677622389
transform 1 0 1016 0 1 770
box -8 -3 16 105
use FILL  FILL_9486
timestamp 1677622389
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_9487
timestamp 1677622389
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_9488
timestamp 1677622389
transform 1 0 1040 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7387
timestamp 1677622389
transform 1 0 1076 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_92
timestamp 1677622389
transform 1 0 1048 0 1 770
box -8 -3 32 105
use FILL  FILL_9489
timestamp 1677622389
transform 1 0 1072 0 1 770
box -8 -3 16 105
use FILL  FILL_9494
timestamp 1677622389
transform 1 0 1080 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_94
timestamp 1677622389
transform 1 0 1088 0 1 770
box -8 -3 32 105
use FILL  FILL_9495
timestamp 1677622389
transform 1 0 1112 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_511
timestamp 1677622389
transform 1 0 1120 0 1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_354
timestamp 1677622389
transform -1 0 1256 0 1 770
box -8 -3 46 105
use FILL  FILL_9496
timestamp 1677622389
transform 1 0 1256 0 1 770
box -8 -3 16 105
use FILL  FILL_9497
timestamp 1677622389
transform 1 0 1264 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7388
timestamp 1677622389
transform 1 0 1292 0 1 775
box -3 -3 3 3
use INVX2  INVX2_598
timestamp 1677622389
transform -1 0 1288 0 1 770
box -9 -3 26 105
use FILL  FILL_9498
timestamp 1677622389
transform 1 0 1288 0 1 770
box -8 -3 16 105
use FILL  FILL_9499
timestamp 1677622389
transform 1 0 1296 0 1 770
box -8 -3 16 105
use FILL  FILL_9500
timestamp 1677622389
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_9508
timestamp 1677622389
transform 1 0 1312 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_356
timestamp 1677622389
transform 1 0 1320 0 1 770
box -8 -3 46 105
use INVX2  INVX2_599
timestamp 1677622389
transform 1 0 1360 0 1 770
box -9 -3 26 105
use FILL  FILL_9510
timestamp 1677622389
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_9511
timestamp 1677622389
transform 1 0 1384 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_513
timestamp 1677622389
transform -1 0 1488 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_7389
timestamp 1677622389
transform 1 0 1516 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_357
timestamp 1677622389
transform -1 0 1528 0 1 770
box -8 -3 46 105
use FILL  FILL_9512
timestamp 1677622389
transform 1 0 1528 0 1 770
box -8 -3 16 105
use INVX2  INVX2_600
timestamp 1677622389
transform 1 0 1536 0 1 770
box -9 -3 26 105
use FILL  FILL_9513
timestamp 1677622389
transform 1 0 1552 0 1 770
box -8 -3 16 105
use FILL  FILL_9514
timestamp 1677622389
transform 1 0 1560 0 1 770
box -8 -3 16 105
use FILL  FILL_9515
timestamp 1677622389
transform 1 0 1568 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_360
timestamp 1677622389
transform 1 0 1576 0 1 770
box -8 -3 46 105
use FILL  FILL_9516
timestamp 1677622389
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_9517
timestamp 1677622389
transform 1 0 1624 0 1 770
box -8 -3 16 105
use FILL  FILL_9518
timestamp 1677622389
transform 1 0 1632 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_109
timestamp 1677622389
transform -1 0 1664 0 1 770
box -5 -3 28 105
use FILL  FILL_9519
timestamp 1677622389
transform 1 0 1664 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_361
timestamp 1677622389
transform 1 0 1672 0 1 770
box -8 -3 46 105
use FILL  FILL_9520
timestamp 1677622389
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_9521
timestamp 1677622389
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_9522
timestamp 1677622389
transform 1 0 1728 0 1 770
box -8 -3 16 105
use INVX2  INVX2_601
timestamp 1677622389
transform -1 0 1752 0 1 770
box -9 -3 26 105
use FILL  FILL_9523
timestamp 1677622389
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_9536
timestamp 1677622389
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_9538
timestamp 1677622389
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_9540
timestamp 1677622389
transform 1 0 1776 0 1 770
box -8 -3 16 105
use INVX2  INVX2_603
timestamp 1677622389
transform 1 0 1784 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_7390
timestamp 1677622389
transform 1 0 1836 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_359
timestamp 1677622389
transform -1 0 1840 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_517
timestamp 1677622389
transform -1 0 1936 0 1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_360
timestamp 1677622389
transform 1 0 1936 0 1 770
box -8 -3 46 105
use FILL  FILL_9542
timestamp 1677622389
transform 1 0 1976 0 1 770
box -8 -3 16 105
use FILL  FILL_9543
timestamp 1677622389
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_9544
timestamp 1677622389
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_9545
timestamp 1677622389
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_9546
timestamp 1677622389
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_9547
timestamp 1677622389
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_9548
timestamp 1677622389
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_9549
timestamp 1677622389
transform 1 0 2032 0 1 770
box -8 -3 16 105
use FILL  FILL_9550
timestamp 1677622389
transform 1 0 2040 0 1 770
box -8 -3 16 105
use FILL  FILL_9551
timestamp 1677622389
transform 1 0 2048 0 1 770
box -8 -3 16 105
use INVX2  INVX2_604
timestamp 1677622389
transform 1 0 2056 0 1 770
box -9 -3 26 105
use FILL  FILL_9552
timestamp 1677622389
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_9553
timestamp 1677622389
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_9554
timestamp 1677622389
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_9555
timestamp 1677622389
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_9556
timestamp 1677622389
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_9557
timestamp 1677622389
transform 1 0 2112 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_71
timestamp 1677622389
transform 1 0 2120 0 1 770
box -8 -3 40 105
use FILL  FILL_9569
timestamp 1677622389
transform 1 0 2152 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_72
timestamp 1677622389
transform 1 0 2160 0 1 770
box -8 -3 40 105
use FILL  FILL_9570
timestamp 1677622389
transform 1 0 2192 0 1 770
box -8 -3 16 105
use FILL  FILL_9571
timestamp 1677622389
transform 1 0 2200 0 1 770
box -8 -3 16 105
use FILL  FILL_9572
timestamp 1677622389
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_9573
timestamp 1677622389
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_9574
timestamp 1677622389
transform 1 0 2224 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7391
timestamp 1677622389
transform 1 0 2252 0 1 775
box -3 -3 3 3
use INVX2  INVX2_606
timestamp 1677622389
transform -1 0 2248 0 1 770
box -9 -3 26 105
use INVX2  INVX2_607
timestamp 1677622389
transform 1 0 2248 0 1 770
box -9 -3 26 105
use FILL  FILL_9575
timestamp 1677622389
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_9576
timestamp 1677622389
transform 1 0 2272 0 1 770
box -8 -3 16 105
use FILL  FILL_9577
timestamp 1677622389
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_9578
timestamp 1677622389
transform 1 0 2288 0 1 770
box -8 -3 16 105
use FILL  FILL_9579
timestamp 1677622389
transform 1 0 2296 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_170
timestamp 1677622389
transform -1 0 2336 0 1 770
box -8 -3 34 105
use FAX1  FAX1_19
timestamp 1677622389
transform 1 0 2336 0 1 770
box -5 -3 126 105
use AOI21X1  AOI21X1_16
timestamp 1677622389
transform 1 0 2456 0 1 770
box -7 -3 39 105
use FILL  FILL_9580
timestamp 1677622389
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_9589
timestamp 1677622389
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_9591
timestamp 1677622389
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_9593
timestamp 1677622389
transform 1 0 2512 0 1 770
box -8 -3 16 105
use INVX2  INVX2_608
timestamp 1677622389
transform -1 0 2536 0 1 770
box -9 -3 26 105
use FILL  FILL_9594
timestamp 1677622389
transform 1 0 2536 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_362
timestamp 1677622389
transform 1 0 2544 0 1 770
box -8 -3 46 105
use FILL  FILL_9595
timestamp 1677622389
transform 1 0 2584 0 1 770
box -8 -3 16 105
use FILL  FILL_9596
timestamp 1677622389
transform 1 0 2592 0 1 770
box -8 -3 16 105
use FILL  FILL_9601
timestamp 1677622389
transform 1 0 2600 0 1 770
box -8 -3 16 105
use FILL  FILL_9603
timestamp 1677622389
transform 1 0 2608 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7392
timestamp 1677622389
transform 1 0 2700 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_522
timestamp 1677622389
transform -1 0 2712 0 1 770
box -8 -3 104 105
use FILL  FILL_9604
timestamp 1677622389
transform 1 0 2712 0 1 770
box -8 -3 16 105
use FILL  FILL_9605
timestamp 1677622389
transform 1 0 2720 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7393
timestamp 1677622389
transform 1 0 2740 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_7394
timestamp 1677622389
transform 1 0 2756 0 1 775
box -3 -3 3 3
use FAX1  FAX1_21
timestamp 1677622389
transform 1 0 2728 0 1 770
box -5 -3 126 105
use FILL  FILL_9606
timestamp 1677622389
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FILL  FILL_9607
timestamp 1677622389
transform 1 0 2856 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7395
timestamp 1677622389
transform 1 0 2876 0 1 775
box -3 -3 3 3
use FILL  FILL_9608
timestamp 1677622389
transform 1 0 2864 0 1 770
box -8 -3 16 105
use FAX1  FAX1_22
timestamp 1677622389
transform 1 0 2872 0 1 770
box -5 -3 126 105
use FILL  FILL_9609
timestamp 1677622389
transform 1 0 2992 0 1 770
box -8 -3 16 105
use FILL  FILL_9629
timestamp 1677622389
transform 1 0 3000 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1677622389
transform 1 0 3008 0 1 770
box -8 -3 32 105
use FILL  FILL_9631
timestamp 1677622389
transform 1 0 3032 0 1 770
box -8 -3 16 105
use FILL  FILL_9632
timestamp 1677622389
transform 1 0 3040 0 1 770
box -8 -3 16 105
use FILL  FILL_9635
timestamp 1677622389
transform 1 0 3048 0 1 770
box -8 -3 16 105
use FILL  FILL_9637
timestamp 1677622389
transform 1 0 3056 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_171
timestamp 1677622389
transform -1 0 3096 0 1 770
box -8 -3 34 105
use AOI21X1  AOI21X1_17
timestamp 1677622389
transform -1 0 3128 0 1 770
box -7 -3 39 105
use FILL  FILL_9638
timestamp 1677622389
transform 1 0 3128 0 1 770
box -8 -3 16 105
use FILL  FILL_9639
timestamp 1677622389
transform 1 0 3136 0 1 770
box -8 -3 16 105
use FILL  FILL_9640
timestamp 1677622389
transform 1 0 3144 0 1 770
box -8 -3 16 105
use FILL  FILL_9647
timestamp 1677622389
transform 1 0 3152 0 1 770
box -8 -3 16 105
use FILL  FILL_9649
timestamp 1677622389
transform 1 0 3160 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7396
timestamp 1677622389
transform 1 0 3180 0 1 775
box -3 -3 3 3
use INVX2  INVX2_610
timestamp 1677622389
transform -1 0 3184 0 1 770
box -9 -3 26 105
use FILL  FILL_9650
timestamp 1677622389
transform 1 0 3184 0 1 770
box -8 -3 16 105
use FILL  FILL_9651
timestamp 1677622389
transform 1 0 3192 0 1 770
box -8 -3 16 105
use FILL  FILL_9652
timestamp 1677622389
transform 1 0 3200 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_363
timestamp 1677622389
transform -1 0 3248 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_7397
timestamp 1677622389
transform 1 0 3260 0 1 775
box -3 -3 3 3
use FILL  FILL_9653
timestamp 1677622389
transform 1 0 3248 0 1 770
box -8 -3 16 105
use FILL  FILL_9654
timestamp 1677622389
transform 1 0 3256 0 1 770
box -8 -3 16 105
use FILL  FILL_9655
timestamp 1677622389
transform 1 0 3264 0 1 770
box -8 -3 16 105
use FILL  FILL_9656
timestamp 1677622389
transform 1 0 3272 0 1 770
box -8 -3 16 105
use FILL  FILL_9657
timestamp 1677622389
transform 1 0 3280 0 1 770
box -8 -3 16 105
use FILL  FILL_9658
timestamp 1677622389
transform 1 0 3288 0 1 770
box -8 -3 16 105
use FILL  FILL_9664
timestamp 1677622389
transform 1 0 3296 0 1 770
box -8 -3 16 105
use FILL  FILL_9666
timestamp 1677622389
transform 1 0 3304 0 1 770
box -8 -3 16 105
use FILL  FILL_9668
timestamp 1677622389
transform 1 0 3312 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7398
timestamp 1677622389
transform 1 0 3348 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_365
timestamp 1677622389
transform 1 0 3320 0 1 770
box -8 -3 46 105
use FILL  FILL_9670
timestamp 1677622389
transform 1 0 3360 0 1 770
box -8 -3 16 105
use FAX1  FAX1_23
timestamp 1677622389
transform -1 0 3488 0 1 770
box -5 -3 126 105
use FILL  FILL_9671
timestamp 1677622389
transform 1 0 3488 0 1 770
box -8 -3 16 105
use FILL  FILL_9672
timestamp 1677622389
transform 1 0 3496 0 1 770
box -8 -3 16 105
use FILL  FILL_9673
timestamp 1677622389
transform 1 0 3504 0 1 770
box -8 -3 16 105
use FILL  FILL_9674
timestamp 1677622389
transform 1 0 3512 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_60
timestamp 1677622389
transform 1 0 3520 0 1 770
box -8 -3 40 105
use FILL  FILL_9680
timestamp 1677622389
transform 1 0 3552 0 1 770
box -8 -3 16 105
use FILL  FILL_9681
timestamp 1677622389
transform 1 0 3560 0 1 770
box -8 -3 16 105
use FILL  FILL_9684
timestamp 1677622389
transform 1 0 3568 0 1 770
box -8 -3 16 105
use FILL  FILL_9686
timestamp 1677622389
transform 1 0 3576 0 1 770
box -8 -3 16 105
use FILL  FILL_9688
timestamp 1677622389
transform 1 0 3584 0 1 770
box -8 -3 16 105
use INVX2  INVX2_611
timestamp 1677622389
transform 1 0 3592 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_7399
timestamp 1677622389
transform 1 0 3628 0 1 775
box -3 -3 3 3
use INVX2  INVX2_612
timestamp 1677622389
transform 1 0 3608 0 1 770
box -9 -3 26 105
use FILL  FILL_9690
timestamp 1677622389
transform 1 0 3624 0 1 770
box -8 -3 16 105
use FILL  FILL_9692
timestamp 1677622389
transform 1 0 3632 0 1 770
box -8 -3 16 105
use FILL  FILL_9694
timestamp 1677622389
transform 1 0 3640 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_362
timestamp 1677622389
transform -1 0 3688 0 1 770
box -8 -3 46 105
use FILL  FILL_9695
timestamp 1677622389
transform 1 0 3688 0 1 770
box -8 -3 16 105
use FILL  FILL_9696
timestamp 1677622389
transform 1 0 3696 0 1 770
box -8 -3 16 105
use FILL  FILL_9700
timestamp 1677622389
transform 1 0 3704 0 1 770
box -8 -3 16 105
use FILL  FILL_9702
timestamp 1677622389
transform 1 0 3712 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7400
timestamp 1677622389
transform 1 0 3756 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_364
timestamp 1677622389
transform 1 0 3720 0 1 770
box -8 -3 46 105
use FILL  FILL_9704
timestamp 1677622389
transform 1 0 3760 0 1 770
box -8 -3 16 105
use FILL  FILL_9706
timestamp 1677622389
transform 1 0 3768 0 1 770
box -8 -3 16 105
use FILL  FILL_9708
timestamp 1677622389
transform 1 0 3776 0 1 770
box -8 -3 16 105
use FILL  FILL_9710
timestamp 1677622389
transform 1 0 3784 0 1 770
box -8 -3 16 105
use FILL  FILL_9712
timestamp 1677622389
transform 1 0 3792 0 1 770
box -8 -3 16 105
use FILL  FILL_9713
timestamp 1677622389
transform 1 0 3800 0 1 770
box -8 -3 16 105
use FILL  FILL_9714
timestamp 1677622389
transform 1 0 3808 0 1 770
box -8 -3 16 105
use FILL  FILL_9715
timestamp 1677622389
transform 1 0 3816 0 1 770
box -8 -3 16 105
use FILL  FILL_9716
timestamp 1677622389
transform 1 0 3824 0 1 770
box -8 -3 16 105
use FILL  FILL_9717
timestamp 1677622389
transform 1 0 3832 0 1 770
box -8 -3 16 105
use FILL  FILL_9719
timestamp 1677622389
transform 1 0 3840 0 1 770
box -8 -3 16 105
use FILL  FILL_9721
timestamp 1677622389
transform 1 0 3848 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_175
timestamp 1677622389
transform 1 0 3856 0 1 770
box -8 -3 34 105
use FILL  FILL_9723
timestamp 1677622389
transform 1 0 3888 0 1 770
box -8 -3 16 105
use FILL  FILL_9724
timestamp 1677622389
transform 1 0 3896 0 1 770
box -8 -3 16 105
use FILL  FILL_9725
timestamp 1677622389
transform 1 0 3904 0 1 770
box -8 -3 16 105
use FILL  FILL_9728
timestamp 1677622389
transform 1 0 3912 0 1 770
box -8 -3 16 105
use FILL  FILL_9730
timestamp 1677622389
transform 1 0 3920 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_35
timestamp 1677622389
transform 1 0 3928 0 1 770
box -8 -3 32 105
use FILL  FILL_9732
timestamp 1677622389
transform 1 0 3952 0 1 770
box -8 -3 16 105
use FILL  FILL_9733
timestamp 1677622389
transform 1 0 3960 0 1 770
box -8 -3 16 105
use FILL  FILL_9734
timestamp 1677622389
transform 1 0 3968 0 1 770
box -8 -3 16 105
use FILL  FILL_9735
timestamp 1677622389
transform 1 0 3976 0 1 770
box -8 -3 16 105
use FILL  FILL_9738
timestamp 1677622389
transform 1 0 3984 0 1 770
box -8 -3 16 105
use FILL  FILL_9740
timestamp 1677622389
transform 1 0 3992 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_176
timestamp 1677622389
transform -1 0 4032 0 1 770
box -8 -3 34 105
use FILL  FILL_9741
timestamp 1677622389
transform 1 0 4032 0 1 770
box -8 -3 16 105
use FILL  FILL_9742
timestamp 1677622389
transform 1 0 4040 0 1 770
box -8 -3 16 105
use FILL  FILL_9743
timestamp 1677622389
transform 1 0 4048 0 1 770
box -8 -3 16 105
use FILL  FILL_9744
timestamp 1677622389
transform 1 0 4056 0 1 770
box -8 -3 16 105
use FILL  FILL_9749
timestamp 1677622389
transform 1 0 4064 0 1 770
box -8 -3 16 105
use FILL  FILL_9751
timestamp 1677622389
transform 1 0 4072 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_36
timestamp 1677622389
transform -1 0 4104 0 1 770
box -8 -3 32 105
use FILL  FILL_9752
timestamp 1677622389
transform 1 0 4104 0 1 770
box -8 -3 16 105
use FILL  FILL_9753
timestamp 1677622389
transform 1 0 4112 0 1 770
box -8 -3 16 105
use FILL  FILL_9754
timestamp 1677622389
transform 1 0 4120 0 1 770
box -8 -3 16 105
use FILL  FILL_9755
timestamp 1677622389
transform 1 0 4128 0 1 770
box -8 -3 16 105
use FILL  FILL_9759
timestamp 1677622389
transform 1 0 4136 0 1 770
box -8 -3 16 105
use FILL  FILL_9761
timestamp 1677622389
transform 1 0 4144 0 1 770
box -8 -3 16 105
use FILL  FILL_9763
timestamp 1677622389
transform 1 0 4152 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_371
timestamp 1677622389
transform 1 0 4160 0 1 770
box -8 -3 46 105
use FILL  FILL_9765
timestamp 1677622389
transform 1 0 4200 0 1 770
box -8 -3 16 105
use FILL  FILL_9772
timestamp 1677622389
transform 1 0 4208 0 1 770
box -8 -3 16 105
use FILL  FILL_9774
timestamp 1677622389
transform 1 0 4216 0 1 770
box -8 -3 16 105
use FILL  FILL_9776
timestamp 1677622389
transform 1 0 4224 0 1 770
box -8 -3 16 105
use FILL  FILL_9777
timestamp 1677622389
transform 1 0 4232 0 1 770
box -8 -3 16 105
use FILL  FILL_9778
timestamp 1677622389
transform 1 0 4240 0 1 770
box -8 -3 16 105
use FILL  FILL_9779
timestamp 1677622389
transform 1 0 4248 0 1 770
box -8 -3 16 105
use FILL  FILL_9780
timestamp 1677622389
transform 1 0 4256 0 1 770
box -8 -3 16 105
use FILL  FILL_9781
timestamp 1677622389
transform 1 0 4264 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_373
timestamp 1677622389
transform 1 0 4272 0 1 770
box -8 -3 46 105
use FILL  FILL_9783
timestamp 1677622389
transform 1 0 4312 0 1 770
box -8 -3 16 105
use FILL  FILL_9785
timestamp 1677622389
transform 1 0 4320 0 1 770
box -8 -3 16 105
use FILL  FILL_9786
timestamp 1677622389
transform 1 0 4328 0 1 770
box -8 -3 16 105
use FILL  FILL_9787
timestamp 1677622389
transform 1 0 4336 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_375
timestamp 1677622389
transform 1 0 4344 0 1 770
box -8 -3 46 105
use FILL  FILL_9788
timestamp 1677622389
transform 1 0 4384 0 1 770
box -8 -3 16 105
use FILL  FILL_9789
timestamp 1677622389
transform 1 0 4392 0 1 770
box -8 -3 16 105
use FILL  FILL_9790
timestamp 1677622389
transform 1 0 4400 0 1 770
box -8 -3 16 105
use FILL  FILL_9791
timestamp 1677622389
transform 1 0 4408 0 1 770
box -8 -3 16 105
use FILL  FILL_9792
timestamp 1677622389
transform 1 0 4416 0 1 770
box -8 -3 16 105
use FILL  FILL_9794
timestamp 1677622389
transform 1 0 4424 0 1 770
box -8 -3 16 105
use FILL  FILL_9796
timestamp 1677622389
transform 1 0 4432 0 1 770
box -8 -3 16 105
use FILL  FILL_9798
timestamp 1677622389
transform 1 0 4440 0 1 770
box -8 -3 16 105
use FILL  FILL_9799
timestamp 1677622389
transform 1 0 4448 0 1 770
box -8 -3 16 105
use FILL  FILL_9800
timestamp 1677622389
transform 1 0 4456 0 1 770
box -8 -3 16 105
use FILL  FILL_9801
timestamp 1677622389
transform 1 0 4464 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_378
timestamp 1677622389
transform 1 0 4472 0 1 770
box -8 -3 46 105
use FILL  FILL_9802
timestamp 1677622389
transform 1 0 4512 0 1 770
box -8 -3 16 105
use FILL  FILL_9803
timestamp 1677622389
transform 1 0 4520 0 1 770
box -8 -3 16 105
use FILL  FILL_9804
timestamp 1677622389
transform 1 0 4528 0 1 770
box -8 -3 16 105
use FILL  FILL_9805
timestamp 1677622389
transform 1 0 4536 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_379
timestamp 1677622389
transform 1 0 4544 0 1 770
box -8 -3 46 105
use FILL  FILL_9806
timestamp 1677622389
transform 1 0 4584 0 1 770
box -8 -3 16 105
use FILL  FILL_9807
timestamp 1677622389
transform 1 0 4592 0 1 770
box -8 -3 16 105
use FILL  FILL_9808
timestamp 1677622389
transform 1 0 4600 0 1 770
box -8 -3 16 105
use FILL  FILL_9809
timestamp 1677622389
transform 1 0 4608 0 1 770
box -8 -3 16 105
use FILL  FILL_9810
timestamp 1677622389
transform 1 0 4616 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_380
timestamp 1677622389
transform -1 0 4664 0 1 770
box -8 -3 46 105
use FILL  FILL_9811
timestamp 1677622389
transform 1 0 4664 0 1 770
box -8 -3 16 105
use FILL  FILL_9812
timestamp 1677622389
transform 1 0 4672 0 1 770
box -8 -3 16 105
use FILL  FILL_9813
timestamp 1677622389
transform 1 0 4680 0 1 770
box -8 -3 16 105
use FILL  FILL_9814
timestamp 1677622389
transform 1 0 4688 0 1 770
box -8 -3 16 105
use FILL  FILL_9827
timestamp 1677622389
transform 1 0 4696 0 1 770
box -8 -3 16 105
use FILL  FILL_9829
timestamp 1677622389
transform 1 0 4704 0 1 770
box -8 -3 16 105
use INVX2  INVX2_614
timestamp 1677622389
transform -1 0 4728 0 1 770
box -9 -3 26 105
use FILL  FILL_9830
timestamp 1677622389
transform 1 0 4728 0 1 770
box -8 -3 16 105
use FILL  FILL_9831
timestamp 1677622389
transform 1 0 4736 0 1 770
box -8 -3 16 105
use FILL  FILL_9832
timestamp 1677622389
transform 1 0 4744 0 1 770
box -8 -3 16 105
use FILL  FILL_9833
timestamp 1677622389
transform 1 0 4752 0 1 770
box -8 -3 16 105
use FILL  FILL_9834
timestamp 1677622389
transform 1 0 4760 0 1 770
box -8 -3 16 105
use FILL  FILL_9835
timestamp 1677622389
transform 1 0 4768 0 1 770
box -8 -3 16 105
use FILL  FILL_9836
timestamp 1677622389
transform 1 0 4776 0 1 770
box -8 -3 16 105
use FILL  FILL_9840
timestamp 1677622389
transform 1 0 4784 0 1 770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_79
timestamp 1677622389
transform 1 0 4819 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_7440
timestamp 1677622389
transform 1 0 164 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8395
timestamp 1677622389
transform 1 0 84 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7441
timestamp 1677622389
transform 1 0 196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8396
timestamp 1677622389
transform 1 0 188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8397
timestamp 1677622389
transform 1 0 196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8398
timestamp 1677622389
transform 1 0 220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8513
timestamp 1677622389
transform 1 0 132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8514
timestamp 1677622389
transform 1 0 164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8515
timestamp 1677622389
transform 1 0 172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8516
timestamp 1677622389
transform 1 0 180 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7541
timestamp 1677622389
transform 1 0 132 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7542
timestamp 1677622389
transform 1 0 172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7543
timestamp 1677622389
transform 1 0 188 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7579
timestamp 1677622389
transform 1 0 180 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8399
timestamp 1677622389
transform 1 0 244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8517
timestamp 1677622389
transform 1 0 212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8518
timestamp 1677622389
transform 1 0 228 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7544
timestamp 1677622389
transform 1 0 212 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7513
timestamp 1677622389
transform 1 0 244 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8519
timestamp 1677622389
transform 1 0 252 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7580
timestamp 1677622389
transform 1 0 236 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7626
timestamp 1677622389
transform 1 0 228 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7442
timestamp 1677622389
transform 1 0 292 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7421
timestamp 1677622389
transform 1 0 348 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7443
timestamp 1677622389
transform 1 0 316 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7444
timestamp 1677622389
transform 1 0 340 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8400
timestamp 1677622389
transform 1 0 292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8401
timestamp 1677622389
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8402
timestamp 1677622389
transform 1 0 316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8403
timestamp 1677622389
transform 1 0 332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8520
timestamp 1677622389
transform 1 0 292 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7514
timestamp 1677622389
transform 1 0 300 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7491
timestamp 1677622389
transform 1 0 340 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8404
timestamp 1677622389
transform 1 0 348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8521
timestamp 1677622389
transform 1 0 308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8522
timestamp 1677622389
transform 1 0 324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8523
timestamp 1677622389
transform 1 0 340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7545
timestamp 1677622389
transform 1 0 324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7613
timestamp 1677622389
transform 1 0 340 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8524
timestamp 1677622389
transform 1 0 356 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7581
timestamp 1677622389
transform 1 0 356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7546
timestamp 1677622389
transform 1 0 372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7445
timestamp 1677622389
transform 1 0 388 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7614
timestamp 1677622389
transform 1 0 380 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7401
timestamp 1677622389
transform 1 0 420 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8405
timestamp 1677622389
transform 1 0 396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8406
timestamp 1677622389
transform 1 0 412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8407
timestamp 1677622389
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8408
timestamp 1677622389
transform 1 0 428 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7515
timestamp 1677622389
transform 1 0 396 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8525
timestamp 1677622389
transform 1 0 404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7547
timestamp 1677622389
transform 1 0 404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7615
timestamp 1677622389
transform 1 0 396 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7548
timestamp 1677622389
transform 1 0 428 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7446
timestamp 1677622389
transform 1 0 452 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8526
timestamp 1677622389
transform 1 0 452 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7402
timestamp 1677622389
transform 1 0 492 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7422
timestamp 1677622389
transform 1 0 548 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7447
timestamp 1677622389
transform 1 0 484 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8409
timestamp 1677622389
transform 1 0 484 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7516
timestamp 1677622389
transform 1 0 508 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8527
timestamp 1677622389
transform 1 0 532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8528
timestamp 1677622389
transform 1 0 564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8529
timestamp 1677622389
transform 1 0 572 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7549
timestamp 1677622389
transform 1 0 532 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7550
timestamp 1677622389
transform 1 0 572 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7423
timestamp 1677622389
transform 1 0 588 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8410
timestamp 1677622389
transform 1 0 588 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7517
timestamp 1677622389
transform 1 0 596 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7551
timestamp 1677622389
transform 1 0 644 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7448
timestamp 1677622389
transform 1 0 660 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8411
timestamp 1677622389
transform 1 0 660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8530
timestamp 1677622389
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8531
timestamp 1677622389
transform 1 0 740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7552
timestamp 1677622389
transform 1 0 708 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7616
timestamp 1677622389
transform 1 0 684 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8532
timestamp 1677622389
transform 1 0 756 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7553
timestamp 1677622389
transform 1 0 756 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7424
timestamp 1677622389
transform 1 0 780 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8412
timestamp 1677622389
transform 1 0 772 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7403
timestamp 1677622389
transform 1 0 828 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7425
timestamp 1677622389
transform 1 0 836 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7449
timestamp 1677622389
transform 1 0 796 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7450
timestamp 1677622389
transform 1 0 812 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8413
timestamp 1677622389
transform 1 0 796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8414
timestamp 1677622389
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8415
timestamp 1677622389
transform 1 0 836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8533
timestamp 1677622389
transform 1 0 804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8534
timestamp 1677622389
transform 1 0 812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8535
timestamp 1677622389
transform 1 0 828 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7518
timestamp 1677622389
transform 1 0 836 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8416
timestamp 1677622389
transform 1 0 852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8536
timestamp 1677622389
transform 1 0 844 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7554
timestamp 1677622389
transform 1 0 804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7519
timestamp 1677622389
transform 1 0 852 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7555
timestamp 1677622389
transform 1 0 844 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7582
timestamp 1677622389
transform 1 0 820 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7583
timestamp 1677622389
transform 1 0 836 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7617
timestamp 1677622389
transform 1 0 812 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7556
timestamp 1677622389
transform 1 0 860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7618
timestamp 1677622389
transform 1 0 876 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7426
timestamp 1677622389
transform 1 0 916 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7451
timestamp 1677622389
transform 1 0 964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7452
timestamp 1677622389
transform 1 0 996 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8417
timestamp 1677622389
transform 1 0 996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8537
timestamp 1677622389
transform 1 0 908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8538
timestamp 1677622389
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8539
timestamp 1677622389
transform 1 0 948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7557
timestamp 1677622389
transform 1 0 908 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7558
timestamp 1677622389
transform 1 0 948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7619
timestamp 1677622389
transform 1 0 980 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8392
timestamp 1677622389
transform 1 0 1012 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_7492
timestamp 1677622389
transform 1 0 1012 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7427
timestamp 1677622389
transform 1 0 1076 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8418
timestamp 1677622389
transform 1 0 1068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8540
timestamp 1677622389
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7404
timestamp 1677622389
transform 1 0 1132 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7453
timestamp 1677622389
transform 1 0 1092 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7454
timestamp 1677622389
transform 1 0 1132 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8419
timestamp 1677622389
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8541
timestamp 1677622389
transform 1 0 1140 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7620
timestamp 1677622389
transform 1 0 1108 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7621
timestamp 1677622389
transform 1 0 1156 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7455
timestamp 1677622389
transform 1 0 1196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8420
timestamp 1677622389
transform 1 0 1180 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7493
timestamp 1677622389
transform 1 0 1188 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8421
timestamp 1677622389
transform 1 0 1196 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7494
timestamp 1677622389
transform 1 0 1212 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8422
timestamp 1677622389
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8542
timestamp 1677622389
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8543
timestamp 1677622389
transform 1 0 1196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8544
timestamp 1677622389
transform 1 0 1212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8545
timestamp 1677622389
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7584
timestamp 1677622389
transform 1 0 1196 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7456
timestamp 1677622389
transform 1 0 1244 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8423
timestamp 1677622389
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8546
timestamp 1677622389
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8547
timestamp 1677622389
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7457
timestamp 1677622389
transform 1 0 1324 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8424
timestamp 1677622389
transform 1 0 1324 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7405
timestamp 1677622389
transform 1 0 1340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7406
timestamp 1677622389
transform 1 0 1372 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7407
timestamp 1677622389
transform 1 0 1420 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8425
timestamp 1677622389
transform 1 0 1340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8426
timestamp 1677622389
transform 1 0 1428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8548
timestamp 1677622389
transform 1 0 1364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8549
timestamp 1677622389
transform 1 0 1420 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7585
timestamp 1677622389
transform 1 0 1428 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7458
timestamp 1677622389
transform 1 0 1476 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8427
timestamp 1677622389
transform 1 0 1476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8550
timestamp 1677622389
transform 1 0 1452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8551
timestamp 1677622389
transform 1 0 1468 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7520
timestamp 1677622389
transform 1 0 1476 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8428
timestamp 1677622389
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8552
timestamp 1677622389
transform 1 0 1484 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7521
timestamp 1677622389
transform 1 0 1492 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7408
timestamp 1677622389
transform 1 0 1612 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7428
timestamp 1677622389
transform 1 0 1596 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7495
timestamp 1677622389
transform 1 0 1540 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7496
timestamp 1677622389
transform 1 0 1580 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8429
timestamp 1677622389
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8553
timestamp 1677622389
transform 1 0 1532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8554
timestamp 1677622389
transform 1 0 1540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8555
timestamp 1677622389
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7559
timestamp 1677622389
transform 1 0 1532 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7560
timestamp 1677622389
transform 1 0 1572 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7429
timestamp 1677622389
transform 1 0 1636 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7409
timestamp 1677622389
transform 1 0 1660 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7430
timestamp 1677622389
transform 1 0 1740 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8430
timestamp 1677622389
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8556
timestamp 1677622389
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8557
timestamp 1677622389
transform 1 0 1740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8558
timestamp 1677622389
transform 1 0 1764 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7586
timestamp 1677622389
transform 1 0 1788 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8431
timestamp 1677622389
transform 1 0 1828 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7522
timestamp 1677622389
transform 1 0 1828 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7410
timestamp 1677622389
transform 1 0 1876 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8432
timestamp 1677622389
transform 1 0 1876 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7497
timestamp 1677622389
transform 1 0 1884 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8433
timestamp 1677622389
transform 1 0 1892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8559
timestamp 1677622389
transform 1 0 1860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8560
timestamp 1677622389
transform 1 0 1868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7561
timestamp 1677622389
transform 1 0 1860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7523
timestamp 1677622389
transform 1 0 1876 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8561
timestamp 1677622389
transform 1 0 1884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8562
timestamp 1677622389
transform 1 0 1900 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7587
timestamp 1677622389
transform 1 0 1868 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7588
timestamp 1677622389
transform 1 0 1900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7411
timestamp 1677622389
transform 1 0 1940 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7412
timestamp 1677622389
transform 1 0 1956 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7459
timestamp 1677622389
transform 1 0 1996 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8434
timestamp 1677622389
transform 1 0 1996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8563
timestamp 1677622389
transform 1 0 1948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7524
timestamp 1677622389
transform 1 0 1996 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7562
timestamp 1677622389
transform 1 0 1948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7589
timestamp 1677622389
transform 1 0 1932 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7590
timestamp 1677622389
transform 1 0 1972 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7460
timestamp 1677622389
transform 1 0 2012 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8435
timestamp 1677622389
transform 1 0 2100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8564
timestamp 1677622389
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7525
timestamp 1677622389
transform 1 0 2036 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8565
timestamp 1677622389
transform 1 0 2068 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7526
timestamp 1677622389
transform 1 0 2100 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7461
timestamp 1677622389
transform 1 0 2204 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8436
timestamp 1677622389
transform 1 0 2140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8566
timestamp 1677622389
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8567
timestamp 1677622389
transform 1 0 2220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8568
timestamp 1677622389
transform 1 0 2228 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7627
timestamp 1677622389
transform 1 0 2148 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7462
timestamp 1677622389
transform 1 0 2316 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8437
timestamp 1677622389
transform 1 0 2316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8569
timestamp 1677622389
transform 1 0 2292 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7591
timestamp 1677622389
transform 1 0 2276 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7628
timestamp 1677622389
transform 1 0 2252 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8393
timestamp 1677622389
transform 1 0 2356 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_7463
timestamp 1677622389
transform 1 0 2364 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7464
timestamp 1677622389
transform 1 0 2460 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8438
timestamp 1677622389
transform 1 0 2348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8570
timestamp 1677622389
transform 1 0 2444 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7592
timestamp 1677622389
transform 1 0 2380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7593
timestamp 1677622389
transform 1 0 2420 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8439
timestamp 1677622389
transform 1 0 2468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8440
timestamp 1677622389
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8441
timestamp 1677622389
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7594
timestamp 1677622389
transform 1 0 2500 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8394
timestamp 1677622389
transform 1 0 2524 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_7498
timestamp 1677622389
transform 1 0 2524 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8571
timestamp 1677622389
transform 1 0 2524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7563
timestamp 1677622389
transform 1 0 2524 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8572
timestamp 1677622389
transform 1 0 2556 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7595
timestamp 1677622389
transform 1 0 2556 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7499
timestamp 1677622389
transform 1 0 2572 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8573
timestamp 1677622389
transform 1 0 2572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8574
timestamp 1677622389
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8575
timestamp 1677622389
transform 1 0 2604 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7564
timestamp 1677622389
transform 1 0 2604 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7596
timestamp 1677622389
transform 1 0 2596 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8638
timestamp 1677622389
transform 1 0 2644 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7597
timestamp 1677622389
transform 1 0 2668 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7413
timestamp 1677622389
transform 1 0 2748 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8442
timestamp 1677622389
transform 1 0 2756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8576
timestamp 1677622389
transform 1 0 2732 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7414
timestamp 1677622389
transform 1 0 2772 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8577
timestamp 1677622389
transform 1 0 2772 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7465
timestamp 1677622389
transform 1 0 2812 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8443
timestamp 1677622389
transform 1 0 2812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8444
timestamp 1677622389
transform 1 0 2820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8578
timestamp 1677622389
transform 1 0 2804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7466
timestamp 1677622389
transform 1 0 2876 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8445
timestamp 1677622389
transform 1 0 2876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8579
timestamp 1677622389
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7565
timestamp 1677622389
transform 1 0 2852 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8580
timestamp 1677622389
transform 1 0 2892 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7467
timestamp 1677622389
transform 1 0 2924 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8446
timestamp 1677622389
transform 1 0 2924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8581
timestamp 1677622389
transform 1 0 2916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7598
timestamp 1677622389
transform 1 0 2916 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8447
timestamp 1677622389
transform 1 0 2972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8448
timestamp 1677622389
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7527
timestamp 1677622389
transform 1 0 2988 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8639
timestamp 1677622389
transform 1 0 2988 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7566
timestamp 1677622389
transform 1 0 2996 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8582
timestamp 1677622389
transform 1 0 3020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7567
timestamp 1677622389
transform 1 0 3020 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8449
timestamp 1677622389
transform 1 0 3044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8640
timestamp 1677622389
transform 1 0 3036 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7528
timestamp 1677622389
transform 1 0 3052 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7599
timestamp 1677622389
transform 1 0 3044 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7415
timestamp 1677622389
transform 1 0 3060 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7468
timestamp 1677622389
transform 1 0 3068 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8450
timestamp 1677622389
transform 1 0 3068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8583
timestamp 1677622389
transform 1 0 3068 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7600
timestamp 1677622389
transform 1 0 3068 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7416
timestamp 1677622389
transform 1 0 3092 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8641
timestamp 1677622389
transform 1 0 3084 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7622
timestamp 1677622389
transform 1 0 3076 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8584
timestamp 1677622389
transform 1 0 3100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8585
timestamp 1677622389
transform 1 0 3132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7568
timestamp 1677622389
transform 1 0 3132 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7601
timestamp 1677622389
transform 1 0 3116 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8647
timestamp 1677622389
transform 1 0 3124 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_7417
timestamp 1677622389
transform 1 0 3164 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7431
timestamp 1677622389
transform 1 0 3188 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7432
timestamp 1677622389
transform 1 0 3204 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7469
timestamp 1677622389
transform 1 0 3172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8451
timestamp 1677622389
transform 1 0 3172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8642
timestamp 1677622389
transform 1 0 3164 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7623
timestamp 1677622389
transform 1 0 3164 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8586
timestamp 1677622389
transform 1 0 3196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8587
timestamp 1677622389
transform 1 0 3220 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7569
timestamp 1677622389
transform 1 0 3196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7570
timestamp 1677622389
transform 1 0 3220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7433
timestamp 1677622389
transform 1 0 3252 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7470
timestamp 1677622389
transform 1 0 3244 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8452
timestamp 1677622389
transform 1 0 3244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8453
timestamp 1677622389
transform 1 0 3260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8588
timestamp 1677622389
transform 1 0 3268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8589
timestamp 1677622389
transform 1 0 3300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8454
timestamp 1677622389
transform 1 0 3316 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7418
timestamp 1677622389
transform 1 0 3340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7419
timestamp 1677622389
transform 1 0 3420 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7471
timestamp 1677622389
transform 1 0 3420 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8512
timestamp 1677622389
transform 1 0 3332 0 1 733
box -2 -2 2 2
use M2_M1  M2_M1_8455
timestamp 1677622389
transform 1 0 3420 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7500
timestamp 1677622389
transform 1 0 3428 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8590
timestamp 1677622389
transform 1 0 3380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8591
timestamp 1677622389
transform 1 0 3412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8592
timestamp 1677622389
transform 1 0 3428 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7624
timestamp 1677622389
transform 1 0 3380 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8456
timestamp 1677622389
transform 1 0 3468 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7472
timestamp 1677622389
transform 1 0 3484 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8457
timestamp 1677622389
transform 1 0 3484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8593
timestamp 1677622389
transform 1 0 3476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7473
timestamp 1677622389
transform 1 0 3516 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8458
timestamp 1677622389
transform 1 0 3508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8459
timestamp 1677622389
transform 1 0 3516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8594
timestamp 1677622389
transform 1 0 3516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8643
timestamp 1677622389
transform 1 0 3524 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7602
timestamp 1677622389
transform 1 0 3524 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7474
timestamp 1677622389
transform 1 0 3564 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8460
timestamp 1677622389
transform 1 0 3556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8644
timestamp 1677622389
transform 1 0 3556 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7603
timestamp 1677622389
transform 1 0 3556 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8461
timestamp 1677622389
transform 1 0 3564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8595
timestamp 1677622389
transform 1 0 3572 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7501
timestamp 1677622389
transform 1 0 3588 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8462
timestamp 1677622389
transform 1 0 3596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8463
timestamp 1677622389
transform 1 0 3620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8645
timestamp 1677622389
transform 1 0 3620 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7604
timestamp 1677622389
transform 1 0 3612 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7475
timestamp 1677622389
transform 1 0 3660 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8464
timestamp 1677622389
transform 1 0 3660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8465
timestamp 1677622389
transform 1 0 3676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8596
timestamp 1677622389
transform 1 0 3644 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7571
timestamp 1677622389
transform 1 0 3636 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7529
timestamp 1677622389
transform 1 0 3652 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8646
timestamp 1677622389
transform 1 0 3644 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7572
timestamp 1677622389
transform 1 0 3652 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7502
timestamp 1677622389
transform 1 0 3684 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7476
timestamp 1677622389
transform 1 0 3700 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8466
timestamp 1677622389
transform 1 0 3692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8467
timestamp 1677622389
transform 1 0 3700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8597
timestamp 1677622389
transform 1 0 3668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7530
timestamp 1677622389
transform 1 0 3676 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8598
timestamp 1677622389
transform 1 0 3684 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7605
timestamp 1677622389
transform 1 0 3668 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7503
timestamp 1677622389
transform 1 0 3724 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8468
timestamp 1677622389
transform 1 0 3740 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7504
timestamp 1677622389
transform 1 0 3748 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8469
timestamp 1677622389
transform 1 0 3756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8599
timestamp 1677622389
transform 1 0 3732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8600
timestamp 1677622389
transform 1 0 3748 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7531
timestamp 1677622389
transform 1 0 3756 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8601
timestamp 1677622389
transform 1 0 3764 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7629
timestamp 1677622389
transform 1 0 3732 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7606
timestamp 1677622389
transform 1 0 3764 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7477
timestamp 1677622389
transform 1 0 3796 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8470
timestamp 1677622389
transform 1 0 3796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8471
timestamp 1677622389
transform 1 0 3812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8602
timestamp 1677622389
transform 1 0 3788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7532
timestamp 1677622389
transform 1 0 3812 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8603
timestamp 1677622389
transform 1 0 3820 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7420
timestamp 1677622389
transform 1 0 3900 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8472
timestamp 1677622389
transform 1 0 3868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8473
timestamp 1677622389
transform 1 0 3884 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7505
timestamp 1677622389
transform 1 0 3892 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8474
timestamp 1677622389
transform 1 0 3900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8604
timestamp 1677622389
transform 1 0 3876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8605
timestamp 1677622389
transform 1 0 3892 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7630
timestamp 1677622389
transform 1 0 3892 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7478
timestamp 1677622389
transform 1 0 3940 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8475
timestamp 1677622389
transform 1 0 3940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8476
timestamp 1677622389
transform 1 0 3956 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7506
timestamp 1677622389
transform 1 0 3964 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7479
timestamp 1677622389
transform 1 0 3980 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8477
timestamp 1677622389
transform 1 0 3972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8478
timestamp 1677622389
transform 1 0 3980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8606
timestamp 1677622389
transform 1 0 3948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7533
timestamp 1677622389
transform 1 0 3956 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8607
timestamp 1677622389
transform 1 0 3964 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7607
timestamp 1677622389
transform 1 0 3948 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8479
timestamp 1677622389
transform 1 0 4004 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7534
timestamp 1677622389
transform 1 0 4012 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8480
timestamp 1677622389
transform 1 0 4036 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7507
timestamp 1677622389
transform 1 0 4044 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8481
timestamp 1677622389
transform 1 0 4052 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8608
timestamp 1677622389
transform 1 0 4020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8609
timestamp 1677622389
transform 1 0 4044 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7608
timestamp 1677622389
transform 1 0 4028 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7631
timestamp 1677622389
transform 1 0 4020 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8610
timestamp 1677622389
transform 1 0 4076 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7609
timestamp 1677622389
transform 1 0 4076 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7480
timestamp 1677622389
transform 1 0 4092 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8482
timestamp 1677622389
transform 1 0 4092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8483
timestamp 1677622389
transform 1 0 4108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8484
timestamp 1677622389
transform 1 0 4124 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7535
timestamp 1677622389
transform 1 0 4108 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8611
timestamp 1677622389
transform 1 0 4116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7632
timestamp 1677622389
transform 1 0 4108 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8612
timestamp 1677622389
transform 1 0 4132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7481
timestamp 1677622389
transform 1 0 4140 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7610
timestamp 1677622389
transform 1 0 4132 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7482
timestamp 1677622389
transform 1 0 4156 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7536
timestamp 1677622389
transform 1 0 4172 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7633
timestamp 1677622389
transform 1 0 4164 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8485
timestamp 1677622389
transform 1 0 4196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8613
timestamp 1677622389
transform 1 0 4188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7483
timestamp 1677622389
transform 1 0 4228 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8486
timestamp 1677622389
transform 1 0 4228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8487
timestamp 1677622389
transform 1 0 4244 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7508
timestamp 1677622389
transform 1 0 4252 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7434
timestamp 1677622389
transform 1 0 4276 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7484
timestamp 1677622389
transform 1 0 4268 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8488
timestamp 1677622389
transform 1 0 4260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8489
timestamp 1677622389
transform 1 0 4268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8614
timestamp 1677622389
transform 1 0 4236 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7537
timestamp 1677622389
transform 1 0 4244 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8615
timestamp 1677622389
transform 1 0 4252 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7573
timestamp 1677622389
transform 1 0 4236 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8616
timestamp 1677622389
transform 1 0 4268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7435
timestamp 1677622389
transform 1 0 4308 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8490
timestamp 1677622389
transform 1 0 4292 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7509
timestamp 1677622389
transform 1 0 4300 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8491
timestamp 1677622389
transform 1 0 4308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8617
timestamp 1677622389
transform 1 0 4300 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7634
timestamp 1677622389
transform 1 0 4268 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7436
timestamp 1677622389
transform 1 0 4340 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7485
timestamp 1677622389
transform 1 0 4332 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7510
timestamp 1677622389
transform 1 0 4324 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7437
timestamp 1677622389
transform 1 0 4380 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7486
timestamp 1677622389
transform 1 0 4372 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7487
timestamp 1677622389
transform 1 0 4412 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8492
timestamp 1677622389
transform 1 0 4340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8493
timestamp 1677622389
transform 1 0 4356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8494
timestamp 1677622389
transform 1 0 4372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8495
timestamp 1677622389
transform 1 0 4380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8496
timestamp 1677622389
transform 1 0 4396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8497
timestamp 1677622389
transform 1 0 4412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8618
timestamp 1677622389
transform 1 0 4324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8619
timestamp 1677622389
transform 1 0 4332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8620
timestamp 1677622389
transform 1 0 4340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8621
timestamp 1677622389
transform 1 0 4348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8622
timestamp 1677622389
transform 1 0 4364 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7635
timestamp 1677622389
transform 1 0 4340 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8623
timestamp 1677622389
transform 1 0 4388 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7538
timestamp 1677622389
transform 1 0 4396 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8624
timestamp 1677622389
transform 1 0 4404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7574
timestamp 1677622389
transform 1 0 4388 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7636
timestamp 1677622389
transform 1 0 4388 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8625
timestamp 1677622389
transform 1 0 4428 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7637
timestamp 1677622389
transform 1 0 4428 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8498
timestamp 1677622389
transform 1 0 4444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8499
timestamp 1677622389
transform 1 0 4460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8626
timestamp 1677622389
transform 1 0 4468 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7575
timestamp 1677622389
transform 1 0 4444 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8500
timestamp 1677622389
transform 1 0 4484 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7611
timestamp 1677622389
transform 1 0 4476 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8627
timestamp 1677622389
transform 1 0 4492 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7612
timestamp 1677622389
transform 1 0 4492 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7488
timestamp 1677622389
transform 1 0 4508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7438
timestamp 1677622389
transform 1 0 4540 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7489
timestamp 1677622389
transform 1 0 4548 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8501
timestamp 1677622389
transform 1 0 4508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8502
timestamp 1677622389
transform 1 0 4524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8503
timestamp 1677622389
transform 1 0 4540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8504
timestamp 1677622389
transform 1 0 4548 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7539
timestamp 1677622389
transform 1 0 4524 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8628
timestamp 1677622389
transform 1 0 4532 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7576
timestamp 1677622389
transform 1 0 4532 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8629
timestamp 1677622389
transform 1 0 4564 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7540
timestamp 1677622389
transform 1 0 4572 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7638
timestamp 1677622389
transform 1 0 4564 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7439
timestamp 1677622389
transform 1 0 4612 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8505
timestamp 1677622389
transform 1 0 4596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8506
timestamp 1677622389
transform 1 0 4612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8630
timestamp 1677622389
transform 1 0 4604 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7639
timestamp 1677622389
transform 1 0 4628 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8507
timestamp 1677622389
transform 1 0 4652 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7511
timestamp 1677622389
transform 1 0 4660 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8508
timestamp 1677622389
transform 1 0 4668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8631
timestamp 1677622389
transform 1 0 4660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8632
timestamp 1677622389
transform 1 0 4676 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7640
timestamp 1677622389
transform 1 0 4652 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7490
timestamp 1677622389
transform 1 0 4692 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8509
timestamp 1677622389
transform 1 0 4700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8633
timestamp 1677622389
transform 1 0 4692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8510
timestamp 1677622389
transform 1 0 4732 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7512
timestamp 1677622389
transform 1 0 4740 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8511
timestamp 1677622389
transform 1 0 4748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8634
timestamp 1677622389
transform 1 0 4724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8635
timestamp 1677622389
transform 1 0 4740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7577
timestamp 1677622389
transform 1 0 4724 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7641
timestamp 1677622389
transform 1 0 4716 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7642
timestamp 1677622389
transform 1 0 4740 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8636
timestamp 1677622389
transform 1 0 4756 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7578
timestamp 1677622389
transform 1 0 4756 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8637
timestamp 1677622389
transform 1 0 4788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7625
timestamp 1677622389
transform 1 0 4868 0 1 695
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_80
timestamp 1677622389
transform 1 0 24 0 1 670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_506
timestamp 1677622389
transform 1 0 72 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_590
timestamp 1677622389
transform -1 0 184 0 -1 770
box -9 -3 26 105
use FILL  FILL_9433
timestamp 1677622389
transform 1 0 184 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_347
timestamp 1677622389
transform -1 0 232 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_348
timestamp 1677622389
transform 1 0 232 0 -1 770
box -8 -3 46 105
use FILL  FILL_9434
timestamp 1677622389
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_9435
timestamp 1677622389
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_9436
timestamp 1677622389
transform 1 0 288 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_591
timestamp 1677622389
transform 1 0 296 0 -1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_355
timestamp 1677622389
transform 1 0 312 0 -1 770
box -8 -3 46 105
use FILL  FILL_9437
timestamp 1677622389
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_9438
timestamp 1677622389
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_9439
timestamp 1677622389
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_9440
timestamp 1677622389
transform 1 0 376 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_349
timestamp 1677622389
transform -1 0 424 0 -1 770
box -8 -3 46 105
use FILL  FILL_9441
timestamp 1677622389
transform 1 0 424 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_593
timestamp 1677622389
transform 1 0 432 0 -1 770
box -9 -3 26 105
use FILL  FILL_9460
timestamp 1677622389
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_9461
timestamp 1677622389
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_9462
timestamp 1677622389
transform 1 0 464 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_507
timestamp 1677622389
transform 1 0 472 0 -1 770
box -8 -3 104 105
use FILL  FILL_9463
timestamp 1677622389
transform 1 0 568 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_594
timestamp 1677622389
transform -1 0 592 0 -1 770
box -9 -3 26 105
use FILL  FILL_9464
timestamp 1677622389
transform 1 0 592 0 -1 770
box -8 -3 16 105
use FILL  FILL_9465
timestamp 1677622389
transform 1 0 600 0 -1 770
box -8 -3 16 105
use FILL  FILL_9466
timestamp 1677622389
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9467
timestamp 1677622389
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_9468
timestamp 1677622389
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9469
timestamp 1677622389
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9470
timestamp 1677622389
transform 1 0 640 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_508
timestamp 1677622389
transform 1 0 648 0 -1 770
box -8 -3 104 105
use FILL  FILL_9471
timestamp 1677622389
transform 1 0 744 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_108
timestamp 1677622389
transform 1 0 752 0 -1 770
box -5 -3 28 105
use FILL  FILL_9472
timestamp 1677622389
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9473
timestamp 1677622389
transform 1 0 784 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_595
timestamp 1677622389
transform 1 0 792 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_353
timestamp 1677622389
transform 1 0 808 0 -1 770
box -8 -3 46 105
use FILL  FILL_9474
timestamp 1677622389
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_9476
timestamp 1677622389
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_9479
timestamp 1677622389
transform 1 0 864 0 -1 770
box -8 -3 16 105
use FILL  FILL_9480
timestamp 1677622389
transform 1 0 872 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_597
timestamp 1677622389
transform 1 0 880 0 -1 770
box -9 -3 26 105
use FILL  FILL_9481
timestamp 1677622389
transform 1 0 896 0 -1 770
box -8 -3 16 105
use FILL  FILL_9482
timestamp 1677622389
transform 1 0 904 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_510
timestamp 1677622389
transform -1 0 1008 0 -1 770
box -8 -3 104 105
use FILL  FILL_9483
timestamp 1677622389
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_9485
timestamp 1677622389
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_93
timestamp 1677622389
transform 1 0 1024 0 -1 770
box -8 -3 32 105
use FILL  FILL_9490
timestamp 1677622389
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use FILL  FILL_9491
timestamp 1677622389
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_9492
timestamp 1677622389
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_9493
timestamp 1677622389
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_512
timestamp 1677622389
transform 1 0 1080 0 -1 770
box -8 -3 104 105
use FILL  FILL_9501
timestamp 1677622389
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_9502
timestamp 1677622389
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_355
timestamp 1677622389
transform 1 0 1192 0 -1 770
box -8 -3 46 105
use FILL  FILL_9503
timestamp 1677622389
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_9504
timestamp 1677622389
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_9505
timestamp 1677622389
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_9506
timestamp 1677622389
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_359
timestamp 1677622389
transform -1 0 1304 0 -1 770
box -8 -3 46 105
use FILL  FILL_9507
timestamp 1677622389
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_9509
timestamp 1677622389
transform 1 0 1312 0 -1 770
box -8 -3 16 105
use FILL  FILL_9524
timestamp 1677622389
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_514
timestamp 1677622389
transform 1 0 1328 0 -1 770
box -8 -3 104 105
use FILL  FILL_9525
timestamp 1677622389
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_9526
timestamp 1677622389
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_9527
timestamp 1677622389
transform 1 0 1440 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_358
timestamp 1677622389
transform 1 0 1448 0 -1 770
box -8 -3 46 105
use FILL  FILL_9528
timestamp 1677622389
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_9529
timestamp 1677622389
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_602
timestamp 1677622389
transform 1 0 1504 0 -1 770
box -9 -3 26 105
use FILL  FILL_9530
timestamp 1677622389
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_9531
timestamp 1677622389
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_515
timestamp 1677622389
transform -1 0 1632 0 -1 770
box -8 -3 104 105
use FILL  FILL_9532
timestamp 1677622389
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9533
timestamp 1677622389
transform 1 0 1640 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_516
timestamp 1677622389
transform 1 0 1648 0 -1 770
box -8 -3 104 105
use FILL  FILL_9534
timestamp 1677622389
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_9535
timestamp 1677622389
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_9537
timestamp 1677622389
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_9539
timestamp 1677622389
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_9541
timestamp 1677622389
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9558
timestamp 1677622389
transform 1 0 1784 0 -1 770
box -8 -3 16 105
use FILL  FILL_9559
timestamp 1677622389
transform 1 0 1792 0 -1 770
box -8 -3 16 105
use FILL  FILL_9560
timestamp 1677622389
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_9561
timestamp 1677622389
transform 1 0 1808 0 -1 770
box -8 -3 16 105
use FILL  FILL_9562
timestamp 1677622389
transform 1 0 1816 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_605
timestamp 1677622389
transform 1 0 1824 0 -1 770
box -9 -3 26 105
use FILL  FILL_9563
timestamp 1677622389
transform 1 0 1840 0 -1 770
box -8 -3 16 105
use FILL  FILL_9564
timestamp 1677622389
transform 1 0 1848 0 -1 770
box -8 -3 16 105
use FILL  FILL_9565
timestamp 1677622389
transform 1 0 1856 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_361
timestamp 1677622389
transform 1 0 1864 0 -1 770
box -8 -3 46 105
use FILL  FILL_9566
timestamp 1677622389
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_518
timestamp 1677622389
transform -1 0 2008 0 -1 770
box -8 -3 104 105
use FILL  FILL_9567
timestamp 1677622389
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_519
timestamp 1677622389
transform -1 0 2112 0 -1 770
box -8 -3 104 105
use FILL  FILL_9568
timestamp 1677622389
transform 1 0 2112 0 -1 770
box -8 -3 16 105
use FILL  FILL_9581
timestamp 1677622389
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_520
timestamp 1677622389
transform 1 0 2128 0 -1 770
box -8 -3 104 105
use FILL  FILL_9582
timestamp 1677622389
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_521
timestamp 1677622389
transform -1 0 2328 0 -1 770
box -8 -3 104 105
use FILL  FILL_9583
timestamp 1677622389
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_9584
timestamp 1677622389
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FAX1  FAX1_20
timestamp 1677622389
transform -1 0 2464 0 -1 770
box -5 -3 126 105
use FILL  FILL_9585
timestamp 1677622389
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9586
timestamp 1677622389
transform 1 0 2472 0 -1 770
box -8 -3 16 105
use FILL  FILL_9587
timestamp 1677622389
transform 1 0 2480 0 -1 770
box -8 -3 16 105
use FILL  FILL_9588
timestamp 1677622389
transform 1 0 2488 0 -1 770
box -8 -3 16 105
use FILL  FILL_9590
timestamp 1677622389
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_9592
timestamp 1677622389
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_9597
timestamp 1677622389
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_95
timestamp 1677622389
transform 1 0 2520 0 -1 770
box -8 -3 32 105
use FILL  FILL_9598
timestamp 1677622389
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use FILL  FILL_9599
timestamp 1677622389
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_56
timestamp 1677622389
transform 1 0 2560 0 -1 770
box -8 -3 40 105
use FILL  FILL_9600
timestamp 1677622389
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7643
timestamp 1677622389
transform 1 0 2612 0 1 675
box -3 -3 3 3
use FILL  FILL_9602
timestamp 1677622389
transform 1 0 2600 0 -1 770
box -8 -3 16 105
use FILL  FILL_9610
timestamp 1677622389
transform 1 0 2608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9611
timestamp 1677622389
transform 1 0 2616 0 -1 770
box -8 -3 16 105
use FILL  FILL_9612
timestamp 1677622389
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9613
timestamp 1677622389
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9614
timestamp 1677622389
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_9615
timestamp 1677622389
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_9616
timestamp 1677622389
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use FILL  FILL_9617
timestamp 1677622389
transform 1 0 2664 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_523
timestamp 1677622389
transform -1 0 2768 0 -1 770
box -8 -3 104 105
use FILL  FILL_9618
timestamp 1677622389
transform 1 0 2768 0 -1 770
box -8 -3 16 105
use FILL  FILL_9619
timestamp 1677622389
transform 1 0 2776 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7644
timestamp 1677622389
transform 1 0 2804 0 1 675
box -3 -3 3 3
use AND2X2  AND2X2_57
timestamp 1677622389
transform -1 0 2816 0 -1 770
box -8 -3 40 105
use FILL  FILL_9620
timestamp 1677622389
transform 1 0 2816 0 -1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_4
timestamp 1677622389
transform -1 0 2880 0 -1 770
box -8 -3 64 105
use FILL  FILL_9621
timestamp 1677622389
transform 1 0 2880 0 -1 770
box -8 -3 16 105
use FILL  FILL_9622
timestamp 1677622389
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_58
timestamp 1677622389
transform -1 0 2928 0 -1 770
box -8 -3 40 105
use FILL  FILL_9623
timestamp 1677622389
transform 1 0 2928 0 -1 770
box -8 -3 16 105
use FILL  FILL_9624
timestamp 1677622389
transform 1 0 2936 0 -1 770
box -8 -3 16 105
use FILL  FILL_9625
timestamp 1677622389
transform 1 0 2944 0 -1 770
box -8 -3 16 105
use FILL  FILL_9626
timestamp 1677622389
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_9627
timestamp 1677622389
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_32
timestamp 1677622389
transform 1 0 2968 0 -1 770
box -8 -3 32 105
use FILL  FILL_9628
timestamp 1677622389
transform 1 0 2992 0 -1 770
box -8 -3 16 105
use FILL  FILL_9630
timestamp 1677622389
transform 1 0 3000 0 -1 770
box -8 -3 16 105
use FILL  FILL_9633
timestamp 1677622389
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1677622389
transform 1 0 3016 0 -1 770
box -8 -3 32 105
use FILL  FILL_9634
timestamp 1677622389
transform 1 0 3040 0 -1 770
box -8 -3 16 105
use FILL  FILL_9636
timestamp 1677622389
transform 1 0 3048 0 -1 770
box -8 -3 16 105
use FILL  FILL_9641
timestamp 1677622389
transform 1 0 3056 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_609
timestamp 1677622389
transform 1 0 3064 0 -1 770
box -9 -3 26 105
use FILL  FILL_9642
timestamp 1677622389
transform 1 0 3080 0 -1 770
box -8 -3 16 105
use FILL  FILL_9643
timestamp 1677622389
transform 1 0 3088 0 -1 770
box -8 -3 16 105
use FILL  FILL_9644
timestamp 1677622389
transform 1 0 3096 0 -1 770
box -8 -3 16 105
use FILL  FILL_9645
timestamp 1677622389
transform 1 0 3104 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1677622389
transform -1 0 3144 0 -1 770
box -8 -3 40 105
use FILL  FILL_9646
timestamp 1677622389
transform 1 0 3144 0 -1 770
box -8 -3 16 105
use FILL  FILL_9648
timestamp 1677622389
transform 1 0 3152 0 -1 770
box -8 -3 16 105
use FILL  FILL_9659
timestamp 1677622389
transform 1 0 3160 0 -1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_5
timestamp 1677622389
transform -1 0 3224 0 -1 770
box -8 -3 64 105
use FILL  FILL_9660
timestamp 1677622389
transform 1 0 3224 0 -1 770
box -8 -3 16 105
use FILL  FILL_9661
timestamp 1677622389
transform 1 0 3232 0 -1 770
box -8 -3 16 105
use FILL  FILL_9662
timestamp 1677622389
transform 1 0 3240 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_364
timestamp 1677622389
transform -1 0 3288 0 -1 770
box -8 -3 46 105
use FILL  FILL_9663
timestamp 1677622389
transform 1 0 3288 0 -1 770
box -8 -3 16 105
use FILL  FILL_9665
timestamp 1677622389
transform 1 0 3296 0 -1 770
box -8 -3 16 105
use FILL  FILL_9667
timestamp 1677622389
transform 1 0 3304 0 -1 770
box -8 -3 16 105
use FILL  FILL_9669
timestamp 1677622389
transform 1 0 3312 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7645
timestamp 1677622389
transform 1 0 3412 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_524
timestamp 1677622389
transform 1 0 3320 0 -1 770
box -8 -3 104 105
use AND2X2  AND2X2_59
timestamp 1677622389
transform 1 0 3416 0 -1 770
box -8 -3 40 105
use FILL  FILL_9675
timestamp 1677622389
transform 1 0 3448 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7646
timestamp 1677622389
transform 1 0 3468 0 1 675
box -3 -3 3 3
use FILL  FILL_9676
timestamp 1677622389
transform 1 0 3456 0 -1 770
box -8 -3 16 105
use FILL  FILL_9677
timestamp 1677622389
transform 1 0 3464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9678
timestamp 1677622389
transform 1 0 3472 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_172
timestamp 1677622389
transform 1 0 3480 0 -1 770
box -8 -3 34 105
use FILL  FILL_9679
timestamp 1677622389
transform 1 0 3512 0 -1 770
box -8 -3 16 105
use FILL  FILL_9682
timestamp 1677622389
transform 1 0 3520 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_173
timestamp 1677622389
transform 1 0 3528 0 -1 770
box -8 -3 34 105
use FILL  FILL_9683
timestamp 1677622389
transform 1 0 3560 0 -1 770
box -8 -3 16 105
use FILL  FILL_9685
timestamp 1677622389
transform 1 0 3568 0 -1 770
box -8 -3 16 105
use FILL  FILL_9687
timestamp 1677622389
transform 1 0 3576 0 -1 770
box -8 -3 16 105
use FILL  FILL_9689
timestamp 1677622389
transform 1 0 3584 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_174
timestamp 1677622389
transform 1 0 3592 0 -1 770
box -8 -3 34 105
use FILL  FILL_9691
timestamp 1677622389
transform 1 0 3624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9693
timestamp 1677622389
transform 1 0 3632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9697
timestamp 1677622389
transform 1 0 3640 0 -1 770
box -8 -3 16 105
use FILL  FILL_9698
timestamp 1677622389
transform 1 0 3648 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_363
timestamp 1677622389
transform 1 0 3656 0 -1 770
box -8 -3 46 105
use FILL  FILL_9699
timestamp 1677622389
transform 1 0 3696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9701
timestamp 1677622389
transform 1 0 3704 0 -1 770
box -8 -3 16 105
use FILL  FILL_9703
timestamp 1677622389
transform 1 0 3712 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7647
timestamp 1677622389
transform 1 0 3748 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_365
timestamp 1677622389
transform 1 0 3720 0 -1 770
box -8 -3 46 105
use FILL  FILL_9705
timestamp 1677622389
transform 1 0 3760 0 -1 770
box -8 -3 16 105
use FILL  FILL_9707
timestamp 1677622389
transform 1 0 3768 0 -1 770
box -8 -3 16 105
use FILL  FILL_9709
timestamp 1677622389
transform 1 0 3776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9711
timestamp 1677622389
transform 1 0 3784 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7648
timestamp 1677622389
transform 1 0 3804 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_366
timestamp 1677622389
transform 1 0 3792 0 -1 770
box -8 -3 46 105
use FILL  FILL_9718
timestamp 1677622389
transform 1 0 3832 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7649
timestamp 1677622389
transform 1 0 3852 0 1 675
box -3 -3 3 3
use FILL  FILL_9720
timestamp 1677622389
transform 1 0 3840 0 -1 770
box -8 -3 16 105
use FILL  FILL_9722
timestamp 1677622389
transform 1 0 3848 0 -1 770
box -8 -3 16 105
use FILL  FILL_9726
timestamp 1677622389
transform 1 0 3856 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7650
timestamp 1677622389
transform 1 0 3876 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_367
timestamp 1677622389
transform -1 0 3904 0 -1 770
box -8 -3 46 105
use FILL  FILL_9727
timestamp 1677622389
transform 1 0 3904 0 -1 770
box -8 -3 16 105
use FILL  FILL_9729
timestamp 1677622389
transform 1 0 3912 0 -1 770
box -8 -3 16 105
use FILL  FILL_9731
timestamp 1677622389
transform 1 0 3920 0 -1 770
box -8 -3 16 105
use FILL  FILL_9736
timestamp 1677622389
transform 1 0 3928 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7651
timestamp 1677622389
transform 1 0 3948 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_368
timestamp 1677622389
transform 1 0 3936 0 -1 770
box -8 -3 46 105
use FILL  FILL_9737
timestamp 1677622389
transform 1 0 3976 0 -1 770
box -8 -3 16 105
use FILL  FILL_9739
timestamp 1677622389
transform 1 0 3984 0 -1 770
box -8 -3 16 105
use FILL  FILL_9745
timestamp 1677622389
transform 1 0 3992 0 -1 770
box -8 -3 16 105
use FILL  FILL_9746
timestamp 1677622389
transform 1 0 4000 0 -1 770
box -8 -3 16 105
use FILL  FILL_9747
timestamp 1677622389
transform 1 0 4008 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7652
timestamp 1677622389
transform 1 0 4044 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_369
timestamp 1677622389
transform 1 0 4016 0 -1 770
box -8 -3 46 105
use FILL  FILL_9748
timestamp 1677622389
transform 1 0 4056 0 -1 770
box -8 -3 16 105
use FILL  FILL_9750
timestamp 1677622389
transform 1 0 4064 0 -1 770
box -8 -3 16 105
use FILL  FILL_9756
timestamp 1677622389
transform 1 0 4072 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7653
timestamp 1677622389
transform 1 0 4092 0 1 675
box -3 -3 3 3
use FILL  FILL_9757
timestamp 1677622389
transform 1 0 4080 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_370
timestamp 1677622389
transform 1 0 4088 0 -1 770
box -8 -3 46 105
use FILL  FILL_9758
timestamp 1677622389
transform 1 0 4128 0 -1 770
box -8 -3 16 105
use FILL  FILL_9760
timestamp 1677622389
transform 1 0 4136 0 -1 770
box -8 -3 16 105
use FILL  FILL_9762
timestamp 1677622389
transform 1 0 4144 0 -1 770
box -8 -3 16 105
use FILL  FILL_9764
timestamp 1677622389
transform 1 0 4152 0 -1 770
box -8 -3 16 105
use FILL  FILL_9766
timestamp 1677622389
transform 1 0 4160 0 -1 770
box -8 -3 16 105
use FILL  FILL_9767
timestamp 1677622389
transform 1 0 4168 0 -1 770
box -8 -3 16 105
use FILL  FILL_9768
timestamp 1677622389
transform 1 0 4176 0 -1 770
box -8 -3 16 105
use FILL  FILL_9769
timestamp 1677622389
transform 1 0 4184 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7654
timestamp 1677622389
transform 1 0 4204 0 1 675
box -3 -3 3 3
use FILL  FILL_9770
timestamp 1677622389
transform 1 0 4192 0 -1 770
box -8 -3 16 105
use FILL  FILL_9771
timestamp 1677622389
transform 1 0 4200 0 -1 770
box -8 -3 16 105
use FILL  FILL_9773
timestamp 1677622389
transform 1 0 4208 0 -1 770
box -8 -3 16 105
use FILL  FILL_9775
timestamp 1677622389
transform 1 0 4216 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_372
timestamp 1677622389
transform 1 0 4224 0 -1 770
box -8 -3 46 105
use FILL  FILL_9782
timestamp 1677622389
transform 1 0 4264 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7655
timestamp 1677622389
transform 1 0 4300 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_374
timestamp 1677622389
transform 1 0 4272 0 -1 770
box -8 -3 46 105
use FILL  FILL_9784
timestamp 1677622389
transform 1 0 4312 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_613
timestamp 1677622389
transform 1 0 4320 0 -1 770
box -9 -3 26 105
use M3_M2  M3_M2_7656
timestamp 1677622389
transform 1 0 4364 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_376
timestamp 1677622389
transform 1 0 4336 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_377
timestamp 1677622389
transform 1 0 4376 0 -1 770
box -8 -3 46 105
use FILL  FILL_9793
timestamp 1677622389
transform 1 0 4416 0 -1 770
box -8 -3 16 105
use FILL  FILL_9795
timestamp 1677622389
transform 1 0 4424 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7657
timestamp 1677622389
transform 1 0 4444 0 1 675
box -3 -3 3 3
use FILL  FILL_9797
timestamp 1677622389
transform 1 0 4432 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7658
timestamp 1677622389
transform 1 0 4468 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_381
timestamp 1677622389
transform 1 0 4440 0 -1 770
box -8 -3 46 105
use FILL  FILL_9815
timestamp 1677622389
transform 1 0 4480 0 -1 770
box -8 -3 16 105
use FILL  FILL_9816
timestamp 1677622389
transform 1 0 4488 0 -1 770
box -8 -3 16 105
use FILL  FILL_9817
timestamp 1677622389
transform 1 0 4496 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_382
timestamp 1677622389
transform 1 0 4504 0 -1 770
box -8 -3 46 105
use FILL  FILL_9818
timestamp 1677622389
transform 1 0 4544 0 -1 770
box -8 -3 16 105
use FILL  FILL_9819
timestamp 1677622389
transform 1 0 4552 0 -1 770
box -8 -3 16 105
use FILL  FILL_9820
timestamp 1677622389
transform 1 0 4560 0 -1 770
box -8 -3 16 105
use FILL  FILL_9821
timestamp 1677622389
transform 1 0 4568 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7659
timestamp 1677622389
transform 1 0 4604 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_383
timestamp 1677622389
transform 1 0 4576 0 -1 770
box -8 -3 46 105
use FILL  FILL_9822
timestamp 1677622389
transform 1 0 4616 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7660
timestamp 1677622389
transform 1 0 4636 0 1 675
box -3 -3 3 3
use FILL  FILL_9823
timestamp 1677622389
transform 1 0 4624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9824
timestamp 1677622389
transform 1 0 4632 0 -1 770
box -8 -3 16 105
use FILL  FILL_9825
timestamp 1677622389
transform 1 0 4640 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_384
timestamp 1677622389
transform -1 0 4688 0 -1 770
box -8 -3 46 105
use FILL  FILL_9826
timestamp 1677622389
transform 1 0 4688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9828
timestamp 1677622389
transform 1 0 4696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9837
timestamp 1677622389
transform 1 0 4704 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_385
timestamp 1677622389
transform 1 0 4712 0 -1 770
box -8 -3 46 105
use FILL  FILL_9838
timestamp 1677622389
transform 1 0 4752 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_615
timestamp 1677622389
transform -1 0 4776 0 -1 770
box -9 -3 26 105
use FILL  FILL_9839
timestamp 1677622389
transform 1 0 4776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9841
timestamp 1677622389
transform 1 0 4784 0 -1 770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_81
timestamp 1677622389
transform 1 0 4843 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_8661
timestamp 1677622389
transform 1 0 108 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7716
timestamp 1677622389
transform 1 0 164 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7665
timestamp 1677622389
transform 1 0 204 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8662
timestamp 1677622389
transform 1 0 172 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7717
timestamp 1677622389
transform 1 0 180 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8663
timestamp 1677622389
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8664
timestamp 1677622389
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8783
timestamp 1677622389
transform 1 0 172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8784
timestamp 1677622389
transform 1 0 180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8785
timestamp 1677622389
transform 1 0 196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8786
timestamp 1677622389
transform 1 0 220 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7796
timestamp 1677622389
transform 1 0 228 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8665
timestamp 1677622389
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8787
timestamp 1677622389
transform 1 0 260 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7736
timestamp 1677622389
transform 1 0 308 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7737
timestamp 1677622389
transform 1 0 348 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7669
timestamp 1677622389
transform 1 0 396 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7691
timestamp 1677622389
transform 1 0 372 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8666
timestamp 1677622389
transform 1 0 364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8667
timestamp 1677622389
transform 1 0 372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8668
timestamp 1677622389
transform 1 0 396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8788
timestamp 1677622389
transform 1 0 356 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7753
timestamp 1677622389
transform 1 0 364 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7797
timestamp 1677622389
transform 1 0 356 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7718
timestamp 1677622389
transform 1 0 404 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8789
timestamp 1677622389
transform 1 0 388 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7738
timestamp 1677622389
transform 1 0 396 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8790
timestamp 1677622389
transform 1 0 404 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7692
timestamp 1677622389
transform 1 0 516 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8669
timestamp 1677622389
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8670
timestamp 1677622389
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8671
timestamp 1677622389
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8791
timestamp 1677622389
transform 1 0 428 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7754
timestamp 1677622389
transform 1 0 412 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8792
timestamp 1677622389
transform 1 0 516 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7755
timestamp 1677622389
transform 1 0 516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7670
timestamp 1677622389
transform 1 0 548 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7674
timestamp 1677622389
transform 1 0 556 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8672
timestamp 1677622389
transform 1 0 532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8673
timestamp 1677622389
transform 1 0 556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8793
timestamp 1677622389
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8794
timestamp 1677622389
transform 1 0 564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8795
timestamp 1677622389
transform 1 0 572 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7756
timestamp 1677622389
transform 1 0 572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7798
timestamp 1677622389
transform 1 0 556 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7675
timestamp 1677622389
transform 1 0 596 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8796
timestamp 1677622389
transform 1 0 588 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7799
timestamp 1677622389
transform 1 0 588 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8674
timestamp 1677622389
transform 1 0 596 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7666
timestamp 1677622389
transform 1 0 612 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7676
timestamp 1677622389
transform 1 0 644 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8675
timestamp 1677622389
transform 1 0 612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8676
timestamp 1677622389
transform 1 0 628 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7719
timestamp 1677622389
transform 1 0 636 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8677
timestamp 1677622389
transform 1 0 644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8797
timestamp 1677622389
transform 1 0 612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8798
timestamp 1677622389
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8799
timestamp 1677622389
transform 1 0 644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7757
timestamp 1677622389
transform 1 0 604 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7758
timestamp 1677622389
transform 1 0 628 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7800
timestamp 1677622389
transform 1 0 620 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7801
timestamp 1677622389
transform 1 0 644 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8678
timestamp 1677622389
transform 1 0 684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8679
timestamp 1677622389
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8800
timestamp 1677622389
transform 1 0 692 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7759
timestamp 1677622389
transform 1 0 692 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8680
timestamp 1677622389
transform 1 0 708 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7693
timestamp 1677622389
transform 1 0 748 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7720
timestamp 1677622389
transform 1 0 740 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8681
timestamp 1677622389
transform 1 0 748 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8801
timestamp 1677622389
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8802
timestamp 1677622389
transform 1 0 740 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7671
timestamp 1677622389
transform 1 0 780 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8682
timestamp 1677622389
transform 1 0 780 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8803
timestamp 1677622389
transform 1 0 772 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7760
timestamp 1677622389
transform 1 0 772 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7667
timestamp 1677622389
transform 1 0 812 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8683
timestamp 1677622389
transform 1 0 812 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7721
timestamp 1677622389
transform 1 0 820 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8804
timestamp 1677622389
transform 1 0 820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7694
timestamp 1677622389
transform 1 0 868 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8684
timestamp 1677622389
transform 1 0 844 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7722
timestamp 1677622389
transform 1 0 852 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8685
timestamp 1677622389
transform 1 0 860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8686
timestamp 1677622389
transform 1 0 868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8805
timestamp 1677622389
transform 1 0 836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8806
timestamp 1677622389
transform 1 0 852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8807
timestamp 1677622389
transform 1 0 860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7695
timestamp 1677622389
transform 1 0 916 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8687
timestamp 1677622389
transform 1 0 884 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7723
timestamp 1677622389
transform 1 0 892 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8688
timestamp 1677622389
transform 1 0 916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8808
timestamp 1677622389
transform 1 0 964 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7802
timestamp 1677622389
transform 1 0 892 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7803
timestamp 1677622389
transform 1 0 964 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8809
timestamp 1677622389
transform 1 0 980 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8897
timestamp 1677622389
transform 1 0 980 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7739
timestamp 1677622389
transform 1 0 1004 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8898
timestamp 1677622389
transform 1 0 1004 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_8689
timestamp 1677622389
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7804
timestamp 1677622389
transform 1 0 1020 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7761
timestamp 1677622389
transform 1 0 1036 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8899
timestamp 1677622389
transform 1 0 1044 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_8690
timestamp 1677622389
transform 1 0 1068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8810
timestamp 1677622389
transform 1 0 1060 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7724
timestamp 1677622389
transform 1 0 1076 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8691
timestamp 1677622389
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8692
timestamp 1677622389
transform 1 0 1100 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7740
timestamp 1677622389
transform 1 0 1092 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8811
timestamp 1677622389
transform 1 0 1116 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7696
timestamp 1677622389
transform 1 0 1132 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8693
timestamp 1677622389
transform 1 0 1140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8812
timestamp 1677622389
transform 1 0 1132 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7668
timestamp 1677622389
transform 1 0 1148 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8694
timestamp 1677622389
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7762
timestamp 1677622389
transform 1 0 1148 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7677
timestamp 1677622389
transform 1 0 1188 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8695
timestamp 1677622389
transform 1 0 1180 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7678
timestamp 1677622389
transform 1 0 1212 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7697
timestamp 1677622389
transform 1 0 1212 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7698
timestamp 1677622389
transform 1 0 1228 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8696
timestamp 1677622389
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8697
timestamp 1677622389
transform 1 0 1228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8813
timestamp 1677622389
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8814
timestamp 1677622389
transform 1 0 1196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8815
timestamp 1677622389
transform 1 0 1220 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7763
timestamp 1677622389
transform 1 0 1220 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7699
timestamp 1677622389
transform 1 0 1308 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8698
timestamp 1677622389
transform 1 0 1284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8699
timestamp 1677622389
transform 1 0 1300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8700
timestamp 1677622389
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7741
timestamp 1677622389
transform 1 0 1284 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8816
timestamp 1677622389
transform 1 0 1292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8701
timestamp 1677622389
transform 1 0 1340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8702
timestamp 1677622389
transform 1 0 1348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8817
timestamp 1677622389
transform 1 0 1324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8818
timestamp 1677622389
transform 1 0 1332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7764
timestamp 1677622389
transform 1 0 1324 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7765
timestamp 1677622389
transform 1 0 1348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7679
timestamp 1677622389
transform 1 0 1476 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8703
timestamp 1677622389
transform 1 0 1428 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7680
timestamp 1677622389
transform 1 0 1492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7700
timestamp 1677622389
transform 1 0 1484 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8704
timestamp 1677622389
transform 1 0 1484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8705
timestamp 1677622389
transform 1 0 1492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8819
timestamp 1677622389
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8820
timestamp 1677622389
transform 1 0 1476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7766
timestamp 1677622389
transform 1 0 1460 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7701
timestamp 1677622389
transform 1 0 1532 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8706
timestamp 1677622389
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8707
timestamp 1677622389
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8821
timestamp 1677622389
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8822
timestamp 1677622389
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8708
timestamp 1677622389
transform 1 0 1612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8709
timestamp 1677622389
transform 1 0 1660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8823
timestamp 1677622389
transform 1 0 1644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7742
timestamp 1677622389
transform 1 0 1660 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7767
timestamp 1677622389
transform 1 0 1620 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7768
timestamp 1677622389
transform 1 0 1644 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8824
timestamp 1677622389
transform 1 0 1676 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7743
timestamp 1677622389
transform 1 0 1684 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7744
timestamp 1677622389
transform 1 0 1708 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7702
timestamp 1677622389
transform 1 0 1748 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7725
timestamp 1677622389
transform 1 0 1732 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8710
timestamp 1677622389
transform 1 0 1740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8711
timestamp 1677622389
transform 1 0 1756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8712
timestamp 1677622389
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8713
timestamp 1677622389
transform 1 0 1788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8825
timestamp 1677622389
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8826
timestamp 1677622389
transform 1 0 1732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8827
timestamp 1677622389
transform 1 0 1748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8828
timestamp 1677622389
transform 1 0 1764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8829
timestamp 1677622389
transform 1 0 1780 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7769
timestamp 1677622389
transform 1 0 1716 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7805
timestamp 1677622389
transform 1 0 1740 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8714
timestamp 1677622389
transform 1 0 1812 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7703
timestamp 1677622389
transform 1 0 1836 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8715
timestamp 1677622389
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8716
timestamp 1677622389
transform 1 0 1836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8830
timestamp 1677622389
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7726
timestamp 1677622389
transform 1 0 1876 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8717
timestamp 1677622389
transform 1 0 1892 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7727
timestamp 1677622389
transform 1 0 1916 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8831
timestamp 1677622389
transform 1 0 1916 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7770
timestamp 1677622389
transform 1 0 1916 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8718
timestamp 1677622389
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7681
timestamp 1677622389
transform 1 0 2052 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8719
timestamp 1677622389
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8720
timestamp 1677622389
transform 1 0 2012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8832
timestamp 1677622389
transform 1 0 1956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8833
timestamp 1677622389
transform 1 0 2044 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7771
timestamp 1677622389
transform 1 0 1964 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8721
timestamp 1677622389
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7806
timestamp 1677622389
transform 1 0 2052 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8722
timestamp 1677622389
transform 1 0 2100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8834
timestamp 1677622389
transform 1 0 2148 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8723
timestamp 1677622389
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7672
timestamp 1677622389
transform 1 0 2236 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8724
timestamp 1677622389
transform 1 0 2228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8835
timestamp 1677622389
transform 1 0 2252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8836
timestamp 1677622389
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7682
timestamp 1677622389
transform 1 0 2332 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8649
timestamp 1677622389
transform 1 0 2332 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7683
timestamp 1677622389
transform 1 0 2356 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8725
timestamp 1677622389
transform 1 0 2348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8726
timestamp 1677622389
transform 1 0 2356 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7745
timestamp 1677622389
transform 1 0 2348 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8650
timestamp 1677622389
transform 1 0 2380 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8837
timestamp 1677622389
transform 1 0 2356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8838
timestamp 1677622389
transform 1 0 2364 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7746
timestamp 1677622389
transform 1 0 2372 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7772
timestamp 1677622389
transform 1 0 2356 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7807
timestamp 1677622389
transform 1 0 2364 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7673
timestamp 1677622389
transform 1 0 2396 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8651
timestamp 1677622389
transform 1 0 2412 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8839
timestamp 1677622389
transform 1 0 2404 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7808
timestamp 1677622389
transform 1 0 2404 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8727
timestamp 1677622389
transform 1 0 2428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8728
timestamp 1677622389
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8729
timestamp 1677622389
transform 1 0 2452 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7809
timestamp 1677622389
transform 1 0 2428 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8730
timestamp 1677622389
transform 1 0 2484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8731
timestamp 1677622389
transform 1 0 2492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8840
timestamp 1677622389
transform 1 0 2468 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7773
timestamp 1677622389
transform 1 0 2476 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8900
timestamp 1677622389
transform 1 0 2484 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7810
timestamp 1677622389
transform 1 0 2492 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8732
timestamp 1677622389
transform 1 0 2524 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7704
timestamp 1677622389
transform 1 0 2540 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8841
timestamp 1677622389
transform 1 0 2540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8733
timestamp 1677622389
transform 1 0 2580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8842
timestamp 1677622389
transform 1 0 2596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8734
timestamp 1677622389
transform 1 0 2612 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7705
timestamp 1677622389
transform 1 0 2636 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8735
timestamp 1677622389
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8736
timestamp 1677622389
transform 1 0 2652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8843
timestamp 1677622389
transform 1 0 2644 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8737
timestamp 1677622389
transform 1 0 2756 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7811
timestamp 1677622389
transform 1 0 2756 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8738
timestamp 1677622389
transform 1 0 2820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8844
timestamp 1677622389
transform 1 0 2844 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7774
timestamp 1677622389
transform 1 0 2820 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8845
timestamp 1677622389
transform 1 0 2860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7775
timestamp 1677622389
transform 1 0 2860 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8739
timestamp 1677622389
transform 1 0 2876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8846
timestamp 1677622389
transform 1 0 2924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8652
timestamp 1677622389
transform 1 0 2988 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7706
timestamp 1677622389
transform 1 0 2996 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8740
timestamp 1677622389
transform 1 0 2996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8741
timestamp 1677622389
transform 1 0 3012 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7684
timestamp 1677622389
transform 1 0 3036 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8648
timestamp 1677622389
transform 1 0 3052 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_8653
timestamp 1677622389
transform 1 0 3036 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8847
timestamp 1677622389
transform 1 0 3028 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7776
timestamp 1677622389
transform 1 0 3028 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7707
timestamp 1677622389
transform 1 0 3044 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8742
timestamp 1677622389
transform 1 0 3044 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7728
timestamp 1677622389
transform 1 0 3052 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8743
timestamp 1677622389
transform 1 0 3068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8654
timestamp 1677622389
transform 1 0 3076 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7708
timestamp 1677622389
transform 1 0 3100 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8655
timestamp 1677622389
transform 1 0 3116 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7729
timestamp 1677622389
transform 1 0 3084 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8744
timestamp 1677622389
transform 1 0 3108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8848
timestamp 1677622389
transform 1 0 3100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8849
timestamp 1677622389
transform 1 0 3108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8901
timestamp 1677622389
transform 1 0 3084 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7812
timestamp 1677622389
transform 1 0 3084 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7813
timestamp 1677622389
transform 1 0 3108 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7709
timestamp 1677622389
transform 1 0 3140 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8745
timestamp 1677622389
transform 1 0 3140 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7730
timestamp 1677622389
transform 1 0 3172 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8746
timestamp 1677622389
transform 1 0 3188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8850
timestamp 1677622389
transform 1 0 3172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8851
timestamp 1677622389
transform 1 0 3180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8902
timestamp 1677622389
transform 1 0 3164 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7777
timestamp 1677622389
transform 1 0 3188 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7685
timestamp 1677622389
transform 1 0 3268 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7710
timestamp 1677622389
transform 1 0 3268 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7711
timestamp 1677622389
transform 1 0 3292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7731
timestamp 1677622389
transform 1 0 3228 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8747
timestamp 1677622389
transform 1 0 3252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8852
timestamp 1677622389
transform 1 0 3228 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7778
timestamp 1677622389
transform 1 0 3252 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7814
timestamp 1677622389
transform 1 0 3228 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7815
timestamp 1677622389
transform 1 0 3300 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8748
timestamp 1677622389
transform 1 0 3332 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7779
timestamp 1677622389
transform 1 0 3332 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8749
timestamp 1677622389
transform 1 0 3372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8853
timestamp 1677622389
transform 1 0 3348 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7816
timestamp 1677622389
transform 1 0 3348 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8854
timestamp 1677622389
transform 1 0 3452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8656
timestamp 1677622389
transform 1 0 3468 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7732
timestamp 1677622389
transform 1 0 3468 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8750
timestamp 1677622389
transform 1 0 3476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8855
timestamp 1677622389
transform 1 0 3468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8856
timestamp 1677622389
transform 1 0 3476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7780
timestamp 1677622389
transform 1 0 3460 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7686
timestamp 1677622389
transform 1 0 3508 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7733
timestamp 1677622389
transform 1 0 3500 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8657
timestamp 1677622389
transform 1 0 3524 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8751
timestamp 1677622389
transform 1 0 3508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8752
timestamp 1677622389
transform 1 0 3516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8857
timestamp 1677622389
transform 1 0 3492 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7781
timestamp 1677622389
transform 1 0 3500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7734
timestamp 1677622389
transform 1 0 3524 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8858
timestamp 1677622389
transform 1 0 3532 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7782
timestamp 1677622389
transform 1 0 3532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7687
timestamp 1677622389
transform 1 0 3548 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8658
timestamp 1677622389
transform 1 0 3548 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7712
timestamp 1677622389
transform 1 0 3564 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7735
timestamp 1677622389
transform 1 0 3556 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7688
timestamp 1677622389
transform 1 0 3580 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8659
timestamp 1677622389
transform 1 0 3580 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8753
timestamp 1677622389
transform 1 0 3564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8754
timestamp 1677622389
transform 1 0 3572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8859
timestamp 1677622389
transform 1 0 3556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7713
timestamp 1677622389
transform 1 0 3588 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8755
timestamp 1677622389
transform 1 0 3588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8860
timestamp 1677622389
transform 1 0 3596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8861
timestamp 1677622389
transform 1 0 3612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8660
timestamp 1677622389
transform 1 0 3644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8756
timestamp 1677622389
transform 1 0 3668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8757
timestamp 1677622389
transform 1 0 3700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8862
timestamp 1677622389
transform 1 0 3716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8863
timestamp 1677622389
transform 1 0 3732 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7661
timestamp 1677622389
transform 1 0 3748 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7662
timestamp 1677622389
transform 1 0 3772 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_8758
timestamp 1677622389
transform 1 0 3772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8759
timestamp 1677622389
transform 1 0 3788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8864
timestamp 1677622389
transform 1 0 3764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8865
timestamp 1677622389
transform 1 0 3780 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7817
timestamp 1677622389
transform 1 0 3764 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7818
timestamp 1677622389
transform 1 0 3788 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8866
timestamp 1677622389
transform 1 0 3820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8867
timestamp 1677622389
transform 1 0 3828 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7783
timestamp 1677622389
transform 1 0 3820 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7819
timestamp 1677622389
transform 1 0 3828 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8760
timestamp 1677622389
transform 1 0 3852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8868
timestamp 1677622389
transform 1 0 3860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8869
timestamp 1677622389
transform 1 0 3876 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7784
timestamp 1677622389
transform 1 0 3876 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8761
timestamp 1677622389
transform 1 0 3892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8762
timestamp 1677622389
transform 1 0 3948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8870
timestamp 1677622389
transform 1 0 3924 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7747
timestamp 1677622389
transform 1 0 3932 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8871
timestamp 1677622389
transform 1 0 3940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8872
timestamp 1677622389
transform 1 0 3972 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7663
timestamp 1677622389
transform 1 0 4020 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_7664
timestamp 1677622389
transform 1 0 4036 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_8763
timestamp 1677622389
transform 1 0 4012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8764
timestamp 1677622389
transform 1 0 4028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8873
timestamp 1677622389
transform 1 0 4020 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7748
timestamp 1677622389
transform 1 0 4028 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8874
timestamp 1677622389
transform 1 0 4036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8765
timestamp 1677622389
transform 1 0 4092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8766
timestamp 1677622389
transform 1 0 4108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8875
timestamp 1677622389
transform 1 0 4084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8876
timestamp 1677622389
transform 1 0 4100 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7820
timestamp 1677622389
transform 1 0 4084 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7821
timestamp 1677622389
transform 1 0 4132 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8767
timestamp 1677622389
transform 1 0 4172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8768
timestamp 1677622389
transform 1 0 4188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8877
timestamp 1677622389
transform 1 0 4156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8878
timestamp 1677622389
transform 1 0 4164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8879
timestamp 1677622389
transform 1 0 4180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8880
timestamp 1677622389
transform 1 0 4196 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7785
timestamp 1677622389
transform 1 0 4156 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7822
timestamp 1677622389
transform 1 0 4164 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7786
timestamp 1677622389
transform 1 0 4196 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8769
timestamp 1677622389
transform 1 0 4284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8881
timestamp 1677622389
transform 1 0 4236 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7749
timestamp 1677622389
transform 1 0 4308 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7787
timestamp 1677622389
transform 1 0 4284 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8770
timestamp 1677622389
transform 1 0 4324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8771
timestamp 1677622389
transform 1 0 4332 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7750
timestamp 1677622389
transform 1 0 4332 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8772
timestamp 1677622389
transform 1 0 4364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8882
timestamp 1677622389
transform 1 0 4340 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8883
timestamp 1677622389
transform 1 0 4356 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7788
timestamp 1677622389
transform 1 0 4356 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8773
timestamp 1677622389
transform 1 0 4388 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7751
timestamp 1677622389
transform 1 0 4380 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8884
timestamp 1677622389
transform 1 0 4388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8774
timestamp 1677622389
transform 1 0 4444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8885
timestamp 1677622389
transform 1 0 4420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8886
timestamp 1677622389
transform 1 0 4436 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7752
timestamp 1677622389
transform 1 0 4444 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8887
timestamp 1677622389
transform 1 0 4452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8888
timestamp 1677622389
transform 1 0 4460 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7789
timestamp 1677622389
transform 1 0 4420 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7790
timestamp 1677622389
transform 1 0 4460 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7823
timestamp 1677622389
transform 1 0 4452 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7689
timestamp 1677622389
transform 1 0 4516 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7714
timestamp 1677622389
transform 1 0 4492 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8775
timestamp 1677622389
transform 1 0 4492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8776
timestamp 1677622389
transform 1 0 4516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8889
timestamp 1677622389
transform 1 0 4508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8890
timestamp 1677622389
transform 1 0 4524 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7824
timestamp 1677622389
transform 1 0 4524 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7715
timestamp 1677622389
transform 1 0 4540 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8777
timestamp 1677622389
transform 1 0 4540 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7690
timestamp 1677622389
transform 1 0 4588 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8778
timestamp 1677622389
transform 1 0 4588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8891
timestamp 1677622389
transform 1 0 4564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8892
timestamp 1677622389
transform 1 0 4580 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7791
timestamp 1677622389
transform 1 0 4564 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7825
timestamp 1677622389
transform 1 0 4580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7826
timestamp 1677622389
transform 1 0 4612 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8779
timestamp 1677622389
transform 1 0 4636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8780
timestamp 1677622389
transform 1 0 4652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8893
timestamp 1677622389
transform 1 0 4628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8894
timestamp 1677622389
transform 1 0 4644 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8895
timestamp 1677622389
transform 1 0 4660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7792
timestamp 1677622389
transform 1 0 4660 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7827
timestamp 1677622389
transform 1 0 4644 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7793
timestamp 1677622389
transform 1 0 4684 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8781
timestamp 1677622389
transform 1 0 4732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8782
timestamp 1677622389
transform 1 0 4788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8896
timestamp 1677622389
transform 1 0 4708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7794
timestamp 1677622389
transform 1 0 4724 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7795
timestamp 1677622389
transform 1 0 4756 0 1 595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_82
timestamp 1677622389
transform 1 0 48 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_7828
timestamp 1677622389
transform 1 0 84 0 1 575
box -3 -3 3 3
use FILL  FILL_9842
timestamp 1677622389
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_9843
timestamp 1677622389
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_9844
timestamp 1677622389
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_9845
timestamp 1677622389
transform 1 0 96 0 1 570
box -8 -3 16 105
use INVX2  INVX2_616
timestamp 1677622389
transform -1 0 120 0 1 570
box -9 -3 26 105
use FILL  FILL_9846
timestamp 1677622389
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_9847
timestamp 1677622389
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_9848
timestamp 1677622389
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_9849
timestamp 1677622389
transform 1 0 144 0 1 570
box -8 -3 16 105
use FILL  FILL_9850
timestamp 1677622389
transform 1 0 152 0 1 570
box -8 -3 16 105
use FILL  FILL_9851
timestamp 1677622389
transform 1 0 160 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_366
timestamp 1677622389
transform -1 0 208 0 1 570
box -8 -3 46 105
use FILL  FILL_9852
timestamp 1677622389
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_9853
timestamp 1677622389
transform 1 0 216 0 1 570
box -8 -3 16 105
use FILL  FILL_9854
timestamp 1677622389
transform 1 0 224 0 1 570
box -8 -3 16 105
use FILL  FILL_9855
timestamp 1677622389
transform 1 0 232 0 1 570
box -8 -3 16 105
use FILL  FILL_9856
timestamp 1677622389
transform 1 0 240 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_526
timestamp 1677622389
transform 1 0 248 0 1 570
box -8 -3 104 105
use FILL  FILL_9860
timestamp 1677622389
transform 1 0 344 0 1 570
box -8 -3 16 105
use FILL  FILL_9861
timestamp 1677622389
transform 1 0 352 0 1 570
box -8 -3 16 105
use FILL  FILL_9862
timestamp 1677622389
transform 1 0 360 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_386
timestamp 1677622389
transform 1 0 368 0 1 570
box -8 -3 46 105
use FILL  FILL_9863
timestamp 1677622389
transform 1 0 408 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7829
timestamp 1677622389
transform 1 0 428 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_528
timestamp 1677622389
transform 1 0 416 0 1 570
box -8 -3 104 105
use FILL  FILL_9864
timestamp 1677622389
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_9873
timestamp 1677622389
transform 1 0 520 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7830
timestamp 1677622389
transform 1 0 548 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_387
timestamp 1677622389
transform 1 0 528 0 1 570
box -8 -3 46 105
use INVX2  INVX2_620
timestamp 1677622389
transform 1 0 568 0 1 570
box -9 -3 26 105
use FILL  FILL_9875
timestamp 1677622389
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_9876
timestamp 1677622389
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_9877
timestamp 1677622389
transform 1 0 600 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_370
timestamp 1677622389
transform 1 0 608 0 1 570
box -8 -3 46 105
use FILL  FILL_9878
timestamp 1677622389
transform 1 0 648 0 1 570
box -8 -3 16 105
use FILL  FILL_9879
timestamp 1677622389
transform 1 0 656 0 1 570
box -8 -3 16 105
use FILL  FILL_9880
timestamp 1677622389
transform 1 0 664 0 1 570
box -8 -3 16 105
use INVX2  INVX2_621
timestamp 1677622389
transform 1 0 672 0 1 570
box -9 -3 26 105
use INVX2  INVX2_622
timestamp 1677622389
transform 1 0 688 0 1 570
box -9 -3 26 105
use FILL  FILL_9881
timestamp 1677622389
transform 1 0 704 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_110
timestamp 1677622389
transform 1 0 712 0 1 570
box -5 -3 28 105
use FILL  FILL_9882
timestamp 1677622389
transform 1 0 736 0 1 570
box -8 -3 16 105
use FILL  FILL_9888
timestamp 1677622389
transform 1 0 744 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_389
timestamp 1677622389
transform 1 0 752 0 1 570
box -8 -3 46 105
use FILL  FILL_9890
timestamp 1677622389
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_9892
timestamp 1677622389
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_9894
timestamp 1677622389
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_9896
timestamp 1677622389
transform 1 0 816 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_372
timestamp 1677622389
transform 1 0 824 0 1 570
box -8 -3 46 105
use INVX2  INVX2_623
timestamp 1677622389
transform 1 0 864 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_7831
timestamp 1677622389
transform 1 0 980 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_530
timestamp 1677622389
transform -1 0 976 0 1 570
box -8 -3 104 105
use FILL  FILL_9897
timestamp 1677622389
transform 1 0 976 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_96
timestamp 1677622389
transform 1 0 984 0 1 570
box -8 -3 32 105
use FILL  FILL_9898
timestamp 1677622389
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_9899
timestamp 1677622389
transform 1 0 1016 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_99
timestamp 1677622389
transform 1 0 1024 0 1 570
box -8 -3 32 105
use FILL  FILL_9910
timestamp 1677622389
transform 1 0 1048 0 1 570
box -8 -3 16 105
use FILL  FILL_9911
timestamp 1677622389
transform 1 0 1056 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_100
timestamp 1677622389
transform 1 0 1064 0 1 570
box -8 -3 32 105
use FILL  FILL_9912
timestamp 1677622389
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_9913
timestamp 1677622389
transform 1 0 1096 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7832
timestamp 1677622389
transform 1 0 1116 0 1 575
box -3 -3 3 3
use FILL  FILL_9914
timestamp 1677622389
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_9915
timestamp 1677622389
transform 1 0 1112 0 1 570
box -8 -3 16 105
use INVX2  INVX2_624
timestamp 1677622389
transform -1 0 1136 0 1 570
box -9 -3 26 105
use INVX2  INVX2_625
timestamp 1677622389
transform -1 0 1152 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_7833
timestamp 1677622389
transform 1 0 1164 0 1 575
box -3 -3 3 3
use FILL  FILL_9916
timestamp 1677622389
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_9917
timestamp 1677622389
transform 1 0 1160 0 1 570
box -8 -3 16 105
use FILL  FILL_9918
timestamp 1677622389
transform 1 0 1168 0 1 570
box -8 -3 16 105
use FILL  FILL_9921
timestamp 1677622389
transform 1 0 1176 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7834
timestamp 1677622389
transform 1 0 1196 0 1 575
box -3 -3 3 3
use FILL  FILL_9923
timestamp 1677622389
transform 1 0 1184 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_374
timestamp 1677622389
transform 1 0 1192 0 1 570
box -8 -3 46 105
use FILL  FILL_9925
timestamp 1677622389
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_9926
timestamp 1677622389
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_9929
timestamp 1677622389
transform 1 0 1248 0 1 570
box -8 -3 16 105
use FILL  FILL_9931
timestamp 1677622389
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_9932
timestamp 1677622389
transform 1 0 1264 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7835
timestamp 1677622389
transform 1 0 1292 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_392
timestamp 1677622389
transform -1 0 1312 0 1 570
box -8 -3 46 105
use FILL  FILL_9933
timestamp 1677622389
transform 1 0 1312 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7836
timestamp 1677622389
transform 1 0 1332 0 1 575
box -3 -3 3 3
use FILL  FILL_9937
timestamp 1677622389
transform 1 0 1320 0 1 570
box -8 -3 16 105
use INVX2  INVX2_627
timestamp 1677622389
transform 1 0 1328 0 1 570
box -9 -3 26 105
use FILL  FILL_9938
timestamp 1677622389
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_9939
timestamp 1677622389
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_9940
timestamp 1677622389
transform 1 0 1360 0 1 570
box -8 -3 16 105
use FILL  FILL_9941
timestamp 1677622389
transform 1 0 1368 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_532
timestamp 1677622389
transform -1 0 1472 0 1 570
box -8 -3 104 105
use INVX2  INVX2_628
timestamp 1677622389
transform 1 0 1472 0 1 570
box -9 -3 26 105
use FILL  FILL_9942
timestamp 1677622389
transform 1 0 1488 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_376
timestamp 1677622389
transform 1 0 1496 0 1 570
box -8 -3 46 105
use FILL  FILL_9943
timestamp 1677622389
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_9960
timestamp 1677622389
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_9962
timestamp 1677622389
transform 1 0 1552 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_533
timestamp 1677622389
transform -1 0 1656 0 1 570
box -8 -3 104 105
use BUFX2  BUFX2_111
timestamp 1677622389
transform 1 0 1656 0 1 570
box -5 -3 28 105
use FILL  FILL_9963
timestamp 1677622389
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_9964
timestamp 1677622389
transform 1 0 1688 0 1 570
box -8 -3 16 105
use FILL  FILL_9965
timestamp 1677622389
transform 1 0 1696 0 1 570
box -8 -3 16 105
use FILL  FILL_9966
timestamp 1677622389
transform 1 0 1704 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_394
timestamp 1677622389
transform 1 0 1712 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_379
timestamp 1677622389
transform -1 0 1792 0 1 570
box -8 -3 46 105
use FILL  FILL_9967
timestamp 1677622389
transform 1 0 1792 0 1 570
box -8 -3 16 105
use FILL  FILL_9968
timestamp 1677622389
transform 1 0 1800 0 1 570
box -8 -3 16 105
use FILL  FILL_9969
timestamp 1677622389
transform 1 0 1808 0 1 570
box -8 -3 16 105
use INVX2  INVX2_630
timestamp 1677622389
transform 1 0 1816 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_534
timestamp 1677622389
transform -1 0 1928 0 1 570
box -8 -3 104 105
use FILL  FILL_9970
timestamp 1677622389
transform 1 0 1928 0 1 570
box -8 -3 16 105
use FILL  FILL_9971
timestamp 1677622389
transform 1 0 1936 0 1 570
box -8 -3 16 105
use INVX2  INVX2_631
timestamp 1677622389
transform -1 0 1960 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_535
timestamp 1677622389
transform -1 0 2056 0 1 570
box -8 -3 104 105
use FILL  FILL_9972
timestamp 1677622389
transform 1 0 2056 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7837
timestamp 1677622389
transform 1 0 2140 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_536
timestamp 1677622389
transform -1 0 2160 0 1 570
box -8 -3 104 105
use FILL  FILL_9973
timestamp 1677622389
transform 1 0 2160 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7838
timestamp 1677622389
transform 1 0 2180 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_537
timestamp 1677622389
transform -1 0 2264 0 1 570
box -8 -3 104 105
use FILL  FILL_9974
timestamp 1677622389
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_9975
timestamp 1677622389
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_9976
timestamp 1677622389
transform 1 0 2280 0 1 570
box -8 -3 16 105
use FILL  FILL_9977
timestamp 1677622389
transform 1 0 2288 0 1 570
box -8 -3 16 105
use FILL  FILL_9978
timestamp 1677622389
transform 1 0 2296 0 1 570
box -8 -3 16 105
use FILL  FILL_9979
timestamp 1677622389
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_9980
timestamp 1677622389
transform 1 0 2312 0 1 570
box -8 -3 16 105
use FILL  FILL_9981
timestamp 1677622389
transform 1 0 2320 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_177
timestamp 1677622389
transform -1 0 2360 0 1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_37
timestamp 1677622389
transform 1 0 2360 0 1 570
box -8 -3 32 105
use FILL  FILL_9982
timestamp 1677622389
transform 1 0 2384 0 1 570
box -8 -3 16 105
use FILL  FILL_9983
timestamp 1677622389
transform 1 0 2392 0 1 570
box -8 -3 16 105
use FILL  FILL_9984
timestamp 1677622389
transform 1 0 2400 0 1 570
box -8 -3 16 105
use FILL  FILL_9985
timestamp 1677622389
transform 1 0 2408 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7839
timestamp 1677622389
transform 1 0 2428 0 1 575
box -3 -3 3 3
use AND2X2  AND2X2_61
timestamp 1677622389
transform 1 0 2416 0 1 570
box -8 -3 40 105
use FILL  FILL_9986
timestamp 1677622389
transform 1 0 2448 0 1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_18
timestamp 1677622389
transform 1 0 2456 0 1 570
box -7 -3 39 105
use INVX2  INVX2_632
timestamp 1677622389
transform -1 0 2504 0 1 570
box -9 -3 26 105
use FILL  FILL_9987
timestamp 1677622389
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_10025
timestamp 1677622389
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_10027
timestamp 1677622389
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_10028
timestamp 1677622389
transform 1 0 2528 0 1 570
box -8 -3 16 105
use FILL  FILL_10029
timestamp 1677622389
transform 1 0 2536 0 1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_1
timestamp 1677622389
transform 1 0 2544 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_7840
timestamp 1677622389
transform 1 0 2612 0 1 575
box -3 -3 3 3
use FILL  FILL_10031
timestamp 1677622389
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_10032
timestamp 1677622389
transform 1 0 2608 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_383
timestamp 1677622389
transform 1 0 2616 0 1 570
box -8 -3 46 105
use FILL  FILL_10033
timestamp 1677622389
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_10034
timestamp 1677622389
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_10035
timestamp 1677622389
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_10036
timestamp 1677622389
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_10037
timestamp 1677622389
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_10038
timestamp 1677622389
transform 1 0 2696 0 1 570
box -8 -3 16 105
use FILL  FILL_10039
timestamp 1677622389
transform 1 0 2704 0 1 570
box -8 -3 16 105
use FILL  FILL_10040
timestamp 1677622389
transform 1 0 2712 0 1 570
box -8 -3 16 105
use FILL  FILL_10041
timestamp 1677622389
transform 1 0 2720 0 1 570
box -8 -3 16 105
use FILL  FILL_10042
timestamp 1677622389
transform 1 0 2728 0 1 570
box -8 -3 16 105
use FILL  FILL_10043
timestamp 1677622389
transform 1 0 2736 0 1 570
box -8 -3 16 105
use FILL  FILL_10044
timestamp 1677622389
transform 1 0 2744 0 1 570
box -8 -3 16 105
use FILL  FILL_10047
timestamp 1677622389
transform 1 0 2752 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_543
timestamp 1677622389
transform -1 0 2856 0 1 570
box -8 -3 104 105
use FILL  FILL_10048
timestamp 1677622389
transform 1 0 2856 0 1 570
box -8 -3 16 105
use FILL  FILL_10063
timestamp 1677622389
transform 1 0 2864 0 1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_7
timestamp 1677622389
transform 1 0 2872 0 1 570
box -8 -3 64 105
use FILL  FILL_10065
timestamp 1677622389
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_10066
timestamp 1677622389
transform 1 0 2936 0 1 570
box -8 -3 16 105
use FILL  FILL_10067
timestamp 1677622389
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_10068
timestamp 1677622389
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_10069
timestamp 1677622389
transform 1 0 2960 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_38
timestamp 1677622389
transform 1 0 2968 0 1 570
box -8 -3 32 105
use FILL  FILL_10070
timestamp 1677622389
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_10071
timestamp 1677622389
transform 1 0 3000 0 1 570
box -8 -3 16 105
use INVX2  INVX2_638
timestamp 1677622389
transform -1 0 3024 0 1 570
box -9 -3 26 105
use FILL  FILL_10072
timestamp 1677622389
transform 1 0 3024 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_74
timestamp 1677622389
transform 1 0 3032 0 1 570
box -8 -3 40 105
use M3_M2  M3_M2_7841
timestamp 1677622389
transform 1 0 3076 0 1 575
box -3 -3 3 3
use FILL  FILL_10073
timestamp 1677622389
transform 1 0 3064 0 1 570
box -8 -3 16 105
use FILL  FILL_10084
timestamp 1677622389
transform 1 0 3072 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7842
timestamp 1677622389
transform 1 0 3108 0 1 575
box -3 -3 3 3
use AOI21X1  AOI21X1_19
timestamp 1677622389
transform -1 0 3112 0 1 570
box -7 -3 39 105
use FILL  FILL_10085
timestamp 1677622389
transform 1 0 3112 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_178
timestamp 1677622389
transform -1 0 3152 0 1 570
box -8 -3 34 105
use FILL  FILL_10086
timestamp 1677622389
transform 1 0 3152 0 1 570
box -8 -3 16 105
use FILL  FILL_10087
timestamp 1677622389
transform 1 0 3160 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_103
timestamp 1677622389
transform 1 0 3168 0 1 570
box -8 -3 32 105
use FILL  FILL_10088
timestamp 1677622389
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_10098
timestamp 1677622389
transform 1 0 3200 0 1 570
box -8 -3 16 105
use FILL  FILL_10100
timestamp 1677622389
transform 1 0 3208 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_544
timestamp 1677622389
transform 1 0 3216 0 1 570
box -8 -3 104 105
use FILL  FILL_10102
timestamp 1677622389
transform 1 0 3312 0 1 570
box -8 -3 16 105
use FILL  FILL_10103
timestamp 1677622389
transform 1 0 3320 0 1 570
box -8 -3 16 105
use FILL  FILL_10104
timestamp 1677622389
transform 1 0 3328 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_545
timestamp 1677622389
transform 1 0 3336 0 1 570
box -8 -3 104 105
use FILL  FILL_10105
timestamp 1677622389
transform 1 0 3432 0 1 570
box -8 -3 16 105
use FILL  FILL_10116
timestamp 1677622389
transform 1 0 3440 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_41
timestamp 1677622389
transform 1 0 3448 0 1 570
box -8 -3 32 105
use INVX2  INVX2_640
timestamp 1677622389
transform 1 0 3472 0 1 570
box -9 -3 26 105
use FILL  FILL_10117
timestamp 1677622389
transform 1 0 3488 0 1 570
box -8 -3 16 105
use FILL  FILL_10119
timestamp 1677622389
transform 1 0 3496 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_44
timestamp 1677622389
transform 1 0 3504 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1677622389
transform 1 0 3528 0 1 570
box -8 -3 32 105
use FILL  FILL_10121
timestamp 1677622389
transform 1 0 3552 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1677622389
transform 1 0 3560 0 1 570
box -8 -3 32 105
use FILL  FILL_10122
timestamp 1677622389
transform 1 0 3584 0 1 570
box -8 -3 16 105
use FILL  FILL_10128
timestamp 1677622389
transform 1 0 3592 0 1 570
box -8 -3 16 105
use FILL  FILL_10130
timestamp 1677622389
transform 1 0 3600 0 1 570
box -8 -3 16 105
use FILL  FILL_10131
timestamp 1677622389
transform 1 0 3608 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_180
timestamp 1677622389
transform 1 0 3616 0 1 570
box -8 -3 34 105
use FILL  FILL_10132
timestamp 1677622389
transform 1 0 3648 0 1 570
box -8 -3 16 105
use FILL  FILL_10136
timestamp 1677622389
transform 1 0 3656 0 1 570
box -8 -3 16 105
use FILL  FILL_10137
timestamp 1677622389
transform 1 0 3664 0 1 570
box -8 -3 16 105
use FILL  FILL_10138
timestamp 1677622389
transform 1 0 3672 0 1 570
box -8 -3 16 105
use FILL  FILL_10139
timestamp 1677622389
transform 1 0 3680 0 1 570
box -8 -3 16 105
use FILL  FILL_10140
timestamp 1677622389
transform 1 0 3688 0 1 570
box -8 -3 16 105
use FILL  FILL_10141
timestamp 1677622389
transform 1 0 3696 0 1 570
box -8 -3 16 105
use FILL  FILL_10143
timestamp 1677622389
transform 1 0 3704 0 1 570
box -8 -3 16 105
use FILL  FILL_10145
timestamp 1677622389
transform 1 0 3712 0 1 570
box -8 -3 16 105
use INVX2  INVX2_642
timestamp 1677622389
transform -1 0 3736 0 1 570
box -9 -3 26 105
use FILL  FILL_10146
timestamp 1677622389
transform 1 0 3736 0 1 570
box -8 -3 16 105
use FILL  FILL_10147
timestamp 1677622389
transform 1 0 3744 0 1 570
box -8 -3 16 105
use FILL  FILL_10148
timestamp 1677622389
transform 1 0 3752 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_398
timestamp 1677622389
transform -1 0 3800 0 1 570
box -8 -3 46 105
use FILL  FILL_10149
timestamp 1677622389
transform 1 0 3800 0 1 570
box -8 -3 16 105
use FILL  FILL_10150
timestamp 1677622389
transform 1 0 3808 0 1 570
box -8 -3 16 105
use FILL  FILL_10151
timestamp 1677622389
transform 1 0 3816 0 1 570
box -8 -3 16 105
use FILL  FILL_10152
timestamp 1677622389
transform 1 0 3824 0 1 570
box -8 -3 16 105
use FILL  FILL_10156
timestamp 1677622389
transform 1 0 3832 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_399
timestamp 1677622389
transform -1 0 3880 0 1 570
box -8 -3 46 105
use FILL  FILL_10157
timestamp 1677622389
transform 1 0 3880 0 1 570
box -8 -3 16 105
use FILL  FILL_10158
timestamp 1677622389
transform 1 0 3888 0 1 570
box -8 -3 16 105
use FILL  FILL_10159
timestamp 1677622389
transform 1 0 3896 0 1 570
box -8 -3 16 105
use FILL  FILL_10164
timestamp 1677622389
transform 1 0 3904 0 1 570
box -8 -3 16 105
use FILL  FILL_10166
timestamp 1677622389
transform 1 0 3912 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_401
timestamp 1677622389
transform 1 0 3920 0 1 570
box -8 -3 46 105
use FILL  FILL_10168
timestamp 1677622389
transform 1 0 3960 0 1 570
box -8 -3 16 105
use FILL  FILL_10173
timestamp 1677622389
transform 1 0 3968 0 1 570
box -8 -3 16 105
use FILL  FILL_10174
timestamp 1677622389
transform 1 0 3976 0 1 570
box -8 -3 16 105
use FILL  FILL_10175
timestamp 1677622389
transform 1 0 3984 0 1 570
box -8 -3 16 105
use FILL  FILL_10176
timestamp 1677622389
transform 1 0 3992 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_402
timestamp 1677622389
transform -1 0 4040 0 1 570
box -8 -3 46 105
use FILL  FILL_10177
timestamp 1677622389
transform 1 0 4040 0 1 570
box -8 -3 16 105
use FILL  FILL_10181
timestamp 1677622389
transform 1 0 4048 0 1 570
box -8 -3 16 105
use FILL  FILL_10183
timestamp 1677622389
transform 1 0 4056 0 1 570
box -8 -3 16 105
use FILL  FILL_10185
timestamp 1677622389
transform 1 0 4064 0 1 570
box -8 -3 16 105
use FILL  FILL_10186
timestamp 1677622389
transform 1 0 4072 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_404
timestamp 1677622389
transform -1 0 4120 0 1 570
box -8 -3 46 105
use FILL  FILL_10187
timestamp 1677622389
transform 1 0 4120 0 1 570
box -8 -3 16 105
use FILL  FILL_10191
timestamp 1677622389
transform 1 0 4128 0 1 570
box -8 -3 16 105
use FILL  FILL_10193
timestamp 1677622389
transform 1 0 4136 0 1 570
box -8 -3 16 105
use FILL  FILL_10195
timestamp 1677622389
transform 1 0 4144 0 1 570
box -8 -3 16 105
use FILL  FILL_10196
timestamp 1677622389
transform 1 0 4152 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_406
timestamp 1677622389
transform -1 0 4200 0 1 570
box -8 -3 46 105
use FILL  FILL_10197
timestamp 1677622389
transform 1 0 4200 0 1 570
box -8 -3 16 105
use FILL  FILL_10198
timestamp 1677622389
transform 1 0 4208 0 1 570
box -8 -3 16 105
use FILL  FILL_10199
timestamp 1677622389
transform 1 0 4216 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_548
timestamp 1677622389
transform 1 0 4224 0 1 570
box -8 -3 104 105
use FILL  FILL_10200
timestamp 1677622389
transform 1 0 4320 0 1 570
box -8 -3 16 105
use FILL  FILL_10208
timestamp 1677622389
transform 1 0 4328 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_407
timestamp 1677622389
transform 1 0 4336 0 1 570
box -8 -3 46 105
use FILL  FILL_10210
timestamp 1677622389
transform 1 0 4376 0 1 570
box -8 -3 16 105
use FILL  FILL_10211
timestamp 1677622389
transform 1 0 4384 0 1 570
box -8 -3 16 105
use FILL  FILL_10214
timestamp 1677622389
transform 1 0 4392 0 1 570
box -8 -3 16 105
use FILL  FILL_10216
timestamp 1677622389
transform 1 0 4400 0 1 570
box -8 -3 16 105
use FILL  FILL_10218
timestamp 1677622389
transform 1 0 4408 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_409
timestamp 1677622389
transform 1 0 4416 0 1 570
box -8 -3 46 105
use FILL  FILL_10219
timestamp 1677622389
transform 1 0 4456 0 1 570
box -8 -3 16 105
use FILL  FILL_10222
timestamp 1677622389
transform 1 0 4464 0 1 570
box -8 -3 16 105
use FILL  FILL_10224
timestamp 1677622389
transform 1 0 4472 0 1 570
box -8 -3 16 105
use FILL  FILL_10226
timestamp 1677622389
transform 1 0 4480 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_411
timestamp 1677622389
transform 1 0 4488 0 1 570
box -8 -3 46 105
use FILL  FILL_10227
timestamp 1677622389
transform 1 0 4528 0 1 570
box -8 -3 16 105
use FILL  FILL_10230
timestamp 1677622389
transform 1 0 4536 0 1 570
box -8 -3 16 105
use FILL  FILL_10232
timestamp 1677622389
transform 1 0 4544 0 1 570
box -8 -3 16 105
use FILL  FILL_10234
timestamp 1677622389
transform 1 0 4552 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_413
timestamp 1677622389
transform 1 0 4560 0 1 570
box -8 -3 46 105
use FILL  FILL_10236
timestamp 1677622389
transform 1 0 4600 0 1 570
box -8 -3 16 105
use FILL  FILL_10237
timestamp 1677622389
transform 1 0 4608 0 1 570
box -8 -3 16 105
use FILL  FILL_10238
timestamp 1677622389
transform 1 0 4616 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_414
timestamp 1677622389
transform -1 0 4664 0 1 570
box -8 -3 46 105
use FILL  FILL_10239
timestamp 1677622389
transform 1 0 4664 0 1 570
box -8 -3 16 105
use FILL  FILL_10240
timestamp 1677622389
transform 1 0 4672 0 1 570
box -8 -3 16 105
use FILL  FILL_10247
timestamp 1677622389
transform 1 0 4680 0 1 570
box -8 -3 16 105
use FILL  FILL_10249
timestamp 1677622389
transform 1 0 4688 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_550
timestamp 1677622389
transform 1 0 4696 0 1 570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_83
timestamp 1677622389
transform 1 0 4819 0 1 570
box -10 -3 10 3
use M2_M1  M2_M1_8911
timestamp 1677622389
transform 1 0 84 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9023
timestamp 1677622389
transform 1 0 108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9024
timestamp 1677622389
transform 1 0 164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9025
timestamp 1677622389
transform 1 0 172 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7857
timestamp 1677622389
transform 1 0 188 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9026
timestamp 1677622389
transform 1 0 188 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7858
timestamp 1677622389
transform 1 0 204 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8912
timestamp 1677622389
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8913
timestamp 1677622389
transform 1 0 212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8914
timestamp 1677622389
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9027
timestamp 1677622389
transform 1 0 220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9028
timestamp 1677622389
transform 1 0 244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8915
timestamp 1677622389
transform 1 0 260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9029
timestamp 1677622389
transform 1 0 284 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7934
timestamp 1677622389
transform 1 0 332 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9030
timestamp 1677622389
transform 1 0 340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9031
timestamp 1677622389
transform 1 0 348 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7955
timestamp 1677622389
transform 1 0 244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7956
timestamp 1677622389
transform 1 0 292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7983
timestamp 1677622389
transform 1 0 236 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8000
timestamp 1677622389
transform 1 0 212 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8001
timestamp 1677622389
transform 1 0 300 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8002
timestamp 1677622389
transform 1 0 340 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7915
timestamp 1677622389
transform 1 0 380 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8916
timestamp 1677622389
transform 1 0 388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8917
timestamp 1677622389
transform 1 0 396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8918
timestamp 1677622389
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9032
timestamp 1677622389
transform 1 0 380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9033
timestamp 1677622389
transform 1 0 404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9034
timestamp 1677622389
transform 1 0 420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9035
timestamp 1677622389
transform 1 0 428 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7957
timestamp 1677622389
transform 1 0 420 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7879
timestamp 1677622389
transform 1 0 444 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8919
timestamp 1677622389
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8920
timestamp 1677622389
transform 1 0 460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8921
timestamp 1677622389
transform 1 0 468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9036
timestamp 1677622389
transform 1 0 452 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7984
timestamp 1677622389
transform 1 0 428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8003
timestamp 1677622389
transform 1 0 396 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7916
timestamp 1677622389
transform 1 0 476 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9037
timestamp 1677622389
transform 1 0 476 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7985
timestamp 1677622389
transform 1 0 476 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9038
timestamp 1677622389
transform 1 0 500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8922
timestamp 1677622389
transform 1 0 516 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7935
timestamp 1677622389
transform 1 0 516 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7880
timestamp 1677622389
transform 1 0 540 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9039
timestamp 1677622389
transform 1 0 532 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7843
timestamp 1677622389
transform 1 0 580 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7881
timestamp 1677622389
transform 1 0 564 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7859
timestamp 1677622389
transform 1 0 596 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7860
timestamp 1677622389
transform 1 0 628 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7882
timestamp 1677622389
transform 1 0 636 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7883
timestamp 1677622389
transform 1 0 732 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8923
timestamp 1677622389
transform 1 0 580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8924
timestamp 1677622389
transform 1 0 596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8925
timestamp 1677622389
transform 1 0 612 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8926
timestamp 1677622389
transform 1 0 636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8927
timestamp 1677622389
transform 1 0 652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9040
timestamp 1677622389
transform 1 0 588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9041
timestamp 1677622389
transform 1 0 604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9042
timestamp 1677622389
transform 1 0 620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9043
timestamp 1677622389
transform 1 0 636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7958
timestamp 1677622389
transform 1 0 564 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7986
timestamp 1677622389
transform 1 0 604 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7936
timestamp 1677622389
transform 1 0 652 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9044
timestamp 1677622389
transform 1 0 684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7937
timestamp 1677622389
transform 1 0 700 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7917
timestamp 1677622389
transform 1 0 748 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7884
timestamp 1677622389
transform 1 0 772 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8928
timestamp 1677622389
transform 1 0 756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8929
timestamp 1677622389
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9045
timestamp 1677622389
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9046
timestamp 1677622389
transform 1 0 740 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8004
timestamp 1677622389
transform 1 0 636 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8005
timestamp 1677622389
transform 1 0 676 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7959
timestamp 1677622389
transform 1 0 740 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9047
timestamp 1677622389
transform 1 0 780 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7960
timestamp 1677622389
transform 1 0 780 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8930
timestamp 1677622389
transform 1 0 812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9048
timestamp 1677622389
transform 1 0 804 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7861
timestamp 1677622389
transform 1 0 860 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8931
timestamp 1677622389
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8932
timestamp 1677622389
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9049
timestamp 1677622389
transform 1 0 844 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7938
timestamp 1677622389
transform 1 0 852 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7918
timestamp 1677622389
transform 1 0 868 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9050
timestamp 1677622389
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9051
timestamp 1677622389
transform 1 0 868 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7862
timestamp 1677622389
transform 1 0 900 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8933
timestamp 1677622389
transform 1 0 916 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7939
timestamp 1677622389
transform 1 0 916 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9052
timestamp 1677622389
transform 1 0 924 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7961
timestamp 1677622389
transform 1 0 924 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8903
timestamp 1677622389
transform 1 0 940 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8934
timestamp 1677622389
transform 1 0 940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8935
timestamp 1677622389
transform 1 0 948 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7987
timestamp 1677622389
transform 1 0 964 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7844
timestamp 1677622389
transform 1 0 988 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8904
timestamp 1677622389
transform 1 0 988 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_7885
timestamp 1677622389
transform 1 0 1004 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8905
timestamp 1677622389
transform 1 0 1012 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_7919
timestamp 1677622389
transform 1 0 996 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9053
timestamp 1677622389
transform 1 0 996 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7886
timestamp 1677622389
transform 1 0 1036 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8936
timestamp 1677622389
transform 1 0 1028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9054
timestamp 1677622389
transform 1 0 1036 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7863
timestamp 1677622389
transform 1 0 1092 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8937
timestamp 1677622389
transform 1 0 1052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8938
timestamp 1677622389
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8939
timestamp 1677622389
transform 1 0 1156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9055
timestamp 1677622389
transform 1 0 1052 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7940
timestamp 1677622389
transform 1 0 1068 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9056
timestamp 1677622389
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7941
timestamp 1677622389
transform 1 0 1140 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9057
timestamp 1677622389
transform 1 0 1148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9058
timestamp 1677622389
transform 1 0 1164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7962
timestamp 1677622389
transform 1 0 1156 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8940
timestamp 1677622389
transform 1 0 1196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9059
timestamp 1677622389
transform 1 0 1180 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7942
timestamp 1677622389
transform 1 0 1188 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7988
timestamp 1677622389
transform 1 0 1180 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8941
timestamp 1677622389
transform 1 0 1228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9060
timestamp 1677622389
transform 1 0 1220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9061
timestamp 1677622389
transform 1 0 1236 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7963
timestamp 1677622389
transform 1 0 1220 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7920
timestamp 1677622389
transform 1 0 1276 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8942
timestamp 1677622389
transform 1 0 1284 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7845
timestamp 1677622389
transform 1 0 1308 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8943
timestamp 1677622389
transform 1 0 1308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9062
timestamp 1677622389
transform 1 0 1276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9063
timestamp 1677622389
transform 1 0 1300 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7964
timestamp 1677622389
transform 1 0 1300 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8944
timestamp 1677622389
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7921
timestamp 1677622389
transform 1 0 1332 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8945
timestamp 1677622389
transform 1 0 1356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8946
timestamp 1677622389
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9064
timestamp 1677622389
transform 1 0 1332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9065
timestamp 1677622389
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7943
timestamp 1677622389
transform 1 0 1356 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7989
timestamp 1677622389
transform 1 0 1380 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7864
timestamp 1677622389
transform 1 0 1396 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9066
timestamp 1677622389
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8947
timestamp 1677622389
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9067
timestamp 1677622389
transform 1 0 1428 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7922
timestamp 1677622389
transform 1 0 1444 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9068
timestamp 1677622389
transform 1 0 1444 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7865
timestamp 1677622389
transform 1 0 1476 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7866
timestamp 1677622389
transform 1 0 1492 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9069
timestamp 1677622389
transform 1 0 1484 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7846
timestamp 1677622389
transform 1 0 1524 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7867
timestamp 1677622389
transform 1 0 1540 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8948
timestamp 1677622389
transform 1 0 1524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8949
timestamp 1677622389
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9070
timestamp 1677622389
transform 1 0 1516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7990
timestamp 1677622389
transform 1 0 1508 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9071
timestamp 1677622389
transform 1 0 1540 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7944
timestamp 1677622389
transform 1 0 1548 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7965
timestamp 1677622389
transform 1 0 1596 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9072
timestamp 1677622389
transform 1 0 1612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7887
timestamp 1677622389
transform 1 0 1660 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8950
timestamp 1677622389
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7923
timestamp 1677622389
transform 1 0 1652 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8951
timestamp 1677622389
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8952
timestamp 1677622389
transform 1 0 1684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8953
timestamp 1677622389
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9073
timestamp 1677622389
transform 1 0 1652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9074
timestamp 1677622389
transform 1 0 1668 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7966
timestamp 1677622389
transform 1 0 1668 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8954
timestamp 1677622389
transform 1 0 1724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8955
timestamp 1677622389
transform 1 0 1740 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7924
timestamp 1677622389
transform 1 0 1748 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9075
timestamp 1677622389
transform 1 0 1708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9076
timestamp 1677622389
transform 1 0 1716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9077
timestamp 1677622389
transform 1 0 1748 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7967
timestamp 1677622389
transform 1 0 1716 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7991
timestamp 1677622389
transform 1 0 1716 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8956
timestamp 1677622389
transform 1 0 1764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8957
timestamp 1677622389
transform 1 0 1796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8958
timestamp 1677622389
transform 1 0 1804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9078
timestamp 1677622389
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9079
timestamp 1677622389
transform 1 0 1788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9080
timestamp 1677622389
transform 1 0 1804 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7968
timestamp 1677622389
transform 1 0 1772 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7992
timestamp 1677622389
transform 1 0 1796 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8006
timestamp 1677622389
transform 1 0 1804 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8959
timestamp 1677622389
transform 1 0 1836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8960
timestamp 1677622389
transform 1 0 1852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8961
timestamp 1677622389
transform 1 0 1860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9081
timestamp 1677622389
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9082
timestamp 1677622389
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9083
timestamp 1677622389
transform 1 0 1844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9084
timestamp 1677622389
transform 1 0 1860 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7969
timestamp 1677622389
transform 1 0 1828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7970
timestamp 1677622389
transform 1 0 1860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7993
timestamp 1677622389
transform 1 0 1852 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8007
timestamp 1677622389
transform 1 0 1860 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9085
timestamp 1677622389
transform 1 0 1892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8962
timestamp 1677622389
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9086
timestamp 1677622389
transform 1 0 1924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9087
timestamp 1677622389
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8963
timestamp 1677622389
transform 1 0 1964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8964
timestamp 1677622389
transform 1 0 1972 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7945
timestamp 1677622389
transform 1 0 1948 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9088
timestamp 1677622389
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7946
timestamp 1677622389
transform 1 0 1964 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9089
timestamp 1677622389
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7971
timestamp 1677622389
transform 1 0 1972 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8011
timestamp 1677622389
transform 1 0 1972 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_7847
timestamp 1677622389
transform 1 0 1988 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_9090
timestamp 1677622389
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7848
timestamp 1677622389
transform 1 0 2044 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7849
timestamp 1677622389
transform 1 0 2076 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7888
timestamp 1677622389
transform 1 0 2124 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8965
timestamp 1677622389
transform 1 0 2124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9091
timestamp 1677622389
transform 1 0 2044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9092
timestamp 1677622389
transform 1 0 2092 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8012
timestamp 1677622389
transform 1 0 2116 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_7889
timestamp 1677622389
transform 1 0 2148 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7850
timestamp 1677622389
transform 1 0 2244 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7890
timestamp 1677622389
transform 1 0 2164 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8966
timestamp 1677622389
transform 1 0 2164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9093
timestamp 1677622389
transform 1 0 2196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9094
timestamp 1677622389
transform 1 0 2244 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7891
timestamp 1677622389
transform 1 0 2276 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7892
timestamp 1677622389
transform 1 0 2316 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8967
timestamp 1677622389
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9095
timestamp 1677622389
transform 1 0 2308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9096
timestamp 1677622389
transform 1 0 2364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9097
timestamp 1677622389
transform 1 0 2372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8906
timestamp 1677622389
transform 1 0 2412 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8968
timestamp 1677622389
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8969
timestamp 1677622389
transform 1 0 2428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9098
timestamp 1677622389
transform 1 0 2436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8970
timestamp 1677622389
transform 1 0 2492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8971
timestamp 1677622389
transform 1 0 2524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9099
timestamp 1677622389
transform 1 0 2516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7893
timestamp 1677622389
transform 1 0 2556 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8972
timestamp 1677622389
transform 1 0 2556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9100
timestamp 1677622389
transform 1 0 2604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9101
timestamp 1677622389
transform 1 0 2636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7894
timestamp 1677622389
transform 1 0 2660 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7895
timestamp 1677622389
transform 1 0 2732 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7925
timestamp 1677622389
transform 1 0 2708 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8973
timestamp 1677622389
transform 1 0 2732 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9102
timestamp 1677622389
transform 1 0 2652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9103
timestamp 1677622389
transform 1 0 2708 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7896
timestamp 1677622389
transform 1 0 2764 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7897
timestamp 1677622389
transform 1 0 2844 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7868
timestamp 1677622389
transform 1 0 2900 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8907
timestamp 1677622389
transform 1 0 2900 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8974
timestamp 1677622389
transform 1 0 2908 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7926
timestamp 1677622389
transform 1 0 2924 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7947
timestamp 1677622389
transform 1 0 2932 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9143
timestamp 1677622389
transform 1 0 2932 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8975
timestamp 1677622389
transform 1 0 2948 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7948
timestamp 1677622389
transform 1 0 2956 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9144
timestamp 1677622389
transform 1 0 2956 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7869
timestamp 1677622389
transform 1 0 2972 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8976
timestamp 1677622389
transform 1 0 2972 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9104
timestamp 1677622389
transform 1 0 2972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9145
timestamp 1677622389
transform 1 0 2996 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9146
timestamp 1677622389
transform 1 0 3012 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7972
timestamp 1677622389
transform 1 0 3020 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9151
timestamp 1677622389
transform 1 0 3020 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_8908
timestamp 1677622389
transform 1 0 3052 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_7870
timestamp 1677622389
transform 1 0 3084 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7898
timestamp 1677622389
transform 1 0 3076 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8977
timestamp 1677622389
transform 1 0 3076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8978
timestamp 1677622389
transform 1 0 3100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9105
timestamp 1677622389
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9106
timestamp 1677622389
transform 1 0 3116 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7899
timestamp 1677622389
transform 1 0 3164 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8979
timestamp 1677622389
transform 1 0 3180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8980
timestamp 1677622389
transform 1 0 3188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9107
timestamp 1677622389
transform 1 0 3172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8909
timestamp 1677622389
transform 1 0 3228 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_7900
timestamp 1677622389
transform 1 0 3236 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8910
timestamp 1677622389
transform 1 0 3244 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_7927
timestamp 1677622389
transform 1 0 3244 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8981
timestamp 1677622389
transform 1 0 3252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9108
timestamp 1677622389
transform 1 0 3244 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7973
timestamp 1677622389
transform 1 0 3252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7994
timestamp 1677622389
transform 1 0 3244 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9109
timestamp 1677622389
transform 1 0 3276 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7995
timestamp 1677622389
transform 1 0 3276 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8982
timestamp 1677622389
transform 1 0 3300 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7928
timestamp 1677622389
transform 1 0 3324 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9110
timestamp 1677622389
transform 1 0 3324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7996
timestamp 1677622389
transform 1 0 3364 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8983
timestamp 1677622389
transform 1 0 3460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9111
timestamp 1677622389
transform 1 0 3460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9147
timestamp 1677622389
transform 1 0 3468 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8008
timestamp 1677622389
transform 1 0 3460 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9148
timestamp 1677622389
transform 1 0 3484 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8984
timestamp 1677622389
transform 1 0 3500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8985
timestamp 1677622389
transform 1 0 3516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9112
timestamp 1677622389
transform 1 0 3508 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7974
timestamp 1677622389
transform 1 0 3508 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9113
timestamp 1677622389
transform 1 0 3524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9114
timestamp 1677622389
transform 1 0 3540 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7901
timestamp 1677622389
transform 1 0 3556 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8986
timestamp 1677622389
transform 1 0 3556 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7871
timestamp 1677622389
transform 1 0 3580 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7902
timestamp 1677622389
transform 1 0 3588 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8987
timestamp 1677622389
transform 1 0 3580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8988
timestamp 1677622389
transform 1 0 3588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9115
timestamp 1677622389
transform 1 0 3604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9149
timestamp 1677622389
transform 1 0 3596 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7997
timestamp 1677622389
transform 1 0 3596 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9150
timestamp 1677622389
transform 1 0 3628 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7998
timestamp 1677622389
transform 1 0 3628 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7903
timestamp 1677622389
transform 1 0 3676 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8989
timestamp 1677622389
transform 1 0 3676 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7929
timestamp 1677622389
transform 1 0 3684 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9116
timestamp 1677622389
transform 1 0 3660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9117
timestamp 1677622389
transform 1 0 3668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9118
timestamp 1677622389
transform 1 0 3684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8990
timestamp 1677622389
transform 1 0 3716 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7949
timestamp 1677622389
transform 1 0 3716 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7904
timestamp 1677622389
transform 1 0 3764 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8991
timestamp 1677622389
transform 1 0 3812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9119
timestamp 1677622389
transform 1 0 3732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9120
timestamp 1677622389
transform 1 0 3764 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7975
timestamp 1677622389
transform 1 0 3812 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7930
timestamp 1677622389
transform 1 0 3844 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7976
timestamp 1677622389
transform 1 0 3844 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8992
timestamp 1677622389
transform 1 0 3860 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7931
timestamp 1677622389
transform 1 0 3868 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8993
timestamp 1677622389
transform 1 0 3876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8994
timestamp 1677622389
transform 1 0 3892 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7950
timestamp 1677622389
transform 1 0 3860 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9121
timestamp 1677622389
transform 1 0 3868 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7951
timestamp 1677622389
transform 1 0 3892 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9122
timestamp 1677622389
transform 1 0 3900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7999
timestamp 1677622389
transform 1 0 3868 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7932
timestamp 1677622389
transform 1 0 3940 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8995
timestamp 1677622389
transform 1 0 3948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9123
timestamp 1677622389
transform 1 0 3940 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7905
timestamp 1677622389
transform 1 0 3980 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8996
timestamp 1677622389
transform 1 0 3980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8997
timestamp 1677622389
transform 1 0 3996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8998
timestamp 1677622389
transform 1 0 4012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9124
timestamp 1677622389
transform 1 0 3988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9125
timestamp 1677622389
transform 1 0 4004 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7952
timestamp 1677622389
transform 1 0 4012 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8999
timestamp 1677622389
transform 1 0 4036 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7977
timestamp 1677622389
transform 1 0 4028 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7906
timestamp 1677622389
transform 1 0 4044 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9000
timestamp 1677622389
transform 1 0 4044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9001
timestamp 1677622389
transform 1 0 4068 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7907
timestamp 1677622389
transform 1 0 4092 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9002
timestamp 1677622389
transform 1 0 4092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9003
timestamp 1677622389
transform 1 0 4108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9126
timestamp 1677622389
transform 1 0 4084 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7953
timestamp 1677622389
transform 1 0 4108 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7978
timestamp 1677622389
transform 1 0 4092 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8009
timestamp 1677622389
transform 1 0 4084 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8010
timestamp 1677622389
transform 1 0 4100 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9127
timestamp 1677622389
transform 1 0 4140 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7851
timestamp 1677622389
transform 1 0 4148 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7852
timestamp 1677622389
transform 1 0 4172 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7908
timestamp 1677622389
transform 1 0 4212 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9004
timestamp 1677622389
transform 1 0 4260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9128
timestamp 1677622389
transform 1 0 4212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9005
timestamp 1677622389
transform 1 0 4316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9129
timestamp 1677622389
transform 1 0 4324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7872
timestamp 1677622389
transform 1 0 4340 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9006
timestamp 1677622389
transform 1 0 4340 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7853
timestamp 1677622389
transform 1 0 4364 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_9007
timestamp 1677622389
transform 1 0 4364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9130
timestamp 1677622389
transform 1 0 4372 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7909
timestamp 1677622389
transform 1 0 4388 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9008
timestamp 1677622389
transform 1 0 4388 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7873
timestamp 1677622389
transform 1 0 4452 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7910
timestamp 1677622389
transform 1 0 4460 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9009
timestamp 1677622389
transform 1 0 4436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9010
timestamp 1677622389
transform 1 0 4452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9011
timestamp 1677622389
transform 1 0 4460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9131
timestamp 1677622389
transform 1 0 4428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9132
timestamp 1677622389
transform 1 0 4444 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7874
timestamp 1677622389
transform 1 0 4508 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7875
timestamp 1677622389
transform 1 0 4524 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9012
timestamp 1677622389
transform 1 0 4508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9013
timestamp 1677622389
transform 1 0 4524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9133
timestamp 1677622389
transform 1 0 4500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9134
timestamp 1677622389
transform 1 0 4532 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7854
timestamp 1677622389
transform 1 0 4564 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7911
timestamp 1677622389
transform 1 0 4572 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9014
timestamp 1677622389
transform 1 0 4564 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7855
timestamp 1677622389
transform 1 0 4596 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7876
timestamp 1677622389
transform 1 0 4588 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9135
timestamp 1677622389
transform 1 0 4564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9136
timestamp 1677622389
transform 1 0 4572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9137
timestamp 1677622389
transform 1 0 4580 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7979
timestamp 1677622389
transform 1 0 4580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7877
timestamp 1677622389
transform 1 0 4628 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7912
timestamp 1677622389
transform 1 0 4628 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9015
timestamp 1677622389
transform 1 0 4596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9016
timestamp 1677622389
transform 1 0 4612 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7933
timestamp 1677622389
transform 1 0 4620 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9017
timestamp 1677622389
transform 1 0 4628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9138
timestamp 1677622389
transform 1 0 4620 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7954
timestamp 1677622389
transform 1 0 4628 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9139
timestamp 1677622389
transform 1 0 4636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7980
timestamp 1677622389
transform 1 0 4636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7878
timestamp 1677622389
transform 1 0 4660 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9018
timestamp 1677622389
transform 1 0 4676 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7856
timestamp 1677622389
transform 1 0 4692 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_9019
timestamp 1677622389
transform 1 0 4692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9140
timestamp 1677622389
transform 1 0 4684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7981
timestamp 1677622389
transform 1 0 4684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7913
timestamp 1677622389
transform 1 0 4732 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9020
timestamp 1677622389
transform 1 0 4716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9021
timestamp 1677622389
transform 1 0 4732 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9141
timestamp 1677622389
transform 1 0 4724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9142
timestamp 1677622389
transform 1 0 4740 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7914
timestamp 1677622389
transform 1 0 4748 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7982
timestamp 1677622389
transform 1 0 4740 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9022
timestamp 1677622389
transform 1 0 4780 0 1 535
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_84
timestamp 1677622389
transform 1 0 24 0 1 470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_525
timestamp 1677622389
transform 1 0 72 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_617
timestamp 1677622389
transform -1 0 184 0 -1 570
box -9 -3 26 105
use FILL  FILL_9857
timestamp 1677622389
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_9858
timestamp 1677622389
transform 1 0 192 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_367
timestamp 1677622389
transform 1 0 200 0 -1 570
box -8 -3 46 105
use FILL  FILL_9859
timestamp 1677622389
transform 1 0 240 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_527
timestamp 1677622389
transform 1 0 248 0 -1 570
box -8 -3 104 105
use FILL  FILL_9865
timestamp 1677622389
transform 1 0 344 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_618
timestamp 1677622389
transform -1 0 368 0 -1 570
box -9 -3 26 105
use FILL  FILL_9866
timestamp 1677622389
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9867
timestamp 1677622389
transform 1 0 376 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8013
timestamp 1677622389
transform 1 0 396 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_368
timestamp 1677622389
transform 1 0 384 0 -1 570
box -8 -3 46 105
use FILL  FILL_9868
timestamp 1677622389
transform 1 0 424 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8014
timestamp 1677622389
transform 1 0 460 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_369
timestamp 1677622389
transform -1 0 472 0 -1 570
box -8 -3 46 105
use FILL  FILL_9869
timestamp 1677622389
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_9870
timestamp 1677622389
transform 1 0 480 0 -1 570
box -8 -3 16 105
use FILL  FILL_9871
timestamp 1677622389
transform 1 0 488 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_619
timestamp 1677622389
transform 1 0 496 0 -1 570
box -9 -3 26 105
use FILL  FILL_9872
timestamp 1677622389
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_9874
timestamp 1677622389
transform 1 0 520 0 -1 570
box -8 -3 16 105
use FILL  FILL_9883
timestamp 1677622389
transform 1 0 528 0 -1 570
box -8 -3 16 105
use FILL  FILL_9884
timestamp 1677622389
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_9885
timestamp 1677622389
transform 1 0 544 0 -1 570
box -8 -3 16 105
use FILL  FILL_9886
timestamp 1677622389
transform 1 0 552 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_388
timestamp 1677622389
transform 1 0 560 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_371
timestamp 1677622389
transform 1 0 600 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_529
timestamp 1677622389
transform 1 0 640 0 -1 570
box -8 -3 104 105
use FILL  FILL_9887
timestamp 1677622389
transform 1 0 736 0 -1 570
box -8 -3 16 105
use FILL  FILL_9889
timestamp 1677622389
transform 1 0 744 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_390
timestamp 1677622389
transform 1 0 752 0 -1 570
box -8 -3 46 105
use FILL  FILL_9891
timestamp 1677622389
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_9893
timestamp 1677622389
transform 1 0 800 0 -1 570
box -8 -3 16 105
use FILL  FILL_9895
timestamp 1677622389
transform 1 0 808 0 -1 570
box -8 -3 16 105
use FILL  FILL_9900
timestamp 1677622389
transform 1 0 816 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_373
timestamp 1677622389
transform -1 0 864 0 -1 570
box -8 -3 46 105
use FILL  FILL_9901
timestamp 1677622389
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_9902
timestamp 1677622389
transform 1 0 872 0 -1 570
box -8 -3 16 105
use FILL  FILL_9903
timestamp 1677622389
transform 1 0 880 0 -1 570
box -8 -3 16 105
use FILL  FILL_9904
timestamp 1677622389
transform 1 0 888 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_391
timestamp 1677622389
transform 1 0 896 0 -1 570
box -8 -3 46 105
use FILL  FILL_9905
timestamp 1677622389
transform 1 0 936 0 -1 570
box -8 -3 16 105
use FILL  FILL_9906
timestamp 1677622389
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_9907
timestamp 1677622389
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_9908
timestamp 1677622389
transform 1 0 960 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_97
timestamp 1677622389
transform 1 0 968 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1677622389
transform 1 0 992 0 -1 570
box -8 -3 32 105
use FILL  FILL_9909
timestamp 1677622389
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_9919
timestamp 1677622389
transform 1 0 1024 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8015
timestamp 1677622389
transform 1 0 1052 0 1 475
box -3 -3 3 3
use NOR2X1  NOR2X1_101
timestamp 1677622389
transform 1 0 1032 0 -1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_531
timestamp 1677622389
transform 1 0 1056 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_626
timestamp 1677622389
transform 1 0 1152 0 -1 570
box -9 -3 26 105
use FILL  FILL_9920
timestamp 1677622389
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_9922
timestamp 1677622389
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_9924
timestamp 1677622389
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use FILL  FILL_9927
timestamp 1677622389
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_375
timestamp 1677622389
transform 1 0 1200 0 -1 570
box -8 -3 46 105
use FILL  FILL_9928
timestamp 1677622389
transform 1 0 1240 0 -1 570
box -8 -3 16 105
use FILL  FILL_9930
timestamp 1677622389
transform 1 0 1248 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8016
timestamp 1677622389
transform 1 0 1268 0 1 475
box -3 -3 3 3
use FILL  FILL_9934
timestamp 1677622389
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8017
timestamp 1677622389
transform 1 0 1308 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_393
timestamp 1677622389
transform -1 0 1304 0 -1 570
box -8 -3 46 105
use FILL  FILL_9935
timestamp 1677622389
transform 1 0 1304 0 -1 570
box -8 -3 16 105
use FILL  FILL_9936
timestamp 1677622389
transform 1 0 1312 0 -1 570
box -8 -3 16 105
use FILL  FILL_9944
timestamp 1677622389
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_377
timestamp 1677622389
transform -1 0 1368 0 -1 570
box -8 -3 46 105
use FILL  FILL_9945
timestamp 1677622389
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9946
timestamp 1677622389
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_9947
timestamp 1677622389
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_629
timestamp 1677622389
transform 1 0 1392 0 -1 570
box -9 -3 26 105
use FILL  FILL_9948
timestamp 1677622389
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_9949
timestamp 1677622389
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_9950
timestamp 1677622389
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_9951
timestamp 1677622389
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_9952
timestamp 1677622389
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_9953
timestamp 1677622389
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_9954
timestamp 1677622389
transform 1 0 1456 0 -1 570
box -8 -3 16 105
use FILL  FILL_9955
timestamp 1677622389
transform 1 0 1464 0 -1 570
box -8 -3 16 105
use FILL  FILL_9956
timestamp 1677622389
transform 1 0 1472 0 -1 570
box -8 -3 16 105
use FILL  FILL_9957
timestamp 1677622389
transform 1 0 1480 0 -1 570
box -8 -3 16 105
use FILL  FILL_9958
timestamp 1677622389
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8018
timestamp 1677622389
transform 1 0 1524 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_378
timestamp 1677622389
transform -1 0 1536 0 -1 570
box -8 -3 46 105
use FILL  FILL_9959
timestamp 1677622389
transform 1 0 1536 0 -1 570
box -8 -3 16 105
use FILL  FILL_9961
timestamp 1677622389
transform 1 0 1544 0 -1 570
box -8 -3 16 105
use FILL  FILL_9988
timestamp 1677622389
transform 1 0 1552 0 -1 570
box -8 -3 16 105
use FILL  FILL_9989
timestamp 1677622389
transform 1 0 1560 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_633
timestamp 1677622389
transform 1 0 1568 0 -1 570
box -9 -3 26 105
use FILL  FILL_9990
timestamp 1677622389
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_9991
timestamp 1677622389
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_9992
timestamp 1677622389
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_9993
timestamp 1677622389
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_9994
timestamp 1677622389
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_9995
timestamp 1677622389
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_9996
timestamp 1677622389
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8019
timestamp 1677622389
transform 1 0 1668 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_8020
timestamp 1677622389
transform 1 0 1684 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_395
timestamp 1677622389
transform -1 0 1680 0 -1 570
box -8 -3 46 105
use FILL  FILL_9997
timestamp 1677622389
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_112
timestamp 1677622389
transform -1 0 1712 0 -1 570
box -5 -3 28 105
use FILL  FILL_9998
timestamp 1677622389
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_396
timestamp 1677622389
transform 1 0 1720 0 -1 570
box -8 -3 46 105
use FILL  FILL_9999
timestamp 1677622389
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_380
timestamp 1677622389
transform -1 0 1808 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_634
timestamp 1677622389
transform 1 0 1808 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_381
timestamp 1677622389
transform -1 0 1864 0 -1 570
box -8 -3 46 105
use FILL  FILL_10000
timestamp 1677622389
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use FILL  FILL_10001
timestamp 1677622389
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_10002
timestamp 1677622389
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_635
timestamp 1677622389
transform 1 0 1888 0 -1 570
box -9 -3 26 105
use FILL  FILL_10003
timestamp 1677622389
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_10004
timestamp 1677622389
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use FILL  FILL_10005
timestamp 1677622389
transform 1 0 1920 0 -1 570
box -8 -3 16 105
use FILL  FILL_10006
timestamp 1677622389
transform 1 0 1928 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_382
timestamp 1677622389
transform -1 0 1976 0 -1 570
box -8 -3 46 105
use FILL  FILL_10007
timestamp 1677622389
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8021
timestamp 1677622389
transform 1 0 1996 0 1 475
box -3 -3 3 3
use FILL  FILL_10008
timestamp 1677622389
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_636
timestamp 1677622389
transform 1 0 1992 0 -1 570
box -9 -3 26 105
use FILL  FILL_10009
timestamp 1677622389
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_10010
timestamp 1677622389
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use FILL  FILL_10011
timestamp 1677622389
transform 1 0 2024 0 -1 570
box -8 -3 16 105
use FILL  FILL_10012
timestamp 1677622389
transform 1 0 2032 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_538
timestamp 1677622389
transform -1 0 2136 0 -1 570
box -8 -3 104 105
use FILL  FILL_10013
timestamp 1677622389
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_10014
timestamp 1677622389
transform 1 0 2144 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_539
timestamp 1677622389
transform 1 0 2152 0 -1 570
box -8 -3 104 105
use FILL  FILL_10015
timestamp 1677622389
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_10016
timestamp 1677622389
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_540
timestamp 1677622389
transform 1 0 2264 0 -1 570
box -8 -3 104 105
use FILL  FILL_10017
timestamp 1677622389
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_10018
timestamp 1677622389
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_10019
timestamp 1677622389
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use OR2X1  OR2X1_1
timestamp 1677622389
transform -1 0 2416 0 -1 570
box -8 -3 40 105
use FILL  FILL_10020
timestamp 1677622389
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_10021
timestamp 1677622389
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_10022
timestamp 1677622389
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_6
timestamp 1677622389
transform -1 0 2496 0 -1 570
box -8 -3 64 105
use FILL  FILL_10023
timestamp 1677622389
transform 1 0 2496 0 -1 570
box -8 -3 16 105
use FILL  FILL_10024
timestamp 1677622389
transform 1 0 2504 0 -1 570
box -8 -3 16 105
use FILL  FILL_10026
timestamp 1677622389
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_637
timestamp 1677622389
transform 1 0 2520 0 -1 570
box -9 -3 26 105
use FILL  FILL_10030
timestamp 1677622389
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_541
timestamp 1677622389
transform 1 0 2544 0 -1 570
box -8 -3 104 105
use FILL  FILL_10045
timestamp 1677622389
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_542
timestamp 1677622389
transform -1 0 2744 0 -1 570
box -8 -3 104 105
use FILL  FILL_10046
timestamp 1677622389
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use FILL  FILL_10049
timestamp 1677622389
transform 1 0 2752 0 -1 570
box -8 -3 16 105
use FILL  FILL_10050
timestamp 1677622389
transform 1 0 2760 0 -1 570
box -8 -3 16 105
use FILL  FILL_10051
timestamp 1677622389
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use FILL  FILL_10052
timestamp 1677622389
transform 1 0 2776 0 -1 570
box -8 -3 16 105
use FILL  FILL_10053
timestamp 1677622389
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use FILL  FILL_10054
timestamp 1677622389
transform 1 0 2792 0 -1 570
box -8 -3 16 105
use FILL  FILL_10055
timestamp 1677622389
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use FILL  FILL_10056
timestamp 1677622389
transform 1 0 2808 0 -1 570
box -8 -3 16 105
use FILL  FILL_10057
timestamp 1677622389
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_10058
timestamp 1677622389
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_10059
timestamp 1677622389
transform 1 0 2832 0 -1 570
box -8 -3 16 105
use FILL  FILL_10060
timestamp 1677622389
transform 1 0 2840 0 -1 570
box -8 -3 16 105
use FILL  FILL_10061
timestamp 1677622389
transform 1 0 2848 0 -1 570
box -8 -3 16 105
use FILL  FILL_10062
timestamp 1677622389
transform 1 0 2856 0 -1 570
box -8 -3 16 105
use FILL  FILL_10064
timestamp 1677622389
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_10074
timestamp 1677622389
transform 1 0 2872 0 -1 570
box -8 -3 16 105
use FILL  FILL_10075
timestamp 1677622389
transform 1 0 2880 0 -1 570
box -8 -3 16 105
use FILL  FILL_10076
timestamp 1677622389
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_102
timestamp 1677622389
transform 1 0 2896 0 -1 570
box -8 -3 32 105
use FILL  FILL_10077
timestamp 1677622389
transform 1 0 2920 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_39
timestamp 1677622389
transform -1 0 2952 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1677622389
transform -1 0 2976 0 -1 570
box -8 -3 32 105
use FILL  FILL_10078
timestamp 1677622389
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_10079
timestamp 1677622389
transform 1 0 2984 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_75
timestamp 1677622389
transform -1 0 3024 0 -1 570
box -8 -3 40 105
use INVX2  INVX2_639
timestamp 1677622389
transform -1 0 3040 0 -1 570
box -9 -3 26 105
use FILL  FILL_10080
timestamp 1677622389
transform 1 0 3040 0 -1 570
box -8 -3 16 105
use FILL  FILL_10081
timestamp 1677622389
transform 1 0 3048 0 -1 570
box -8 -3 16 105
use FILL  FILL_10082
timestamp 1677622389
transform 1 0 3056 0 -1 570
box -8 -3 16 105
use FILL  FILL_10083
timestamp 1677622389
transform 1 0 3064 0 -1 570
box -8 -3 16 105
use FILL  FILL_10089
timestamp 1677622389
transform 1 0 3072 0 -1 570
box -8 -3 16 105
use FILL  FILL_10090
timestamp 1677622389
transform 1 0 3080 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_104
timestamp 1677622389
transform 1 0 3088 0 -1 570
box -8 -3 32 105
use FILL  FILL_10091
timestamp 1677622389
transform 1 0 3112 0 -1 570
box -8 -3 16 105
use FILL  FILL_10092
timestamp 1677622389
transform 1 0 3120 0 -1 570
box -8 -3 16 105
use FILL  FILL_10093
timestamp 1677622389
transform 1 0 3128 0 -1 570
box -8 -3 16 105
use FILL  FILL_10094
timestamp 1677622389
transform 1 0 3136 0 -1 570
box -8 -3 16 105
use FILL  FILL_10095
timestamp 1677622389
transform 1 0 3144 0 -1 570
box -8 -3 16 105
use AND2X2  AND2X2_62
timestamp 1677622389
transform -1 0 3184 0 -1 570
box -8 -3 40 105
use FILL  FILL_10096
timestamp 1677622389
transform 1 0 3184 0 -1 570
box -8 -3 16 105
use FILL  FILL_10097
timestamp 1677622389
transform 1 0 3192 0 -1 570
box -8 -3 16 105
use FILL  FILL_10099
timestamp 1677622389
transform 1 0 3200 0 -1 570
box -8 -3 16 105
use FILL  FILL_10101
timestamp 1677622389
transform 1 0 3208 0 -1 570
box -8 -3 16 105
use FILL  FILL_10106
timestamp 1677622389
transform 1 0 3216 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_105
timestamp 1677622389
transform 1 0 3224 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1677622389
transform 1 0 3248 0 -1 570
box -8 -3 32 105
use FILL  FILL_10107
timestamp 1677622389
transform 1 0 3272 0 -1 570
box -8 -3 16 105
use FILL  FILL_10108
timestamp 1677622389
transform 1 0 3280 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_546
timestamp 1677622389
transform 1 0 3288 0 -1 570
box -8 -3 104 105
use FILL  FILL_10109
timestamp 1677622389
transform 1 0 3384 0 -1 570
box -8 -3 16 105
use FILL  FILL_10110
timestamp 1677622389
transform 1 0 3392 0 -1 570
box -8 -3 16 105
use FILL  FILL_10111
timestamp 1677622389
transform 1 0 3400 0 -1 570
box -8 -3 16 105
use FILL  FILL_10112
timestamp 1677622389
transform 1 0 3408 0 -1 570
box -8 -3 16 105
use FILL  FILL_10113
timestamp 1677622389
transform 1 0 3416 0 -1 570
box -8 -3 16 105
use FILL  FILL_10114
timestamp 1677622389
transform 1 0 3424 0 -1 570
box -8 -3 16 105
use FILL  FILL_10115
timestamp 1677622389
transform 1 0 3432 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_42
timestamp 1677622389
transform 1 0 3440 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1677622389
transform 1 0 3464 0 -1 570
box -8 -3 32 105
use FILL  FILL_10118
timestamp 1677622389
transform 1 0 3488 0 -1 570
box -8 -3 16 105
use FILL  FILL_10120
timestamp 1677622389
transform 1 0 3496 0 -1 570
box -8 -3 16 105
use FILL  FILL_10123
timestamp 1677622389
transform 1 0 3504 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_641
timestamp 1677622389
transform 1 0 3512 0 -1 570
box -9 -3 26 105
use FILL  FILL_10124
timestamp 1677622389
transform 1 0 3528 0 -1 570
box -8 -3 16 105
use FILL  FILL_10125
timestamp 1677622389
transform 1 0 3536 0 -1 570
box -8 -3 16 105
use FILL  FILL_10126
timestamp 1677622389
transform 1 0 3544 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_179
timestamp 1677622389
transform 1 0 3552 0 -1 570
box -8 -3 34 105
use FILL  FILL_10127
timestamp 1677622389
transform 1 0 3584 0 -1 570
box -8 -3 16 105
use FILL  FILL_10129
timestamp 1677622389
transform 1 0 3592 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_181
timestamp 1677622389
transform 1 0 3600 0 -1 570
box -8 -3 34 105
use FILL  FILL_10133
timestamp 1677622389
transform 1 0 3632 0 -1 570
box -8 -3 16 105
use FILL  FILL_10134
timestamp 1677622389
transform 1 0 3640 0 -1 570
box -8 -3 16 105
use FILL  FILL_10135
timestamp 1677622389
transform 1 0 3648 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_397
timestamp 1677622389
transform 1 0 3656 0 -1 570
box -8 -3 46 105
use FILL  FILL_10142
timestamp 1677622389
transform 1 0 3696 0 -1 570
box -8 -3 16 105
use FILL  FILL_10144
timestamp 1677622389
transform 1 0 3704 0 -1 570
box -8 -3 16 105
use FILL  FILL_10153
timestamp 1677622389
transform 1 0 3712 0 -1 570
box -8 -3 16 105
use FILL  FILL_10154
timestamp 1677622389
transform 1 0 3720 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_547
timestamp 1677622389
transform -1 0 3824 0 -1 570
box -8 -3 104 105
use FILL  FILL_10155
timestamp 1677622389
transform 1 0 3824 0 -1 570
box -8 -3 16 105
use FILL  FILL_10160
timestamp 1677622389
transform 1 0 3832 0 -1 570
box -8 -3 16 105
use FILL  FILL_10161
timestamp 1677622389
transform 1 0 3840 0 -1 570
box -8 -3 16 105
use FILL  FILL_10162
timestamp 1677622389
transform 1 0 3848 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_400
timestamp 1677622389
transform -1 0 3896 0 -1 570
box -8 -3 46 105
use FILL  FILL_10163
timestamp 1677622389
transform 1 0 3896 0 -1 570
box -8 -3 16 105
use FILL  FILL_10165
timestamp 1677622389
transform 1 0 3904 0 -1 570
box -8 -3 16 105
use FILL  FILL_10167
timestamp 1677622389
transform 1 0 3912 0 -1 570
box -8 -3 16 105
use FILL  FILL_10169
timestamp 1677622389
transform 1 0 3920 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_643
timestamp 1677622389
transform -1 0 3944 0 -1 570
box -9 -3 26 105
use FILL  FILL_10170
timestamp 1677622389
transform 1 0 3944 0 -1 570
box -8 -3 16 105
use FILL  FILL_10171
timestamp 1677622389
transform 1 0 3952 0 -1 570
box -8 -3 16 105
use FILL  FILL_10172
timestamp 1677622389
transform 1 0 3960 0 -1 570
box -8 -3 16 105
use FILL  FILL_10178
timestamp 1677622389
transform 1 0 3968 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_403
timestamp 1677622389
transform -1 0 4016 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_644
timestamp 1677622389
transform -1 0 4032 0 -1 570
box -9 -3 26 105
use FILL  FILL_10179
timestamp 1677622389
transform 1 0 4032 0 -1 570
box -8 -3 16 105
use FILL  FILL_10180
timestamp 1677622389
transform 1 0 4040 0 -1 570
box -8 -3 16 105
use FILL  FILL_10182
timestamp 1677622389
transform 1 0 4048 0 -1 570
box -8 -3 16 105
use FILL  FILL_10184
timestamp 1677622389
transform 1 0 4056 0 -1 570
box -8 -3 16 105
use FILL  FILL_10188
timestamp 1677622389
transform 1 0 4064 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_405
timestamp 1677622389
transform -1 0 4112 0 -1 570
box -8 -3 46 105
use FILL  FILL_10189
timestamp 1677622389
transform 1 0 4112 0 -1 570
box -8 -3 16 105
use FILL  FILL_10190
timestamp 1677622389
transform 1 0 4120 0 -1 570
box -8 -3 16 105
use FILL  FILL_10192
timestamp 1677622389
transform 1 0 4128 0 -1 570
box -8 -3 16 105
use FILL  FILL_10194
timestamp 1677622389
transform 1 0 4136 0 -1 570
box -8 -3 16 105
use FILL  FILL_10201
timestamp 1677622389
transform 1 0 4144 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_645
timestamp 1677622389
transform -1 0 4168 0 -1 570
box -9 -3 26 105
use FILL  FILL_10202
timestamp 1677622389
transform 1 0 4168 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_549
timestamp 1677622389
transform -1 0 4272 0 -1 570
box -8 -3 104 105
use FILL  FILL_10203
timestamp 1677622389
transform 1 0 4272 0 -1 570
box -8 -3 16 105
use FILL  FILL_10204
timestamp 1677622389
transform 1 0 4280 0 -1 570
box -8 -3 16 105
use FILL  FILL_10205
timestamp 1677622389
transform 1 0 4288 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_646
timestamp 1677622389
transform -1 0 4312 0 -1 570
box -9 -3 26 105
use FILL  FILL_10206
timestamp 1677622389
transform 1 0 4312 0 -1 570
box -8 -3 16 105
use FILL  FILL_10207
timestamp 1677622389
transform 1 0 4320 0 -1 570
box -8 -3 16 105
use FILL  FILL_10209
timestamp 1677622389
transform 1 0 4328 0 -1 570
box -8 -3 16 105
use FILL  FILL_10212
timestamp 1677622389
transform 1 0 4336 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_408
timestamp 1677622389
transform 1 0 4344 0 -1 570
box -8 -3 46 105
use FILL  FILL_10213
timestamp 1677622389
transform 1 0 4384 0 -1 570
box -8 -3 16 105
use FILL  FILL_10215
timestamp 1677622389
transform 1 0 4392 0 -1 570
box -8 -3 16 105
use FILL  FILL_10217
timestamp 1677622389
transform 1 0 4400 0 -1 570
box -8 -3 16 105
use FILL  FILL_10220
timestamp 1677622389
transform 1 0 4408 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_410
timestamp 1677622389
transform -1 0 4456 0 -1 570
box -8 -3 46 105
use FILL  FILL_10221
timestamp 1677622389
transform 1 0 4456 0 -1 570
box -8 -3 16 105
use FILL  FILL_10223
timestamp 1677622389
transform 1 0 4464 0 -1 570
box -8 -3 16 105
use FILL  FILL_10225
timestamp 1677622389
transform 1 0 4472 0 -1 570
box -8 -3 16 105
use FILL  FILL_10228
timestamp 1677622389
transform 1 0 4480 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_412
timestamp 1677622389
transform -1 0 4528 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_8022
timestamp 1677622389
transform 1 0 4540 0 1 475
box -3 -3 3 3
use FILL  FILL_10229
timestamp 1677622389
transform 1 0 4528 0 -1 570
box -8 -3 16 105
use FILL  FILL_10231
timestamp 1677622389
transform 1 0 4536 0 -1 570
box -8 -3 16 105
use FILL  FILL_10233
timestamp 1677622389
transform 1 0 4544 0 -1 570
box -8 -3 16 105
use FILL  FILL_10235
timestamp 1677622389
transform 1 0 4552 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_647
timestamp 1677622389
transform 1 0 4560 0 -1 570
box -9 -3 26 105
use FILL  FILL_10241
timestamp 1677622389
transform 1 0 4576 0 -1 570
box -8 -3 16 105
use FILL  FILL_10242
timestamp 1677622389
transform 1 0 4584 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8023
timestamp 1677622389
transform 1 0 4620 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_415
timestamp 1677622389
transform 1 0 4592 0 -1 570
box -8 -3 46 105
use FILL  FILL_10243
timestamp 1677622389
transform 1 0 4632 0 -1 570
box -8 -3 16 105
use FILL  FILL_10244
timestamp 1677622389
transform 1 0 4640 0 -1 570
box -8 -3 16 105
use FILL  FILL_10245
timestamp 1677622389
transform 1 0 4648 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_648
timestamp 1677622389
transform -1 0 4672 0 -1 570
box -9 -3 26 105
use FILL  FILL_10246
timestamp 1677622389
transform 1 0 4672 0 -1 570
box -8 -3 16 105
use FILL  FILL_10248
timestamp 1677622389
transform 1 0 4680 0 -1 570
box -8 -3 16 105
use FILL  FILL_10250
timestamp 1677622389
transform 1 0 4688 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_416
timestamp 1677622389
transform 1 0 4696 0 -1 570
box -8 -3 46 105
use FILL  FILL_10251
timestamp 1677622389
transform 1 0 4736 0 -1 570
box -8 -3 16 105
use FILL  FILL_10252
timestamp 1677622389
transform 1 0 4744 0 -1 570
box -8 -3 16 105
use FILL  FILL_10253
timestamp 1677622389
transform 1 0 4752 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_649
timestamp 1677622389
transform -1 0 4776 0 -1 570
box -9 -3 26 105
use FILL  FILL_10254
timestamp 1677622389
transform 1 0 4776 0 -1 570
box -8 -3 16 105
use FILL  FILL_10255
timestamp 1677622389
transform 1 0 4784 0 -1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_85
timestamp 1677622389
transform 1 0 4843 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_8052
timestamp 1677622389
transform 1 0 132 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9166
timestamp 1677622389
transform 1 0 132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9280
timestamp 1677622389
transform 1 0 84 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8179
timestamp 1677622389
transform 1 0 84 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8053
timestamp 1677622389
transform 1 0 172 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8132
timestamp 1677622389
transform 1 0 172 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8054
timestamp 1677622389
transform 1 0 196 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9167
timestamp 1677622389
transform 1 0 196 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8055
timestamp 1677622389
transform 1 0 228 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8096
timestamp 1677622389
transform 1 0 212 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9168
timestamp 1677622389
transform 1 0 220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9169
timestamp 1677622389
transform 1 0 236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9281
timestamp 1677622389
transform 1 0 204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9282
timestamp 1677622389
transform 1 0 212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9283
timestamp 1677622389
transform 1 0 228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8133
timestamp 1677622389
transform 1 0 228 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8180
timestamp 1677622389
transform 1 0 252 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8056
timestamp 1677622389
transform 1 0 276 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9170
timestamp 1677622389
transform 1 0 284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9171
timestamp 1677622389
transform 1 0 292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9284
timestamp 1677622389
transform 1 0 276 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8057
timestamp 1677622389
transform 1 0 332 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9172
timestamp 1677622389
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9285
timestamp 1677622389
transform 1 0 324 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9286
timestamp 1677622389
transform 1 0 340 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8041
timestamp 1677622389
transform 1 0 388 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9173
timestamp 1677622389
transform 1 0 388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9287
timestamp 1677622389
transform 1 0 380 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8097
timestamp 1677622389
transform 1 0 396 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9174
timestamp 1677622389
transform 1 0 404 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8098
timestamp 1677622389
transform 1 0 412 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9288
timestamp 1677622389
transform 1 0 396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9289
timestamp 1677622389
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9290
timestamp 1677622389
transform 1 0 420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9175
timestamp 1677622389
transform 1 0 436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9176
timestamp 1677622389
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9177
timestamp 1677622389
transform 1 0 500 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8099
timestamp 1677622389
transform 1 0 532 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9178
timestamp 1677622389
transform 1 0 540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9291
timestamp 1677622389
transform 1 0 460 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8134
timestamp 1677622389
transform 1 0 444 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8135
timestamp 1677622389
transform 1 0 476 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9292
timestamp 1677622389
transform 1 0 548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9179
timestamp 1677622389
transform 1 0 564 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8058
timestamp 1677622389
transform 1 0 596 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9180
timestamp 1677622389
transform 1 0 596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9293
timestamp 1677622389
transform 1 0 588 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8121
timestamp 1677622389
transform 1 0 596 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9181
timestamp 1677622389
transform 1 0 612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9294
timestamp 1677622389
transform 1 0 604 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8181
timestamp 1677622389
transform 1 0 588 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8042
timestamp 1677622389
transform 1 0 620 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9182
timestamp 1677622389
transform 1 0 620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9183
timestamp 1677622389
transform 1 0 660 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8100
timestamp 1677622389
transform 1 0 668 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9184
timestamp 1677622389
transform 1 0 676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9295
timestamp 1677622389
transform 1 0 652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9296
timestamp 1677622389
transform 1 0 668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9297
timestamp 1677622389
transform 1 0 676 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8059
timestamp 1677622389
transform 1 0 708 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9185
timestamp 1677622389
transform 1 0 708 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8136
timestamp 1677622389
transform 1 0 700 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8060
timestamp 1677622389
transform 1 0 748 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8061
timestamp 1677622389
transform 1 0 804 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9186
timestamp 1677622389
transform 1 0 748 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8101
timestamp 1677622389
transform 1 0 756 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8102
timestamp 1677622389
transform 1 0 796 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9187
timestamp 1677622389
transform 1 0 804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9298
timestamp 1677622389
transform 1 0 724 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8137
timestamp 1677622389
transform 1 0 724 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9299
timestamp 1677622389
transform 1 0 844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8031
timestamp 1677622389
transform 1 0 860 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8043
timestamp 1677622389
transform 1 0 860 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9188
timestamp 1677622389
transform 1 0 860 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8062
timestamp 1677622389
transform 1 0 884 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9189
timestamp 1677622389
transform 1 0 884 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8103
timestamp 1677622389
transform 1 0 916 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8044
timestamp 1677622389
transform 1 0 940 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9190
timestamp 1677622389
transform 1 0 932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9191
timestamp 1677622389
transform 1 0 948 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8104
timestamp 1677622389
transform 1 0 956 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8045
timestamp 1677622389
transform 1 0 988 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8063
timestamp 1677622389
transform 1 0 980 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8064
timestamp 1677622389
transform 1 0 1020 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9192
timestamp 1677622389
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9193
timestamp 1677622389
transform 1 0 980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9194
timestamp 1677622389
transform 1 0 988 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9195
timestamp 1677622389
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9300
timestamp 1677622389
transform 1 0 940 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9301
timestamp 1677622389
transform 1 0 956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9302
timestamp 1677622389
transform 1 0 964 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9303
timestamp 1677622389
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9365
timestamp 1677622389
transform 1 0 1084 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_8182
timestamp 1677622389
transform 1 0 1084 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9196
timestamp 1677622389
transform 1 0 1124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9304
timestamp 1677622389
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8122
timestamp 1677622389
transform 1 0 1124 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9197
timestamp 1677622389
transform 1 0 1164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9305
timestamp 1677622389
transform 1 0 1140 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8138
timestamp 1677622389
transform 1 0 1140 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8139
timestamp 1677622389
transform 1 0 1188 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8183
timestamp 1677622389
transform 1 0 1132 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8032
timestamp 1677622389
transform 1 0 1236 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9198
timestamp 1677622389
transform 1 0 1228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9199
timestamp 1677622389
transform 1 0 1236 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8184
timestamp 1677622389
transform 1 0 1260 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9306
timestamp 1677622389
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8065
timestamp 1677622389
transform 1 0 1332 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9200
timestamp 1677622389
transform 1 0 1308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9201
timestamp 1677622389
transform 1 0 1324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9202
timestamp 1677622389
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9307
timestamp 1677622389
transform 1 0 1308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9308
timestamp 1677622389
transform 1 0 1332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8066
timestamp 1677622389
transform 1 0 1452 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9203
timestamp 1677622389
transform 1 0 1396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9204
timestamp 1677622389
transform 1 0 1452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9205
timestamp 1677622389
transform 1 0 1460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9309
timestamp 1677622389
transform 1 0 1372 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8140
timestamp 1677622389
transform 1 0 1372 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9310
timestamp 1677622389
transform 1 0 1516 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8067
timestamp 1677622389
transform 1 0 1604 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9206
timestamp 1677622389
transform 1 0 1548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9207
timestamp 1677622389
transform 1 0 1604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9311
timestamp 1677622389
transform 1 0 1628 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8141
timestamp 1677622389
transform 1 0 1548 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8185
timestamp 1677622389
transform 1 0 1628 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8068
timestamp 1677622389
transform 1 0 1644 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9208
timestamp 1677622389
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8123
timestamp 1677622389
transform 1 0 1644 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8069
timestamp 1677622389
transform 1 0 1660 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8142
timestamp 1677622389
transform 1 0 1652 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9209
timestamp 1677622389
transform 1 0 1668 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8124
timestamp 1677622389
transform 1 0 1668 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8070
timestamp 1677622389
transform 1 0 1700 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8105
timestamp 1677622389
transform 1 0 1692 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8046
timestamp 1677622389
transform 1 0 1724 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9210
timestamp 1677622389
transform 1 0 1700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9211
timestamp 1677622389
transform 1 0 1716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9312
timestamp 1677622389
transform 1 0 1684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9313
timestamp 1677622389
transform 1 0 1692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9314
timestamp 1677622389
transform 1 0 1708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8143
timestamp 1677622389
transform 1 0 1708 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8106
timestamp 1677622389
transform 1 0 1756 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9212
timestamp 1677622389
transform 1 0 1764 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8107
timestamp 1677622389
transform 1 0 1796 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9213
timestamp 1677622389
transform 1 0 1820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9315
timestamp 1677622389
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8186
timestamp 1677622389
transform 1 0 1844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8026
timestamp 1677622389
transform 1 0 1868 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8033
timestamp 1677622389
transform 1 0 1860 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9214
timestamp 1677622389
transform 1 0 1860 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8047
timestamp 1677622389
transform 1 0 1908 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8071
timestamp 1677622389
transform 1 0 1900 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8072
timestamp 1677622389
transform 1 0 1916 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9215
timestamp 1677622389
transform 1 0 1900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9216
timestamp 1677622389
transform 1 0 1924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9316
timestamp 1677622389
transform 1 0 1892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9317
timestamp 1677622389
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9318
timestamp 1677622389
transform 1 0 1916 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8144
timestamp 1677622389
transform 1 0 1892 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8187
timestamp 1677622389
transform 1 0 1884 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8073
timestamp 1677622389
transform 1 0 1932 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9217
timestamp 1677622389
transform 1 0 1956 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8145
timestamp 1677622389
transform 1 0 1948 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9218
timestamp 1677622389
transform 1 0 1972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9319
timestamp 1677622389
transform 1 0 1964 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8125
timestamp 1677622389
transform 1 0 1972 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8146
timestamp 1677622389
transform 1 0 1964 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8188
timestamp 1677622389
transform 1 0 1972 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8048
timestamp 1677622389
transform 1 0 2004 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8074
timestamp 1677622389
transform 1 0 2012 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9219
timestamp 1677622389
transform 1 0 1996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9220
timestamp 1677622389
transform 1 0 2012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9320
timestamp 1677622389
transform 1 0 2004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9321
timestamp 1677622389
transform 1 0 2012 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8147
timestamp 1677622389
transform 1 0 1988 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8049
timestamp 1677622389
transform 1 0 2076 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8075
timestamp 1677622389
transform 1 0 2068 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8076
timestamp 1677622389
transform 1 0 2108 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9221
timestamp 1677622389
transform 1 0 2068 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9222
timestamp 1677622389
transform 1 0 2076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9223
timestamp 1677622389
transform 1 0 2108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9322
timestamp 1677622389
transform 1 0 2156 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8148
timestamp 1677622389
transform 1 0 2156 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8027
timestamp 1677622389
transform 1 0 2172 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9224
timestamp 1677622389
transform 1 0 2172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9225
timestamp 1677622389
transform 1 0 2228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9323
timestamp 1677622389
transform 1 0 2260 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8149
timestamp 1677622389
transform 1 0 2180 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8150
timestamp 1677622389
transform 1 0 2260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8189
timestamp 1677622389
transform 1 0 2244 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8034
timestamp 1677622389
transform 1 0 2284 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9226
timestamp 1677622389
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9227
timestamp 1677622389
transform 1 0 2348 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9324
timestamp 1677622389
transform 1 0 2372 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8151
timestamp 1677622389
transform 1 0 2340 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8152
timestamp 1677622389
transform 1 0 2372 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9366
timestamp 1677622389
transform 1 0 2388 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_8190
timestamp 1677622389
transform 1 0 2372 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9228
timestamp 1677622389
transform 1 0 2404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9229
timestamp 1677622389
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9230
timestamp 1677622389
transform 1 0 2468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9325
timestamp 1677622389
transform 1 0 2436 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8153
timestamp 1677622389
transform 1 0 2436 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8154
timestamp 1677622389
transform 1 0 2468 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8191
timestamp 1677622389
transform 1 0 2508 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9231
timestamp 1677622389
transform 1 0 2524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9326
timestamp 1677622389
transform 1 0 2524 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8155
timestamp 1677622389
transform 1 0 2524 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8077
timestamp 1677622389
transform 1 0 2556 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9155
timestamp 1677622389
transform 1 0 2564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9232
timestamp 1677622389
transform 1 0 2556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9327
timestamp 1677622389
transform 1 0 2548 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8078
timestamp 1677622389
transform 1 0 2580 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8108
timestamp 1677622389
transform 1 0 2564 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9233
timestamp 1677622389
transform 1 0 2580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9328
timestamp 1677622389
transform 1 0 2588 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8156
timestamp 1677622389
transform 1 0 2588 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9156
timestamp 1677622389
transform 1 0 2604 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8109
timestamp 1677622389
transform 1 0 2604 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9152
timestamp 1677622389
transform 1 0 2628 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_9234
timestamp 1677622389
transform 1 0 2620 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8157
timestamp 1677622389
transform 1 0 2620 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9157
timestamp 1677622389
transform 1 0 2636 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8079
timestamp 1677622389
transform 1 0 2708 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9235
timestamp 1677622389
transform 1 0 2708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9329
timestamp 1677622389
transform 1 0 2660 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8158
timestamp 1677622389
transform 1 0 2660 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9236
timestamp 1677622389
transform 1 0 2748 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8080
timestamp 1677622389
transform 1 0 2788 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9237
timestamp 1677622389
transform 1 0 2788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9238
timestamp 1677622389
transform 1 0 2844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9330
timestamp 1677622389
transform 1 0 2764 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8126
timestamp 1677622389
transform 1 0 2804 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8127
timestamp 1677622389
transform 1 0 2844 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8159
timestamp 1677622389
transform 1 0 2764 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8081
timestamp 1677622389
transform 1 0 2932 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8082
timestamp 1677622389
transform 1 0 2948 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9239
timestamp 1677622389
transform 1 0 2908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9240
timestamp 1677622389
transform 1 0 2948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9331
timestamp 1677622389
transform 1 0 2868 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8160
timestamp 1677622389
transform 1 0 2868 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9241
timestamp 1677622389
transform 1 0 2972 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8083
timestamp 1677622389
transform 1 0 2996 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9332
timestamp 1677622389
transform 1 0 2988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9333
timestamp 1677622389
transform 1 0 2996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9367
timestamp 1677622389
transform 1 0 2996 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9368
timestamp 1677622389
transform 1 0 3004 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_8161
timestamp 1677622389
transform 1 0 3028 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9153
timestamp 1677622389
transform 1 0 3068 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_8084
timestamp 1677622389
transform 1 0 3068 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9158
timestamp 1677622389
transform 1 0 3076 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9159
timestamp 1677622389
transform 1 0 3084 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9160
timestamp 1677622389
transform 1 0 3100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9242
timestamp 1677622389
transform 1 0 3060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9243
timestamp 1677622389
transform 1 0 3100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9154
timestamp 1677622389
transform 1 0 3116 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_9334
timestamp 1677622389
transform 1 0 3116 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8085
timestamp 1677622389
transform 1 0 3132 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9370
timestamp 1677622389
transform 1 0 3124 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_9369
timestamp 1677622389
transform 1 0 3140 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9244
timestamp 1677622389
transform 1 0 3156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9245
timestamp 1677622389
transform 1 0 3236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9335
timestamp 1677622389
transform 1 0 3204 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8086
timestamp 1677622389
transform 1 0 3316 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9246
timestamp 1677622389
transform 1 0 3316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9247
timestamp 1677622389
transform 1 0 3364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9336
timestamp 1677622389
transform 1 0 3340 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8087
timestamp 1677622389
transform 1 0 3428 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9248
timestamp 1677622389
transform 1 0 3436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9337
timestamp 1677622389
transform 1 0 3428 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8162
timestamp 1677622389
transform 1 0 3436 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8028
timestamp 1677622389
transform 1 0 3460 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9161
timestamp 1677622389
transform 1 0 3468 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9249
timestamp 1677622389
transform 1 0 3460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9338
timestamp 1677622389
transform 1 0 3468 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8163
timestamp 1677622389
transform 1 0 3468 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9162
timestamp 1677622389
transform 1 0 3492 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9250
timestamp 1677622389
transform 1 0 3508 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8128
timestamp 1677622389
transform 1 0 3508 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9163
timestamp 1677622389
transform 1 0 3532 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8110
timestamp 1677622389
transform 1 0 3524 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9339
timestamp 1677622389
transform 1 0 3516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9251
timestamp 1677622389
transform 1 0 3540 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8164
timestamp 1677622389
transform 1 0 3532 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9164
timestamp 1677622389
transform 1 0 3556 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8111
timestamp 1677622389
transform 1 0 3556 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9165
timestamp 1677622389
transform 1 0 3572 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9252
timestamp 1677622389
transform 1 0 3564 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8112
timestamp 1677622389
transform 1 0 3572 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9340
timestamp 1677622389
transform 1 0 3572 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8165
timestamp 1677622389
transform 1 0 3572 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9253
timestamp 1677622389
transform 1 0 3604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9341
timestamp 1677622389
transform 1 0 3596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8166
timestamp 1677622389
transform 1 0 3596 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8113
timestamp 1677622389
transform 1 0 3652 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8035
timestamp 1677622389
transform 1 0 3684 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8088
timestamp 1677622389
transform 1 0 3668 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9254
timestamp 1677622389
transform 1 0 3668 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8114
timestamp 1677622389
transform 1 0 3676 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9255
timestamp 1677622389
transform 1 0 3684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9342
timestamp 1677622389
transform 1 0 3660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9343
timestamp 1677622389
transform 1 0 3676 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8167
timestamp 1677622389
transform 1 0 3660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8036
timestamp 1677622389
transform 1 0 3708 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8089
timestamp 1677622389
transform 1 0 3700 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9256
timestamp 1677622389
transform 1 0 3700 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8090
timestamp 1677622389
transform 1 0 3716 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9344
timestamp 1677622389
transform 1 0 3716 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8091
timestamp 1677622389
transform 1 0 3732 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9257
timestamp 1677622389
transform 1 0 3732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9345
timestamp 1677622389
transform 1 0 3740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8115
timestamp 1677622389
transform 1 0 3748 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9346
timestamp 1677622389
transform 1 0 3748 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8168
timestamp 1677622389
transform 1 0 3748 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9258
timestamp 1677622389
transform 1 0 3788 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8129
timestamp 1677622389
transform 1 0 3788 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9347
timestamp 1677622389
transform 1 0 3796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9348
timestamp 1677622389
transform 1 0 3812 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8169
timestamp 1677622389
transform 1 0 3812 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9259
timestamp 1677622389
transform 1 0 3828 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8116
timestamp 1677622389
transform 1 0 3844 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9260
timestamp 1677622389
transform 1 0 3876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9349
timestamp 1677622389
transform 1 0 3844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8170
timestamp 1677622389
transform 1 0 3892 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9261
timestamp 1677622389
transform 1 0 3940 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8029
timestamp 1677622389
transform 1 0 3988 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8030
timestamp 1677622389
transform 1 0 4004 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8037
timestamp 1677622389
transform 1 0 3972 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8038
timestamp 1677622389
transform 1 0 3988 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8117
timestamp 1677622389
transform 1 0 3956 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9262
timestamp 1677622389
transform 1 0 3996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9263
timestamp 1677622389
transform 1 0 4036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9350
timestamp 1677622389
transform 1 0 3956 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8118
timestamp 1677622389
transform 1 0 4060 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8050
timestamp 1677622389
transform 1 0 4076 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9264
timestamp 1677622389
transform 1 0 4076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9265
timestamp 1677622389
transform 1 0 4092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9351
timestamp 1677622389
transform 1 0 4068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9352
timestamp 1677622389
transform 1 0 4084 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8171
timestamp 1677622389
transform 1 0 4068 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8119
timestamp 1677622389
transform 1 0 4108 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9353
timestamp 1677622389
transform 1 0 4108 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8092
timestamp 1677622389
transform 1 0 4156 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8120
timestamp 1677622389
transform 1 0 4148 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9266
timestamp 1677622389
transform 1 0 4156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9267
timestamp 1677622389
transform 1 0 4172 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8093
timestamp 1677622389
transform 1 0 4188 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9268
timestamp 1677622389
transform 1 0 4188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9354
timestamp 1677622389
transform 1 0 4140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9355
timestamp 1677622389
transform 1 0 4148 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9356
timestamp 1677622389
transform 1 0 4164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9357
timestamp 1677622389
transform 1 0 4180 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8172
timestamp 1677622389
transform 1 0 4180 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9358
timestamp 1677622389
transform 1 0 4212 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8039
timestamp 1677622389
transform 1 0 4284 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9269
timestamp 1677622389
transform 1 0 4284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9270
timestamp 1677622389
transform 1 0 4316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9359
timestamp 1677622389
transform 1 0 4236 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8130
timestamp 1677622389
transform 1 0 4276 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8131
timestamp 1677622389
transform 1 0 4316 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8173
timestamp 1677622389
transform 1 0 4236 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8174
timestamp 1677622389
transform 1 0 4260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8040
timestamp 1677622389
transform 1 0 4364 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8051
timestamp 1677622389
transform 1 0 4428 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8094
timestamp 1677622389
transform 1 0 4396 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8095
timestamp 1677622389
transform 1 0 4436 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9271
timestamp 1677622389
transform 1 0 4396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9360
timestamp 1677622389
transform 1 0 4348 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8175
timestamp 1677622389
transform 1 0 4348 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9272
timestamp 1677622389
transform 1 0 4444 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8024
timestamp 1677622389
transform 1 0 4460 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_8025
timestamp 1677622389
transform 1 0 4500 0 1 465
box -3 -3 3 3
use M2_M1  M2_M1_9273
timestamp 1677622389
transform 1 0 4508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9274
timestamp 1677622389
transform 1 0 4556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9275
timestamp 1677622389
transform 1 0 4564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9361
timestamp 1677622389
transform 1 0 4476 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8176
timestamp 1677622389
transform 1 0 4476 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9362
timestamp 1677622389
transform 1 0 4572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9276
timestamp 1677622389
transform 1 0 4620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9277
timestamp 1677622389
transform 1 0 4676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9363
timestamp 1677622389
transform 1 0 4596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8177
timestamp 1677622389
transform 1 0 4596 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9278
timestamp 1677622389
transform 1 0 4724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9279
timestamp 1677622389
transform 1 0 4780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9364
timestamp 1677622389
transform 1 0 4700 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8178
timestamp 1677622389
transform 1 0 4700 0 1 395
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_86
timestamp 1677622389
transform 1 0 48 0 1 370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_551
timestamp 1677622389
transform 1 0 72 0 1 370
box -8 -3 104 105
use FILL  FILL_10256
timestamp 1677622389
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_10257
timestamp 1677622389
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_10258
timestamp 1677622389
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_10259
timestamp 1677622389
transform 1 0 192 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_384
timestamp 1677622389
transform 1 0 200 0 1 370
box -8 -3 46 105
use FILL  FILL_10262
timestamp 1677622389
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_10263
timestamp 1677622389
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_10264
timestamp 1677622389
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_10265
timestamp 1677622389
transform 1 0 264 0 1 370
box -8 -3 16 105
use INVX2  INVX2_651
timestamp 1677622389
transform 1 0 272 0 1 370
box -9 -3 26 105
use FILL  FILL_10266
timestamp 1677622389
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_10267
timestamp 1677622389
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_10268
timestamp 1677622389
transform 1 0 304 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_385
timestamp 1677622389
transform -1 0 352 0 1 370
box -8 -3 46 105
use FILL  FILL_10269
timestamp 1677622389
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_10270
timestamp 1677622389
transform 1 0 360 0 1 370
box -8 -3 16 105
use FILL  FILL_10271
timestamp 1677622389
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_10272
timestamp 1677622389
transform 1 0 376 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_386
timestamp 1677622389
transform 1 0 384 0 1 370
box -8 -3 46 105
use FILL  FILL_10282
timestamp 1677622389
transform 1 0 424 0 1 370
box -8 -3 16 105
use INVX2  INVX2_653
timestamp 1677622389
transform 1 0 432 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_554
timestamp 1677622389
transform 1 0 448 0 1 370
box -8 -3 104 105
use FILL  FILL_10284
timestamp 1677622389
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_10285
timestamp 1677622389
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_10286
timestamp 1677622389
transform 1 0 560 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_417
timestamp 1677622389
transform 1 0 568 0 1 370
box -8 -3 46 105
use FILL  FILL_10287
timestamp 1677622389
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_10294
timestamp 1677622389
transform 1 0 616 0 1 370
box -8 -3 16 105
use FILL  FILL_10296
timestamp 1677622389
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_10297
timestamp 1677622389
transform 1 0 632 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_388
timestamp 1677622389
transform 1 0 640 0 1 370
box -8 -3 46 105
use FILL  FILL_10298
timestamp 1677622389
transform 1 0 680 0 1 370
box -8 -3 16 105
use INVX2  INVX2_655
timestamp 1677622389
transform 1 0 688 0 1 370
box -9 -3 26 105
use FILL  FILL_10305
timestamp 1677622389
transform 1 0 704 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_556
timestamp 1677622389
transform 1 0 712 0 1 370
box -8 -3 104 105
use FILL  FILL_10306
timestamp 1677622389
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_10307
timestamp 1677622389
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_10308
timestamp 1677622389
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_10309
timestamp 1677622389
transform 1 0 832 0 1 370
box -8 -3 16 105
use INVX2  INVX2_656
timestamp 1677622389
transform 1 0 840 0 1 370
box -9 -3 26 105
use FILL  FILL_10310
timestamp 1677622389
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_10311
timestamp 1677622389
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_10312
timestamp 1677622389
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_10313
timestamp 1677622389
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_10314
timestamp 1677622389
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_10315
timestamp 1677622389
transform 1 0 896 0 1 370
box -8 -3 16 105
use FILL  FILL_10316
timestamp 1677622389
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_10317
timestamp 1677622389
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_10318
timestamp 1677622389
transform 1 0 920 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_389
timestamp 1677622389
transform -1 0 968 0 1 370
box -8 -3 46 105
use INVX2  INVX2_657
timestamp 1677622389
transform 1 0 968 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_557
timestamp 1677622389
transform -1 0 1080 0 1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_107
timestamp 1677622389
transform 1 0 1080 0 1 370
box -8 -3 32 105
use FILL  FILL_10319
timestamp 1677622389
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_10320
timestamp 1677622389
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_10329
timestamp 1677622389
transform 1 0 1120 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_561
timestamp 1677622389
transform 1 0 1128 0 1 370
box -8 -3 104 105
use FILL  FILL_10330
timestamp 1677622389
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_10336
timestamp 1677622389
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_10338
timestamp 1677622389
transform 1 0 1240 0 1 370
box -8 -3 16 105
use FILL  FILL_10340
timestamp 1677622389
transform 1 0 1248 0 1 370
box -8 -3 16 105
use FILL  FILL_10341
timestamp 1677622389
transform 1 0 1256 0 1 370
box -8 -3 16 105
use FILL  FILL_10342
timestamp 1677622389
transform 1 0 1264 0 1 370
box -8 -3 16 105
use FILL  FILL_10343
timestamp 1677622389
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_10344
timestamp 1677622389
transform 1 0 1280 0 1 370
box -8 -3 16 105
use FILL  FILL_10345
timestamp 1677622389
transform 1 0 1288 0 1 370
box -8 -3 16 105
use FILL  FILL_10347
timestamp 1677622389
transform 1 0 1296 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_391
timestamp 1677622389
transform 1 0 1304 0 1 370
box -8 -3 46 105
use FILL  FILL_10349
timestamp 1677622389
transform 1 0 1344 0 1 370
box -8 -3 16 105
use FILL  FILL_10350
timestamp 1677622389
transform 1 0 1352 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_562
timestamp 1677622389
transform 1 0 1360 0 1 370
box -8 -3 104 105
use FILL  FILL_10351
timestamp 1677622389
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_10352
timestamp 1677622389
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_10353
timestamp 1677622389
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_10354
timestamp 1677622389
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_10355
timestamp 1677622389
transform 1 0 1488 0 1 370
box -8 -3 16 105
use INVX2  INVX2_659
timestamp 1677622389
transform -1 0 1512 0 1 370
box -9 -3 26 105
use FILL  FILL_10356
timestamp 1677622389
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_10357
timestamp 1677622389
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_10358
timestamp 1677622389
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_10359
timestamp 1677622389
transform 1 0 1536 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_563
timestamp 1677622389
transform -1 0 1640 0 1 370
box -8 -3 104 105
use FILL  FILL_10360
timestamp 1677622389
transform 1 0 1640 0 1 370
box -8 -3 16 105
use INVX2  INVX2_660
timestamp 1677622389
transform -1 0 1664 0 1 370
box -9 -3 26 105
use FILL  FILL_10361
timestamp 1677622389
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_10367
timestamp 1677622389
transform 1 0 1672 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_393
timestamp 1677622389
transform 1 0 1680 0 1 370
box -8 -3 46 105
use FILL  FILL_10368
timestamp 1677622389
transform 1 0 1720 0 1 370
box -8 -3 16 105
use FILL  FILL_10371
timestamp 1677622389
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_10373
timestamp 1677622389
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_10375
timestamp 1677622389
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_10376
timestamp 1677622389
transform 1 0 1752 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_566
timestamp 1677622389
transform -1 0 1856 0 1 370
box -8 -3 104 105
use FILL  FILL_10377
timestamp 1677622389
transform 1 0 1856 0 1 370
box -8 -3 16 105
use FILL  FILL_10378
timestamp 1677622389
transform 1 0 1864 0 1 370
box -8 -3 16 105
use FILL  FILL_10379
timestamp 1677622389
transform 1 0 1872 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_394
timestamp 1677622389
transform 1 0 1880 0 1 370
box -8 -3 46 105
use FILL  FILL_10380
timestamp 1677622389
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_10381
timestamp 1677622389
transform 1 0 1928 0 1 370
box -8 -3 16 105
use FILL  FILL_10382
timestamp 1677622389
transform 1 0 1936 0 1 370
box -8 -3 16 105
use INVX2  INVX2_662
timestamp 1677622389
transform 1 0 1944 0 1 370
box -9 -3 26 105
use FILL  FILL_10383
timestamp 1677622389
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_10384
timestamp 1677622389
transform 1 0 1968 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_395
timestamp 1677622389
transform 1 0 1976 0 1 370
box -8 -3 46 105
use FILL  FILL_10385
timestamp 1677622389
transform 1 0 2016 0 1 370
box -8 -3 16 105
use FILL  FILL_10386
timestamp 1677622389
transform 1 0 2024 0 1 370
box -8 -3 16 105
use FILL  FILL_10387
timestamp 1677622389
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_10388
timestamp 1677622389
transform 1 0 2040 0 1 370
box -8 -3 16 105
use INVX2  INVX2_663
timestamp 1677622389
transform 1 0 2048 0 1 370
box -9 -3 26 105
use FILL  FILL_10389
timestamp 1677622389
transform 1 0 2064 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_567
timestamp 1677622389
transform -1 0 2168 0 1 370
box -8 -3 104 105
use FILL  FILL_10390
timestamp 1677622389
transform 1 0 2168 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_568
timestamp 1677622389
transform -1 0 2272 0 1 370
box -8 -3 104 105
use FILL  FILL_10391
timestamp 1677622389
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_10392
timestamp 1677622389
transform 1 0 2280 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_569
timestamp 1677622389
transform -1 0 2384 0 1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_112
timestamp 1677622389
transform 1 0 2384 0 1 370
box -8 -3 32 105
use FILL  FILL_10393
timestamp 1677622389
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_10394
timestamp 1677622389
transform 1 0 2416 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_570
timestamp 1677622389
transform 1 0 2424 0 1 370
box -8 -3 104 105
use FILL  FILL_10395
timestamp 1677622389
transform 1 0 2520 0 1 370
box -8 -3 16 105
use INVX2  INVX2_664
timestamp 1677622389
transform 1 0 2528 0 1 370
box -9 -3 26 105
use FILL  FILL_10396
timestamp 1677622389
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_10397
timestamp 1677622389
transform 1 0 2552 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_182
timestamp 1677622389
transform -1 0 2592 0 1 370
box -8 -3 34 105
use FILL  FILL_10398
timestamp 1677622389
transform 1 0 2592 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_76
timestamp 1677622389
transform -1 0 2632 0 1 370
box -8 -3 40 105
use FILL  FILL_10399
timestamp 1677622389
transform 1 0 2632 0 1 370
box -8 -3 16 105
use FILL  FILL_10425
timestamp 1677622389
transform 1 0 2640 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_577
timestamp 1677622389
transform 1 0 2648 0 1 370
box -8 -3 104 105
use FILL  FILL_10426
timestamp 1677622389
transform 1 0 2744 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_578
timestamp 1677622389
transform 1 0 2752 0 1 370
box -8 -3 104 105
use FILL  FILL_10427
timestamp 1677622389
transform 1 0 2848 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_579
timestamp 1677622389
transform 1 0 2856 0 1 370
box -8 -3 104 105
use FILL  FILL_10428
timestamp 1677622389
transform 1 0 2952 0 1 370
box -8 -3 16 105
use FILL  FILL_10429
timestamp 1677622389
transform 1 0 2960 0 1 370
box -8 -3 16 105
use FILL  FILL_10430
timestamp 1677622389
transform 1 0 2968 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_113
timestamp 1677622389
transform -1 0 3000 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1677622389
transform 1 0 3000 0 1 370
box -8 -3 32 105
use FILL  FILL_10431
timestamp 1677622389
transform 1 0 3024 0 1 370
box -8 -3 16 105
use FILL  FILL_10432
timestamp 1677622389
transform 1 0 3032 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_77
timestamp 1677622389
transform -1 0 3072 0 1 370
box -8 -3 40 105
use FILL  FILL_10433
timestamp 1677622389
transform 1 0 3072 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_78
timestamp 1677622389
transform -1 0 3112 0 1 370
box -8 -3 40 105
use FILL  FILL_10434
timestamp 1677622389
transform 1 0 3112 0 1 370
box -8 -3 16 105
use FILL  FILL_10435
timestamp 1677622389
transform 1 0 3120 0 1 370
box -8 -3 16 105
use FILL  FILL_10436
timestamp 1677622389
transform 1 0 3128 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_115
timestamp 1677622389
transform 1 0 3136 0 1 370
box -8 -3 32 105
use FILL  FILL_10437
timestamp 1677622389
transform 1 0 3160 0 1 370
box -8 -3 16 105
use FILL  FILL_10438
timestamp 1677622389
transform 1 0 3168 0 1 370
box -8 -3 16 105
use FILL  FILL_10439
timestamp 1677622389
transform 1 0 3176 0 1 370
box -8 -3 16 105
use FILL  FILL_10440
timestamp 1677622389
transform 1 0 3184 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_580
timestamp 1677622389
transform 1 0 3192 0 1 370
box -8 -3 104 105
use FILL  FILL_10441
timestamp 1677622389
transform 1 0 3288 0 1 370
box -8 -3 16 105
use FILL  FILL_10442
timestamp 1677622389
transform 1 0 3296 0 1 370
box -8 -3 16 105
use FILL  FILL_10443
timestamp 1677622389
transform 1 0 3304 0 1 370
box -8 -3 16 105
use FILL  FILL_10444
timestamp 1677622389
transform 1 0 3312 0 1 370
box -8 -3 16 105
use FILL  FILL_10445
timestamp 1677622389
transform 1 0 3320 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_581
timestamp 1677622389
transform 1 0 3328 0 1 370
box -8 -3 104 105
use FILL  FILL_10446
timestamp 1677622389
transform 1 0 3424 0 1 370
box -8 -3 16 105
use FILL  FILL_10447
timestamp 1677622389
transform 1 0 3432 0 1 370
box -8 -3 16 105
use FILL  FILL_10448
timestamp 1677622389
transform 1 0 3440 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1677622389
transform 1 0 3448 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1677622389
transform 1 0 3472 0 1 370
box -8 -3 32 105
use FILL  FILL_10470
timestamp 1677622389
transform 1 0 3496 0 1 370
box -8 -3 16 105
use FILL  FILL_10471
timestamp 1677622389
transform 1 0 3504 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_53
timestamp 1677622389
transform 1 0 3512 0 1 370
box -8 -3 32 105
use FILL  FILL_10472
timestamp 1677622389
transform 1 0 3536 0 1 370
box -8 -3 16 105
use FILL  FILL_10476
timestamp 1677622389
transform 1 0 3544 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_55
timestamp 1677622389
transform -1 0 3576 0 1 370
box -8 -3 32 105
use M3_M2  M3_M2_8192
timestamp 1677622389
transform 1 0 3596 0 1 375
box -3 -3 3 3
use NAND2X1  NAND2X1_56
timestamp 1677622389
transform -1 0 3600 0 1 370
box -8 -3 32 105
use FILL  FILL_10477
timestamp 1677622389
transform 1 0 3600 0 1 370
box -8 -3 16 105
use FILL  FILL_10478
timestamp 1677622389
transform 1 0 3608 0 1 370
box -8 -3 16 105
use FILL  FILL_10479
timestamp 1677622389
transform 1 0 3616 0 1 370
box -8 -3 16 105
use FILL  FILL_10480
timestamp 1677622389
transform 1 0 3624 0 1 370
box -8 -3 16 105
use FILL  FILL_10481
timestamp 1677622389
transform 1 0 3632 0 1 370
box -8 -3 16 105
use FILL  FILL_10486
timestamp 1677622389
transform 1 0 3640 0 1 370
box -8 -3 16 105
use FILL  FILL_10488
timestamp 1677622389
transform 1 0 3648 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_423
timestamp 1677622389
transform 1 0 3656 0 1 370
box -8 -3 46 105
use FILL  FILL_10489
timestamp 1677622389
transform 1 0 3696 0 1 370
box -8 -3 16 105
use FILL  FILL_10490
timestamp 1677622389
transform 1 0 3704 0 1 370
box -8 -3 16 105
use FILL  FILL_10491
timestamp 1677622389
transform 1 0 3712 0 1 370
box -8 -3 16 105
use INVX2  INVX2_670
timestamp 1677622389
transform -1 0 3736 0 1 370
box -9 -3 26 105
use FILL  FILL_10492
timestamp 1677622389
transform 1 0 3736 0 1 370
box -8 -3 16 105
use FILL  FILL_10493
timestamp 1677622389
transform 1 0 3744 0 1 370
box -8 -3 16 105
use INVX2  INVX2_671
timestamp 1677622389
transform 1 0 3752 0 1 370
box -9 -3 26 105
use FILL  FILL_10495
timestamp 1677622389
transform 1 0 3768 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_424
timestamp 1677622389
transform -1 0 3816 0 1 370
box -8 -3 46 105
use FILL  FILL_10496
timestamp 1677622389
transform 1 0 3816 0 1 370
box -8 -3 16 105
use FILL  FILL_10497
timestamp 1677622389
transform 1 0 3824 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_588
timestamp 1677622389
transform 1 0 3832 0 1 370
box -8 -3 104 105
use FILL  FILL_10498
timestamp 1677622389
transform 1 0 3928 0 1 370
box -8 -3 16 105
use FILL  FILL_10508
timestamp 1677622389
transform 1 0 3936 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_590
timestamp 1677622389
transform 1 0 3944 0 1 370
box -8 -3 104 105
use FILL  FILL_10510
timestamp 1677622389
transform 1 0 4040 0 1 370
box -8 -3 16 105
use FILL  FILL_10511
timestamp 1677622389
transform 1 0 4048 0 1 370
box -8 -3 16 105
use FILL  FILL_10512
timestamp 1677622389
transform 1 0 4056 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_425
timestamp 1677622389
transform -1 0 4104 0 1 370
box -8 -3 46 105
use FILL  FILL_10513
timestamp 1677622389
transform 1 0 4104 0 1 370
box -8 -3 16 105
use FILL  FILL_10514
timestamp 1677622389
transform 1 0 4112 0 1 370
box -8 -3 16 105
use INVX2  INVX2_673
timestamp 1677622389
transform -1 0 4136 0 1 370
box -9 -3 26 105
use FILL  FILL_10515
timestamp 1677622389
transform 1 0 4136 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_426
timestamp 1677622389
transform 1 0 4144 0 1 370
box -8 -3 46 105
use FILL  FILL_10520
timestamp 1677622389
transform 1 0 4184 0 1 370
box -8 -3 16 105
use FILL  FILL_10522
timestamp 1677622389
transform 1 0 4192 0 1 370
box -8 -3 16 105
use INVX2  INVX2_676
timestamp 1677622389
transform -1 0 4216 0 1 370
box -9 -3 26 105
use FILL  FILL_10523
timestamp 1677622389
transform 1 0 4216 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8193
timestamp 1677622389
transform 1 0 4324 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_592
timestamp 1677622389
transform 1 0 4224 0 1 370
box -8 -3 104 105
use FILL  FILL_10524
timestamp 1677622389
transform 1 0 4320 0 1 370
box -8 -3 16 105
use FILL  FILL_10528
timestamp 1677622389
transform 1 0 4328 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8194
timestamp 1677622389
transform 1 0 4396 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_594
timestamp 1677622389
transform 1 0 4336 0 1 370
box -8 -3 104 105
use INVX2  INVX2_678
timestamp 1677622389
transform 1 0 4432 0 1 370
box -9 -3 26 105
use FILL  FILL_10530
timestamp 1677622389
transform 1 0 4448 0 1 370
box -8 -3 16 105
use FILL  FILL_10531
timestamp 1677622389
transform 1 0 4456 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8195
timestamp 1677622389
transform 1 0 4484 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_595
timestamp 1677622389
transform 1 0 4464 0 1 370
box -8 -3 104 105
use INVX2  INVX2_679
timestamp 1677622389
transform -1 0 4576 0 1 370
box -9 -3 26 105
use FILL  FILL_10532
timestamp 1677622389
transform 1 0 4576 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8196
timestamp 1677622389
transform 1 0 4596 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8197
timestamp 1677622389
transform 1 0 4636 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_596
timestamp 1677622389
transform 1 0 4584 0 1 370
box -8 -3 104 105
use FILL  FILL_10550
timestamp 1677622389
transform 1 0 4680 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_597
timestamp 1677622389
transform 1 0 4688 0 1 370
box -8 -3 104 105
use FILL  FILL_10551
timestamp 1677622389
transform 1 0 4784 0 1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_87
timestamp 1677622389
transform 1 0 4819 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_9379
timestamp 1677622389
transform 1 0 92 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9467
timestamp 1677622389
transform 1 0 140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9468
timestamp 1677622389
transform 1 0 172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9469
timestamp 1677622389
transform 1 0 180 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8291
timestamp 1677622389
transform 1 0 140 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8292
timestamp 1677622389
transform 1 0 180 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8330
timestamp 1677622389
transform 1 0 180 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8258
timestamp 1677622389
transform 1 0 204 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9380
timestamp 1677622389
transform 1 0 220 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8230
timestamp 1677622389
transform 1 0 332 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9381
timestamp 1677622389
transform 1 0 252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9470
timestamp 1677622389
transform 1 0 300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9471
timestamp 1677622389
transform 1 0 332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9472
timestamp 1677622389
transform 1 0 340 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8293
timestamp 1677622389
transform 1 0 300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8294
timestamp 1677622389
transform 1 0 340 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8259
timestamp 1677622389
transform 1 0 372 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9473
timestamp 1677622389
transform 1 0 372 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8231
timestamp 1677622389
transform 1 0 412 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9382
timestamp 1677622389
transform 1 0 388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9383
timestamp 1677622389
transform 1 0 396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9384
timestamp 1677622389
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9474
timestamp 1677622389
transform 1 0 388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9475
timestamp 1677622389
transform 1 0 404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9476
timestamp 1677622389
transform 1 0 420 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8295
timestamp 1677622389
transform 1 0 388 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8211
timestamp 1677622389
transform 1 0 556 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8232
timestamp 1677622389
transform 1 0 548 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9385
timestamp 1677622389
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9386
timestamp 1677622389
transform 1 0 540 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8260
timestamp 1677622389
transform 1 0 548 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9387
timestamp 1677622389
transform 1 0 556 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8261
timestamp 1677622389
transform 1 0 564 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9388
timestamp 1677622389
transform 1 0 572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9477
timestamp 1677622389
transform 1 0 476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9478
timestamp 1677622389
transform 1 0 532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9479
timestamp 1677622389
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9480
timestamp 1677622389
transform 1 0 564 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8296
timestamp 1677622389
transform 1 0 492 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8357
timestamp 1677622389
transform 1 0 492 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8297
timestamp 1677622389
transform 1 0 564 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8298
timestamp 1677622389
transform 1 0 580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8331
timestamp 1677622389
transform 1 0 572 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9481
timestamp 1677622389
transform 1 0 596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9482
timestamp 1677622389
transform 1 0 684 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8299
timestamp 1677622389
transform 1 0 684 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9389
timestamp 1677622389
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9483
timestamp 1677622389
transform 1 0 724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9484
timestamp 1677622389
transform 1 0 780 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8300
timestamp 1677622389
transform 1 0 724 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8301
timestamp 1677622389
transform 1 0 740 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8233
timestamp 1677622389
transform 1 0 892 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9390
timestamp 1677622389
transform 1 0 892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9485
timestamp 1677622389
transform 1 0 812 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8277
timestamp 1677622389
transform 1 0 852 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9391
timestamp 1677622389
transform 1 0 916 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9392
timestamp 1677622389
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9393
timestamp 1677622389
transform 1 0 940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9486
timestamp 1677622389
transform 1 0 860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9487
timestamp 1677622389
transform 1 0 908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9488
timestamp 1677622389
transform 1 0 924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9489
timestamp 1677622389
transform 1 0 940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9490
timestamp 1677622389
transform 1 0 948 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8302
timestamp 1677622389
transform 1 0 908 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8332
timestamp 1677622389
transform 1 0 932 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8303
timestamp 1677622389
transform 1 0 948 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8344
timestamp 1677622389
transform 1 0 948 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8234
timestamp 1677622389
transform 1 0 1060 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9394
timestamp 1677622389
transform 1 0 1060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9491
timestamp 1677622389
transform 1 0 972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9492
timestamp 1677622389
transform 1 0 980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9493
timestamp 1677622389
transform 1 0 1012 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8304
timestamp 1677622389
transform 1 0 972 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8305
timestamp 1677622389
transform 1 0 1012 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8333
timestamp 1677622389
transform 1 0 980 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8358
timestamp 1677622389
transform 1 0 972 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8212
timestamp 1677622389
transform 1 0 1076 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9371
timestamp 1677622389
transform 1 0 1076 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8262
timestamp 1677622389
transform 1 0 1076 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9395
timestamp 1677622389
transform 1 0 1092 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9372
timestamp 1677622389
transform 1 0 1116 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8263
timestamp 1677622389
transform 1 0 1108 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9373
timestamp 1677622389
transform 1 0 1140 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9396
timestamp 1677622389
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9494
timestamp 1677622389
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8334
timestamp 1677622389
transform 1 0 1124 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8264
timestamp 1677622389
transform 1 0 1148 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9495
timestamp 1677622389
transform 1 0 1148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9374
timestamp 1677622389
transform 1 0 1164 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9397
timestamp 1677622389
transform 1 0 1172 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8278
timestamp 1677622389
transform 1 0 1164 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9398
timestamp 1677622389
transform 1 0 1204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9496
timestamp 1677622389
transform 1 0 1204 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8306
timestamp 1677622389
transform 1 0 1204 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9497
timestamp 1677622389
transform 1 0 1220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9498
timestamp 1677622389
transform 1 0 1236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8213
timestamp 1677622389
transform 1 0 1252 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9399
timestamp 1677622389
transform 1 0 1252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9400
timestamp 1677622389
transform 1 0 1268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9499
timestamp 1677622389
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8307
timestamp 1677622389
transform 1 0 1260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8198
timestamp 1677622389
transform 1 0 1316 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8235
timestamp 1677622389
transform 1 0 1324 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8199
timestamp 1677622389
transform 1 0 1340 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8214
timestamp 1677622389
transform 1 0 1396 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8215
timestamp 1677622389
transform 1 0 1436 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8236
timestamp 1677622389
transform 1 0 1380 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9401
timestamp 1677622389
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9402
timestamp 1677622389
transform 1 0 1340 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8265
timestamp 1677622389
transform 1 0 1348 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9403
timestamp 1677622389
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9404
timestamp 1677622389
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9405
timestamp 1677622389
transform 1 0 1380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9500
timestamp 1677622389
transform 1 0 1348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9501
timestamp 1677622389
transform 1 0 1364 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8279
timestamp 1677622389
transform 1 0 1372 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8237
timestamp 1677622389
transform 1 0 1476 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9406
timestamp 1677622389
transform 1 0 1476 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8238
timestamp 1677622389
transform 1 0 1500 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9407
timestamp 1677622389
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8266
timestamp 1677622389
transform 1 0 1508 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9408
timestamp 1677622389
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9502
timestamp 1677622389
transform 1 0 1388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9503
timestamp 1677622389
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9504
timestamp 1677622389
transform 1 0 1452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9505
timestamp 1677622389
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9506
timestamp 1677622389
transform 1 0 1508 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8308
timestamp 1677622389
transform 1 0 1364 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8345
timestamp 1677622389
transform 1 0 1380 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8280
timestamp 1677622389
transform 1 0 1516 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8239
timestamp 1677622389
transform 1 0 1612 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9409
timestamp 1677622389
transform 1 0 1612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9410
timestamp 1677622389
transform 1 0 1628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9411
timestamp 1677622389
transform 1 0 1644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9507
timestamp 1677622389
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9508
timestamp 1677622389
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9509
timestamp 1677622389
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8346
timestamp 1677622389
transform 1 0 1500 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9510
timestamp 1677622389
transform 1 0 1636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9511
timestamp 1677622389
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8309
timestamp 1677622389
transform 1 0 1636 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8347
timestamp 1677622389
transform 1 0 1628 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9412
timestamp 1677622389
transform 1 0 1668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9413
timestamp 1677622389
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9414
timestamp 1677622389
transform 1 0 1692 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8281
timestamp 1677622389
transform 1 0 1676 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9512
timestamp 1677622389
transform 1 0 1684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9513
timestamp 1677622389
transform 1 0 1700 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8310
timestamp 1677622389
transform 1 0 1684 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8335
timestamp 1677622389
transform 1 0 1692 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8267
timestamp 1677622389
transform 1 0 1724 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9514
timestamp 1677622389
transform 1 0 1724 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8240
timestamp 1677622389
transform 1 0 1748 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8241
timestamp 1677622389
transform 1 0 1772 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9415
timestamp 1677622389
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9416
timestamp 1677622389
transform 1 0 1756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9417
timestamp 1677622389
transform 1 0 1772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9515
timestamp 1677622389
transform 1 0 1748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9516
timestamp 1677622389
transform 1 0 1764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9517
timestamp 1677622389
transform 1 0 1780 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8311
timestamp 1677622389
transform 1 0 1748 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9418
timestamp 1677622389
transform 1 0 1884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9518
timestamp 1677622389
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8216
timestamp 1677622389
transform 1 0 1948 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9419
timestamp 1677622389
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9519
timestamp 1677622389
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9520
timestamp 1677622389
transform 1 0 1956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9420
timestamp 1677622389
transform 1 0 2004 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8282
timestamp 1677622389
transform 1 0 2004 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8348
timestamp 1677622389
transform 1 0 2004 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9521
timestamp 1677622389
transform 1 0 2020 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8217
timestamp 1677622389
transform 1 0 2052 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8242
timestamp 1677622389
transform 1 0 2044 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9421
timestamp 1677622389
transform 1 0 2052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9522
timestamp 1677622389
transform 1 0 2044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9523
timestamp 1677622389
transform 1 0 2060 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8312
timestamp 1677622389
transform 1 0 2060 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8218
timestamp 1677622389
transform 1 0 2148 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8219
timestamp 1677622389
transform 1 0 2188 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9422
timestamp 1677622389
transform 1 0 2180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9524
timestamp 1677622389
transform 1 0 2100 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8283
timestamp 1677622389
transform 1 0 2108 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8284
timestamp 1677622389
transform 1 0 2132 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9525
timestamp 1677622389
transform 1 0 2156 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8285
timestamp 1677622389
transform 1 0 2180 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8313
timestamp 1677622389
transform 1 0 2156 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8349
timestamp 1677622389
transform 1 0 2164 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8243
timestamp 1677622389
transform 1 0 2196 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9423
timestamp 1677622389
transform 1 0 2196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9526
timestamp 1677622389
transform 1 0 2196 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8314
timestamp 1677622389
transform 1 0 2196 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8350
timestamp 1677622389
transform 1 0 2212 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8315
timestamp 1677622389
transform 1 0 2236 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8336
timestamp 1677622389
transform 1 0 2236 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9527
timestamp 1677622389
transform 1 0 2244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9424
timestamp 1677622389
transform 1 0 2340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9528
timestamp 1677622389
transform 1 0 2292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8316
timestamp 1677622389
transform 1 0 2260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8200
timestamp 1677622389
transform 1 0 2364 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8201
timestamp 1677622389
transform 1 0 2388 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8220
timestamp 1677622389
transform 1 0 2444 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9425
timestamp 1677622389
transform 1 0 2444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9529
timestamp 1677622389
transform 1 0 2364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9530
timestamp 1677622389
transform 1 0 2412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8317
timestamp 1677622389
transform 1 0 2364 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8318
timestamp 1677622389
transform 1 0 2404 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8337
timestamp 1677622389
transform 1 0 2412 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9531
timestamp 1677622389
transform 1 0 2468 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8244
timestamp 1677622389
transform 1 0 2556 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9426
timestamp 1677622389
transform 1 0 2556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9532
timestamp 1677622389
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9427
timestamp 1677622389
transform 1 0 2572 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8338
timestamp 1677622389
transform 1 0 2572 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9533
timestamp 1677622389
transform 1 0 2588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8359
timestamp 1677622389
transform 1 0 2580 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9576
timestamp 1677622389
transform 1 0 2620 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8221
timestamp 1677622389
transform 1 0 2652 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9428
timestamp 1677622389
transform 1 0 2652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9534
timestamp 1677622389
transform 1 0 2676 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8339
timestamp 1677622389
transform 1 0 2676 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9375
timestamp 1677622389
transform 1 0 2772 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8360
timestamp 1677622389
transform 1 0 2772 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8268
timestamp 1677622389
transform 1 0 2796 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9535
timestamp 1677622389
transform 1 0 2796 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8245
timestamp 1677622389
transform 1 0 2820 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9429
timestamp 1677622389
transform 1 0 2820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9536
timestamp 1677622389
transform 1 0 2860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9537
timestamp 1677622389
transform 1 0 2900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9577
timestamp 1677622389
transform 1 0 2804 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8319
timestamp 1677622389
transform 1 0 2820 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9538
timestamp 1677622389
transform 1 0 2916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8202
timestamp 1677622389
transform 1 0 3028 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9430
timestamp 1677622389
transform 1 0 3028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9539
timestamp 1677622389
transform 1 0 2988 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8320
timestamp 1677622389
transform 1 0 3028 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8246
timestamp 1677622389
transform 1 0 3052 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9431
timestamp 1677622389
transform 1 0 3044 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8361
timestamp 1677622389
transform 1 0 3044 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9540
timestamp 1677622389
transform 1 0 3060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9541
timestamp 1677622389
transform 1 0 3068 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8351
timestamp 1677622389
transform 1 0 3060 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9542
timestamp 1677622389
transform 1 0 3084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8247
timestamp 1677622389
transform 1 0 3100 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9432
timestamp 1677622389
transform 1 0 3100 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8222
timestamp 1677622389
transform 1 0 3124 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9376
timestamp 1677622389
transform 1 0 3124 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9433
timestamp 1677622389
transform 1 0 3116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9434
timestamp 1677622389
transform 1 0 3132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9543
timestamp 1677622389
transform 1 0 3156 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8203
timestamp 1677622389
transform 1 0 3172 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8204
timestamp 1677622389
transform 1 0 3204 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8223
timestamp 1677622389
transform 1 0 3196 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9435
timestamp 1677622389
transform 1 0 3172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9544
timestamp 1677622389
transform 1 0 3196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9545
timestamp 1677622389
transform 1 0 3268 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8321
timestamp 1677622389
transform 1 0 3268 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8205
timestamp 1677622389
transform 1 0 3284 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8206
timestamp 1677622389
transform 1 0 3300 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8207
timestamp 1677622389
transform 1 0 3340 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8248
timestamp 1677622389
transform 1 0 3308 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9436
timestamp 1677622389
transform 1 0 3284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9546
timestamp 1677622389
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8224
timestamp 1677622389
transform 1 0 3420 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8269
timestamp 1677622389
transform 1 0 3412 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9437
timestamp 1677622389
transform 1 0 3420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9547
timestamp 1677622389
transform 1 0 3412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8286
timestamp 1677622389
transform 1 0 3420 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9578
timestamp 1677622389
transform 1 0 3420 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8340
timestamp 1677622389
transform 1 0 3420 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9438
timestamp 1677622389
transform 1 0 3444 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8322
timestamp 1677622389
transform 1 0 3444 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9579
timestamp 1677622389
transform 1 0 3468 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8341
timestamp 1677622389
transform 1 0 3468 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9548
timestamp 1677622389
transform 1 0 3484 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8323
timestamp 1677622389
transform 1 0 3484 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8225
timestamp 1677622389
transform 1 0 3508 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9377
timestamp 1677622389
transform 1 0 3508 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8270
timestamp 1677622389
transform 1 0 3500 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9439
timestamp 1677622389
transform 1 0 3508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9549
timestamp 1677622389
transform 1 0 3500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9440
timestamp 1677622389
transform 1 0 3532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9550
timestamp 1677622389
transform 1 0 3524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9441
timestamp 1677622389
transform 1 0 3556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9551
timestamp 1677622389
transform 1 0 3564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9378
timestamp 1677622389
transform 1 0 3596 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9442
timestamp 1677622389
transform 1 0 3596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9552
timestamp 1677622389
transform 1 0 3588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9580
timestamp 1677622389
transform 1 0 3588 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8352
timestamp 1677622389
transform 1 0 3588 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8271
timestamp 1677622389
transform 1 0 3612 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9581
timestamp 1677622389
transform 1 0 3628 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9443
timestamp 1677622389
transform 1 0 3636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9582
timestamp 1677622389
transform 1 0 3644 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8353
timestamp 1677622389
transform 1 0 3644 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8249
timestamp 1677622389
transform 1 0 3660 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9444
timestamp 1677622389
transform 1 0 3660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9553
timestamp 1677622389
transform 1 0 3684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9554
timestamp 1677622389
transform 1 0 3740 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8324
timestamp 1677622389
transform 1 0 3684 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8325
timestamp 1677622389
transform 1 0 3708 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8250
timestamp 1677622389
transform 1 0 3764 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8251
timestamp 1677622389
transform 1 0 3844 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9445
timestamp 1677622389
transform 1 0 3764 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8272
timestamp 1677622389
transform 1 0 3828 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9555
timestamp 1677622389
transform 1 0 3796 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8342
timestamp 1677622389
transform 1 0 3788 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8273
timestamp 1677622389
transform 1 0 3876 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9556
timestamp 1677622389
transform 1 0 3876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9446
timestamp 1677622389
transform 1 0 3932 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8287
timestamp 1677622389
transform 1 0 3932 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8252
timestamp 1677622389
transform 1 0 3972 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9557
timestamp 1677622389
transform 1 0 3980 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8226
timestamp 1677622389
transform 1 0 4028 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8208
timestamp 1677622389
transform 1 0 4060 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8227
timestamp 1677622389
transform 1 0 4148 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8228
timestamp 1677622389
transform 1 0 4164 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8253
timestamp 1677622389
transform 1 0 4076 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8254
timestamp 1677622389
transform 1 0 4108 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9447
timestamp 1677622389
transform 1 0 4012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9448
timestamp 1677622389
transform 1 0 4028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9449
timestamp 1677622389
transform 1 0 4044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9450
timestamp 1677622389
transform 1 0 4060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9451
timestamp 1677622389
transform 1 0 4148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9452
timestamp 1677622389
transform 1 0 4164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9558
timestamp 1677622389
transform 1 0 4004 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8288
timestamp 1677622389
transform 1 0 4028 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9559
timestamp 1677622389
transform 1 0 4036 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8289
timestamp 1677622389
transform 1 0 4044 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9560
timestamp 1677622389
transform 1 0 4084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8290
timestamp 1677622389
transform 1 0 4100 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8274
timestamp 1677622389
transform 1 0 4172 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9453
timestamp 1677622389
transform 1 0 4180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9561
timestamp 1677622389
transform 1 0 4140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9562
timestamp 1677622389
transform 1 0 4148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9563
timestamp 1677622389
transform 1 0 4172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8354
timestamp 1677622389
transform 1 0 4004 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8362
timestamp 1677622389
transform 1 0 4172 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8209
timestamp 1677622389
transform 1 0 4204 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8210
timestamp 1677622389
transform 1 0 4292 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8229
timestamp 1677622389
transform 1 0 4244 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9454
timestamp 1677622389
transform 1 0 4292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9455
timestamp 1677622389
transform 1 0 4308 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9564
timestamp 1677622389
transform 1 0 4212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9565
timestamp 1677622389
transform 1 0 4244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9456
timestamp 1677622389
transform 1 0 4324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9566
timestamp 1677622389
transform 1 0 4316 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8363
timestamp 1677622389
transform 1 0 4316 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9457
timestamp 1677622389
transform 1 0 4364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9567
timestamp 1677622389
transform 1 0 4372 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8343
timestamp 1677622389
transform 1 0 4372 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9458
timestamp 1677622389
transform 1 0 4396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9568
timestamp 1677622389
transform 1 0 4436 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8255
timestamp 1677622389
transform 1 0 4460 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9459
timestamp 1677622389
transform 1 0 4468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9460
timestamp 1677622389
transform 1 0 4484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9569
timestamp 1677622389
transform 1 0 4460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9570
timestamp 1677622389
transform 1 0 4500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9461
timestamp 1677622389
transform 1 0 4548 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8326
timestamp 1677622389
transform 1 0 4540 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9462
timestamp 1677622389
transform 1 0 4556 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8327
timestamp 1677622389
transform 1 0 4564 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8256
timestamp 1677622389
transform 1 0 4620 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8275
timestamp 1677622389
transform 1 0 4612 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9463
timestamp 1677622389
transform 1 0 4620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9464
timestamp 1677622389
transform 1 0 4636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9571
timestamp 1677622389
transform 1 0 4612 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8355
timestamp 1677622389
transform 1 0 4620 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9572
timestamp 1677622389
transform 1 0 4644 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8328
timestamp 1677622389
transform 1 0 4644 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8356
timestamp 1677622389
transform 1 0 4668 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8257
timestamp 1677622389
transform 1 0 4708 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9465
timestamp 1677622389
transform 1 0 4684 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8276
timestamp 1677622389
transform 1 0 4748 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9466
timestamp 1677622389
transform 1 0 4780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9573
timestamp 1677622389
transform 1 0 4708 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9574
timestamp 1677622389
transform 1 0 4764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9575
timestamp 1677622389
transform 1 0 4772 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8329
timestamp 1677622389
transform 1 0 4772 0 1 315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_88
timestamp 1677622389
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_10260
timestamp 1677622389
transform 1 0 72 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_552
timestamp 1677622389
transform 1 0 80 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_650
timestamp 1677622389
transform -1 0 192 0 -1 370
box -9 -3 26 105
use FILL  FILL_10261
timestamp 1677622389
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_10273
timestamp 1677622389
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_10274
timestamp 1677622389
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_10275
timestamp 1677622389
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_10276
timestamp 1677622389
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_10277
timestamp 1677622389
transform 1 0 232 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_553
timestamp 1677622389
transform 1 0 240 0 -1 370
box -8 -3 104 105
use FILL  FILL_10278
timestamp 1677622389
transform 1 0 336 0 -1 370
box -8 -3 16 105
use FILL  FILL_10279
timestamp 1677622389
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_10280
timestamp 1677622389
transform 1 0 352 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_652
timestamp 1677622389
transform -1 0 376 0 -1 370
box -9 -3 26 105
use FILL  FILL_10281
timestamp 1677622389
transform 1 0 376 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_387
timestamp 1677622389
transform 1 0 384 0 -1 370
box -8 -3 46 105
use FILL  FILL_10283
timestamp 1677622389
transform 1 0 424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10288
timestamp 1677622389
transform 1 0 432 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_555
timestamp 1677622389
transform 1 0 440 0 -1 370
box -8 -3 104 105
use OAI22X1  OAI22X1_418
timestamp 1677622389
transform 1 0 536 0 -1 370
box -8 -3 46 105
use FILL  FILL_10289
timestamp 1677622389
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_10290
timestamp 1677622389
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10291
timestamp 1677622389
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_10292
timestamp 1677622389
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_10293
timestamp 1677622389
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_10295
timestamp 1677622389
transform 1 0 616 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_654
timestamp 1677622389
transform 1 0 624 0 -1 370
box -9 -3 26 105
use FILL  FILL_10299
timestamp 1677622389
transform 1 0 640 0 -1 370
box -8 -3 16 105
use FILL  FILL_10300
timestamp 1677622389
transform 1 0 648 0 -1 370
box -8 -3 16 105
use FILL  FILL_10301
timestamp 1677622389
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_10302
timestamp 1677622389
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_10303
timestamp 1677622389
transform 1 0 672 0 -1 370
box -8 -3 16 105
use FILL  FILL_10304
timestamp 1677622389
transform 1 0 680 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8364
timestamp 1677622389
transform 1 0 732 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_558
timestamp 1677622389
transform 1 0 688 0 -1 370
box -8 -3 104 105
use FILL  FILL_10321
timestamp 1677622389
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_10322
timestamp 1677622389
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_10323
timestamp 1677622389
transform 1 0 800 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_559
timestamp 1677622389
transform -1 0 904 0 -1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_390
timestamp 1677622389
transform 1 0 904 0 -1 370
box -8 -3 46 105
use FILL  FILL_10324
timestamp 1677622389
transform 1 0 944 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_658
timestamp 1677622389
transform 1 0 952 0 -1 370
box -9 -3 26 105
use FILL  FILL_10325
timestamp 1677622389
transform 1 0 968 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_560
timestamp 1677622389
transform -1 0 1072 0 -1 370
box -8 -3 104 105
use FILL  FILL_10326
timestamp 1677622389
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10327
timestamp 1677622389
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_108
timestamp 1677622389
transform 1 0 1088 0 -1 370
box -8 -3 32 105
use FILL  FILL_10328
timestamp 1677622389
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8365
timestamp 1677622389
transform 1 0 1140 0 1 275
box -3 -3 3 3
use NOR2X1  NOR2X1_109
timestamp 1677622389
transform 1 0 1120 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1677622389
transform 1 0 1144 0 -1 370
box -8 -3 32 105
use FILL  FILL_10331
timestamp 1677622389
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_10332
timestamp 1677622389
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use FILL  FILL_10333
timestamp 1677622389
transform 1 0 1184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10334
timestamp 1677622389
transform 1 0 1192 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_111
timestamp 1677622389
transform 1 0 1200 0 -1 370
box -8 -3 32 105
use FILL  FILL_10335
timestamp 1677622389
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_10337
timestamp 1677622389
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8366
timestamp 1677622389
transform 1 0 1252 0 1 275
box -3 -3 3 3
use FILL  FILL_10339
timestamp 1677622389
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_419
timestamp 1677622389
transform 1 0 1248 0 -1 370
box -8 -3 46 105
use FILL  FILL_10346
timestamp 1677622389
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_10348
timestamp 1677622389
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_10362
timestamp 1677622389
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_10363
timestamp 1677622389
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_10364
timestamp 1677622389
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use FILL  FILL_10365
timestamp 1677622389
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8367
timestamp 1677622389
transform 1 0 1348 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_420
timestamp 1677622389
transform -1 0 1376 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_661
timestamp 1677622389
transform 1 0 1376 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_564
timestamp 1677622389
transform -1 0 1488 0 -1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_392
timestamp 1677622389
transform 1 0 1488 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_565
timestamp 1677622389
transform -1 0 1624 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_8368
timestamp 1677622389
transform 1 0 1652 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_421
timestamp 1677622389
transform 1 0 1624 0 -1 370
box -8 -3 46 105
use FILL  FILL_10366
timestamp 1677622389
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8369
timestamp 1677622389
transform 1 0 1700 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_422
timestamp 1677622389
transform 1 0 1672 0 -1 370
box -8 -3 46 105
use FILL  FILL_10369
timestamp 1677622389
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_10370
timestamp 1677622389
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_10372
timestamp 1677622389
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_10374
timestamp 1677622389
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_396
timestamp 1677622389
transform 1 0 1744 0 -1 370
box -8 -3 46 105
use FILL  FILL_10400
timestamp 1677622389
transform 1 0 1784 0 -1 370
box -8 -3 16 105
use FILL  FILL_10401
timestamp 1677622389
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_571
timestamp 1677622389
transform -1 0 1896 0 -1 370
box -8 -3 104 105
use FILL  FILL_10402
timestamp 1677622389
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_572
timestamp 1677622389
transform -1 0 2000 0 -1 370
box -8 -3 104 105
use FILL  FILL_10403
timestamp 1677622389
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use FILL  FILL_10404
timestamp 1677622389
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_10405
timestamp 1677622389
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_397
timestamp 1677622389
transform -1 0 2064 0 -1 370
box -8 -3 46 105
use FILL  FILL_10406
timestamp 1677622389
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_10407
timestamp 1677622389
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10408
timestamp 1677622389
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_10409
timestamp 1677622389
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_573
timestamp 1677622389
transform -1 0 2192 0 -1 370
box -8 -3 104 105
use FILL  FILL_10410
timestamp 1677622389
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_10411
timestamp 1677622389
transform 1 0 2200 0 -1 370
box -8 -3 16 105
use FILL  FILL_10412
timestamp 1677622389
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_665
timestamp 1677622389
transform 1 0 2216 0 -1 370
box -9 -3 26 105
use FILL  FILL_10413
timestamp 1677622389
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_10414
timestamp 1677622389
transform 1 0 2240 0 -1 370
box -8 -3 16 105
use FILL  FILL_10415
timestamp 1677622389
transform 1 0 2248 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_574
timestamp 1677622389
transform -1 0 2352 0 -1 370
box -8 -3 104 105
use FILL  FILL_10416
timestamp 1677622389
transform 1 0 2352 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_575
timestamp 1677622389
transform -1 0 2456 0 -1 370
box -8 -3 104 105
use FILL  FILL_10417
timestamp 1677622389
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_10418
timestamp 1677622389
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_576
timestamp 1677622389
transform -1 0 2568 0 -1 370
box -8 -3 104 105
use FILL  FILL_10419
timestamp 1677622389
transform 1 0 2568 0 -1 370
box -8 -3 16 105
use FILL  FILL_10420
timestamp 1677622389
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_10421
timestamp 1677622389
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10422
timestamp 1677622389
transform 1 0 2592 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1677622389
transform 1 0 2600 0 -1 370
box -8 -3 32 105
use FILL  FILL_10423
timestamp 1677622389
transform 1 0 2624 0 -1 370
box -8 -3 16 105
use FILL  FILL_10424
timestamp 1677622389
transform 1 0 2632 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_582
timestamp 1677622389
transform 1 0 2640 0 -1 370
box -8 -3 104 105
use FILL  FILL_10449
timestamp 1677622389
transform 1 0 2736 0 -1 370
box -8 -3 16 105
use FILL  FILL_10450
timestamp 1677622389
transform 1 0 2744 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_116
timestamp 1677622389
transform -1 0 2776 0 -1 370
box -8 -3 32 105
use FILL  FILL_10451
timestamp 1677622389
transform 1 0 2776 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1677622389
transform 1 0 2784 0 -1 370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_583
timestamp 1677622389
transform 1 0 2808 0 -1 370
box -8 -3 104 105
use FILL  FILL_10452
timestamp 1677622389
transform 1 0 2904 0 -1 370
box -8 -3 16 105
use FILL  FILL_10453
timestamp 1677622389
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_10454
timestamp 1677622389
transform 1 0 2920 0 -1 370
box -8 -3 16 105
use FILL  FILL_10455
timestamp 1677622389
transform 1 0 2928 0 -1 370
box -8 -3 16 105
use FILL  FILL_10456
timestamp 1677622389
transform 1 0 2936 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_584
timestamp 1677622389
transform -1 0 3040 0 -1 370
box -8 -3 104 105
use FILL  FILL_10457
timestamp 1677622389
transform 1 0 3040 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_666
timestamp 1677622389
transform 1 0 3048 0 -1 370
box -9 -3 26 105
use FILL  FILL_10458
timestamp 1677622389
transform 1 0 3064 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_667
timestamp 1677622389
transform -1 0 3088 0 -1 370
box -9 -3 26 105
use FILL  FILL_10459
timestamp 1677622389
transform 1 0 3088 0 -1 370
box -8 -3 16 105
use FILL  FILL_10460
timestamp 1677622389
transform 1 0 3096 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_668
timestamp 1677622389
transform -1 0 3120 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_117
timestamp 1677622389
transform 1 0 3120 0 -1 370
box -8 -3 32 105
use FILL  FILL_10461
timestamp 1677622389
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use FILL  FILL_10462
timestamp 1677622389
transform 1 0 3152 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_585
timestamp 1677622389
transform 1 0 3160 0 -1 370
box -8 -3 104 105
use FILL  FILL_10463
timestamp 1677622389
transform 1 0 3256 0 -1 370
box -8 -3 16 105
use FILL  FILL_10464
timestamp 1677622389
transform 1 0 3264 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_586
timestamp 1677622389
transform 1 0 3272 0 -1 370
box -8 -3 104 105
use FILL  FILL_10465
timestamp 1677622389
transform 1 0 3368 0 -1 370
box -8 -3 16 105
use FILL  FILL_10466
timestamp 1677622389
transform 1 0 3376 0 -1 370
box -8 -3 16 105
use FILL  FILL_10467
timestamp 1677622389
transform 1 0 3384 0 -1 370
box -8 -3 16 105
use FILL  FILL_10468
timestamp 1677622389
transform 1 0 3392 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_49
timestamp 1677622389
transform 1 0 3400 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_669
timestamp 1677622389
transform 1 0 3424 0 -1 370
box -9 -3 26 105
use FILL  FILL_10469
timestamp 1677622389
transform 1 0 3440 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_51
timestamp 1677622389
transform 1 0 3448 0 -1 370
box -8 -3 32 105
use FILL  FILL_10473
timestamp 1677622389
transform 1 0 3472 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_54
timestamp 1677622389
transform -1 0 3504 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1677622389
transform 1 0 3504 0 -1 370
box -8 -3 32 105
use FILL  FILL_10474
timestamp 1677622389
transform 1 0 3528 0 -1 370
box -8 -3 16 105
use FILL  FILL_10475
timestamp 1677622389
transform 1 0 3536 0 -1 370
box -8 -3 16 105
use FILL  FILL_10482
timestamp 1677622389
transform 1 0 3544 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_183
timestamp 1677622389
transform 1 0 3552 0 -1 370
box -8 -3 34 105
use FILL  FILL_10483
timestamp 1677622389
transform 1 0 3584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10484
timestamp 1677622389
transform 1 0 3592 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_184
timestamp 1677622389
transform 1 0 3600 0 -1 370
box -8 -3 34 105
use FILL  FILL_10485
timestamp 1677622389
transform 1 0 3632 0 -1 370
box -8 -3 16 105
use FILL  FILL_10487
timestamp 1677622389
transform 1 0 3640 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_587
timestamp 1677622389
transform 1 0 3648 0 -1 370
box -8 -3 104 105
use FILL  FILL_10494
timestamp 1677622389
transform 1 0 3744 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_589
timestamp 1677622389
transform 1 0 3752 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_8370
timestamp 1677622389
transform 1 0 3860 0 1 275
box -3 -3 3 3
use FILL  FILL_10499
timestamp 1677622389
transform 1 0 3848 0 -1 370
box -8 -3 16 105
use FILL  FILL_10500
timestamp 1677622389
transform 1 0 3856 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_672
timestamp 1677622389
transform 1 0 3864 0 -1 370
box -9 -3 26 105
use FILL  FILL_10501
timestamp 1677622389
transform 1 0 3880 0 -1 370
box -8 -3 16 105
use FILL  FILL_10502
timestamp 1677622389
transform 1 0 3888 0 -1 370
box -8 -3 16 105
use FILL  FILL_10503
timestamp 1677622389
transform 1 0 3896 0 -1 370
box -8 -3 16 105
use FILL  FILL_10504
timestamp 1677622389
transform 1 0 3904 0 -1 370
box -8 -3 16 105
use FILL  FILL_10505
timestamp 1677622389
transform 1 0 3912 0 -1 370
box -8 -3 16 105
use FILL  FILL_10506
timestamp 1677622389
transform 1 0 3920 0 -1 370
box -8 -3 16 105
use FILL  FILL_10507
timestamp 1677622389
transform 1 0 3928 0 -1 370
box -8 -3 16 105
use FILL  FILL_10509
timestamp 1677622389
transform 1 0 3936 0 -1 370
box -8 -3 16 105
use FILL  FILL_10516
timestamp 1677622389
transform 1 0 3944 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_674
timestamp 1677622389
transform 1 0 3952 0 -1 370
box -9 -3 26 105
use FILL  FILL_10517
timestamp 1677622389
transform 1 0 3968 0 -1 370
box -8 -3 16 105
use FILL  FILL_10518
timestamp 1677622389
transform 1 0 3976 0 -1 370
box -8 -3 16 105
use FILL  FILL_10519
timestamp 1677622389
transform 1 0 3984 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_427
timestamp 1677622389
transform -1 0 4032 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_675
timestamp 1677622389
transform -1 0 4048 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_591
timestamp 1677622389
transform 1 0 4048 0 -1 370
box -8 -3 104 105
use OAI22X1  OAI22X1_428
timestamp 1677622389
transform 1 0 4144 0 -1 370
box -8 -3 46 105
use FILL  FILL_10521
timestamp 1677622389
transform 1 0 4184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10525
timestamp 1677622389
transform 1 0 4192 0 -1 370
box -8 -3 16 105
use FILL  FILL_10526
timestamp 1677622389
transform 1 0 4200 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_593
timestamp 1677622389
transform -1 0 4304 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_677
timestamp 1677622389
transform 1 0 4304 0 -1 370
box -9 -3 26 105
use FILL  FILL_10527
timestamp 1677622389
transform 1 0 4320 0 -1 370
box -8 -3 16 105
use FILL  FILL_10529
timestamp 1677622389
transform 1 0 4328 0 -1 370
box -8 -3 16 105
use FILL  FILL_10533
timestamp 1677622389
transform 1 0 4336 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_429
timestamp 1677622389
transform 1 0 4344 0 -1 370
box -8 -3 46 105
use FILL  FILL_10534
timestamp 1677622389
transform 1 0 4384 0 -1 370
box -8 -3 16 105
use FILL  FILL_10535
timestamp 1677622389
transform 1 0 4392 0 -1 370
box -8 -3 16 105
use FILL  FILL_10536
timestamp 1677622389
transform 1 0 4400 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_680
timestamp 1677622389
transform 1 0 4408 0 -1 370
box -9 -3 26 105
use FILL  FILL_10537
timestamp 1677622389
transform 1 0 4424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10538
timestamp 1677622389
transform 1 0 4432 0 -1 370
box -8 -3 16 105
use FILL  FILL_10539
timestamp 1677622389
transform 1 0 4440 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_430
timestamp 1677622389
transform -1 0 4488 0 -1 370
box -8 -3 46 105
use FILL  FILL_10540
timestamp 1677622389
transform 1 0 4488 0 -1 370
box -8 -3 16 105
use FILL  FILL_10541
timestamp 1677622389
transform 1 0 4496 0 -1 370
box -8 -3 16 105
use FILL  FILL_10542
timestamp 1677622389
transform 1 0 4504 0 -1 370
box -8 -3 16 105
use FILL  FILL_10543
timestamp 1677622389
transform 1 0 4512 0 -1 370
box -8 -3 16 105
use FILL  FILL_10544
timestamp 1677622389
transform 1 0 4520 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_681
timestamp 1677622389
transform -1 0 4544 0 -1 370
box -9 -3 26 105
use FILL  FILL_10545
timestamp 1677622389
transform 1 0 4544 0 -1 370
box -8 -3 16 105
use FILL  FILL_10546
timestamp 1677622389
transform 1 0 4552 0 -1 370
box -8 -3 16 105
use FILL  FILL_10547
timestamp 1677622389
transform 1 0 4560 0 -1 370
box -8 -3 16 105
use FILL  FILL_10548
timestamp 1677622389
transform 1 0 4568 0 -1 370
box -8 -3 16 105
use FILL  FILL_10549
timestamp 1677622389
transform 1 0 4576 0 -1 370
box -8 -3 16 105
use FILL  FILL_10552
timestamp 1677622389
transform 1 0 4584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10553
timestamp 1677622389
transform 1 0 4592 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8371
timestamp 1677622389
transform 1 0 4612 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_431
timestamp 1677622389
transform -1 0 4640 0 -1 370
box -8 -3 46 105
use FILL  FILL_10554
timestamp 1677622389
transform 1 0 4640 0 -1 370
box -8 -3 16 105
use FILL  FILL_10555
timestamp 1677622389
transform 1 0 4648 0 -1 370
box -8 -3 16 105
use FILL  FILL_10556
timestamp 1677622389
transform 1 0 4656 0 -1 370
box -8 -3 16 105
use FILL  FILL_10557
timestamp 1677622389
transform 1 0 4664 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_598
timestamp 1677622389
transform 1 0 4672 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_682
timestamp 1677622389
transform -1 0 4784 0 -1 370
box -9 -3 26 105
use FILL  FILL_10558
timestamp 1677622389
transform 1 0 4784 0 -1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_89
timestamp 1677622389
transform 1 0 4843 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_8403
timestamp 1677622389
transform 1 0 124 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9588
timestamp 1677622389
transform 1 0 116 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8431
timestamp 1677622389
transform 1 0 172 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8487
timestamp 1677622389
transform 1 0 164 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8404
timestamp 1677622389
transform 1 0 204 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9589
timestamp 1677622389
transform 1 0 172 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8488
timestamp 1677622389
transform 1 0 180 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9590
timestamp 1677622389
transform 1 0 188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9591
timestamp 1677622389
transform 1 0 204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9746
timestamp 1677622389
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9747
timestamp 1677622389
transform 1 0 180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8489
timestamp 1677622389
transform 1 0 212 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8384
timestamp 1677622389
transform 1 0 228 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8432
timestamp 1677622389
transform 1 0 236 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8433
timestamp 1677622389
transform 1 0 268 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9592
timestamp 1677622389
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9593
timestamp 1677622389
transform 1 0 228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9748
timestamp 1677622389
transform 1 0 212 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8490
timestamp 1677622389
transform 1 0 244 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9594
timestamp 1677622389
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9595
timestamp 1677622389
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9749
timestamp 1677622389
transform 1 0 236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9750
timestamp 1677622389
transform 1 0 244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9751
timestamp 1677622389
transform 1 0 260 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8598
timestamp 1677622389
transform 1 0 260 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8385
timestamp 1677622389
transform 1 0 316 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8434
timestamp 1677622389
transform 1 0 300 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8435
timestamp 1677622389
transform 1 0 332 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9596
timestamp 1677622389
transform 1 0 308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9597
timestamp 1677622389
transform 1 0 316 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8491
timestamp 1677622389
transform 1 0 324 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9598
timestamp 1677622389
transform 1 0 332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9752
timestamp 1677622389
transform 1 0 300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9753
timestamp 1677622389
transform 1 0 324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8436
timestamp 1677622389
transform 1 0 356 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9599
timestamp 1677622389
transform 1 0 356 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8372
timestamp 1677622389
transform 1 0 372 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8405
timestamp 1677622389
transform 1 0 372 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8437
timestamp 1677622389
transform 1 0 404 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9600
timestamp 1677622389
transform 1 0 372 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8492
timestamp 1677622389
transform 1 0 380 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9601
timestamp 1677622389
transform 1 0 388 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8493
timestamp 1677622389
transform 1 0 396 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9602
timestamp 1677622389
transform 1 0 404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9754
timestamp 1677622389
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9755
timestamp 1677622389
transform 1 0 380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9756
timestamp 1677622389
transform 1 0 396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9757
timestamp 1677622389
transform 1 0 404 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8548
timestamp 1677622389
transform 1 0 380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8438
timestamp 1677622389
transform 1 0 420 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9603
timestamp 1677622389
transform 1 0 436 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8439
timestamp 1677622389
transform 1 0 460 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9758
timestamp 1677622389
transform 1 0 460 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8494
timestamp 1677622389
transform 1 0 476 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8406
timestamp 1677622389
transform 1 0 524 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8440
timestamp 1677622389
transform 1 0 508 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8373
timestamp 1677622389
transform 1 0 572 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8377
timestamp 1677622389
transform 1 0 564 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8441
timestamp 1677622389
transform 1 0 548 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9604
timestamp 1677622389
transform 1 0 484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9605
timestamp 1677622389
transform 1 0 492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9606
timestamp 1677622389
transform 1 0 508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9607
timestamp 1677622389
transform 1 0 524 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8528
timestamp 1677622389
transform 1 0 484 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8495
timestamp 1677622389
transform 1 0 532 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9608
timestamp 1677622389
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9609
timestamp 1677622389
transform 1 0 556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9759
timestamp 1677622389
transform 1 0 500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9760
timestamp 1677622389
transform 1 0 516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9761
timestamp 1677622389
transform 1 0 524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9762
timestamp 1677622389
transform 1 0 548 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8529
timestamp 1677622389
transform 1 0 556 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9610
timestamp 1677622389
transform 1 0 572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9763
timestamp 1677622389
transform 1 0 564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9764
timestamp 1677622389
transform 1 0 572 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8549
timestamp 1677622389
transform 1 0 524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8550
timestamp 1677622389
transform 1 0 548 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8599
timestamp 1677622389
transform 1 0 564 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8386
timestamp 1677622389
transform 1 0 620 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8407
timestamp 1677622389
transform 1 0 612 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9611
timestamp 1677622389
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9612
timestamp 1677622389
transform 1 0 612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9613
timestamp 1677622389
transform 1 0 620 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8408
timestamp 1677622389
transform 1 0 676 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9614
timestamp 1677622389
transform 1 0 660 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8496
timestamp 1677622389
transform 1 0 668 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9615
timestamp 1677622389
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9616
timestamp 1677622389
transform 1 0 684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9765
timestamp 1677622389
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9766
timestamp 1677622389
transform 1 0 652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9767
timestamp 1677622389
transform 1 0 668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9768
timestamp 1677622389
transform 1 0 676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8551
timestamp 1677622389
transform 1 0 644 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8442
timestamp 1677622389
transform 1 0 700 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9617
timestamp 1677622389
transform 1 0 700 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8497
timestamp 1677622389
transform 1 0 708 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8374
timestamp 1677622389
transform 1 0 740 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8378
timestamp 1677622389
transform 1 0 740 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8409
timestamp 1677622389
transform 1 0 748 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9618
timestamp 1677622389
transform 1 0 740 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8443
timestamp 1677622389
transform 1 0 756 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9619
timestamp 1677622389
transform 1 0 756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9769
timestamp 1677622389
transform 1 0 708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9770
timestamp 1677622389
transform 1 0 716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9771
timestamp 1677622389
transform 1 0 732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9772
timestamp 1677622389
transform 1 0 748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9773
timestamp 1677622389
transform 1 0 756 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8552
timestamp 1677622389
transform 1 0 756 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9774
timestamp 1677622389
transform 1 0 780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8379
timestamp 1677622389
transform 1 0 828 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8410
timestamp 1677622389
transform 1 0 820 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8411
timestamp 1677622389
transform 1 0 860 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8444
timestamp 1677622389
transform 1 0 836 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8498
timestamp 1677622389
transform 1 0 812 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9620
timestamp 1677622389
transform 1 0 820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9621
timestamp 1677622389
transform 1 0 836 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9622
timestamp 1677622389
transform 1 0 860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9775
timestamp 1677622389
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9776
timestamp 1677622389
transform 1 0 828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9777
timestamp 1677622389
transform 1 0 836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9778
timestamp 1677622389
transform 1 0 852 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8600
timestamp 1677622389
transform 1 0 836 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9623
timestamp 1677622389
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9779
timestamp 1677622389
transform 1 0 876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9780
timestamp 1677622389
transform 1 0 892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9781
timestamp 1677622389
transform 1 0 900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8553
timestamp 1677622389
transform 1 0 876 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8554
timestamp 1677622389
transform 1 0 900 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8380
timestamp 1677622389
transform 1 0 932 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8445
timestamp 1677622389
transform 1 0 924 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9624
timestamp 1677622389
transform 1 0 916 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8387
timestamp 1677622389
transform 1 0 972 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8446
timestamp 1677622389
transform 1 0 964 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9625
timestamp 1677622389
transform 1 0 940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9626
timestamp 1677622389
transform 1 0 956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9627
timestamp 1677622389
transform 1 0 972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9782
timestamp 1677622389
transform 1 0 932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9783
timestamp 1677622389
transform 1 0 964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9784
timestamp 1677622389
transform 1 0 972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9628
timestamp 1677622389
transform 1 0 988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8530
timestamp 1677622389
transform 1 0 1020 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9897
timestamp 1677622389
transform 1 0 1020 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_8388
timestamp 1677622389
transform 1 0 1092 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8412
timestamp 1677622389
transform 1 0 1100 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9629
timestamp 1677622389
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9630
timestamp 1677622389
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9631
timestamp 1677622389
transform 1 0 1108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9785
timestamp 1677622389
transform 1 0 1076 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8531
timestamp 1677622389
transform 1 0 1084 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8499
timestamp 1677622389
transform 1 0 1116 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9786
timestamp 1677622389
transform 1 0 1100 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8447
timestamp 1677622389
transform 1 0 1132 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9632
timestamp 1677622389
transform 1 0 1132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9633
timestamp 1677622389
transform 1 0 1140 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8381
timestamp 1677622389
transform 1 0 1156 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8413
timestamp 1677622389
transform 1 0 1156 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8375
timestamp 1677622389
transform 1 0 1196 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8389
timestamp 1677622389
transform 1 0 1196 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8390
timestamp 1677622389
transform 1 0 1212 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8448
timestamp 1677622389
transform 1 0 1180 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9634
timestamp 1677622389
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8500
timestamp 1677622389
transform 1 0 1172 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9635
timestamp 1677622389
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9787
timestamp 1677622389
transform 1 0 1148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9788
timestamp 1677622389
transform 1 0 1156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9789
timestamp 1677622389
transform 1 0 1172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9790
timestamp 1677622389
transform 1 0 1180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8555
timestamp 1677622389
transform 1 0 1156 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8391
timestamp 1677622389
transform 1 0 1252 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8449
timestamp 1677622389
transform 1 0 1236 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8450
timestamp 1677622389
transform 1 0 1268 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9636
timestamp 1677622389
transform 1 0 1196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9637
timestamp 1677622389
transform 1 0 1212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9638
timestamp 1677622389
transform 1 0 1236 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8501
timestamp 1677622389
transform 1 0 1244 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9639
timestamp 1677622389
transform 1 0 1252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9640
timestamp 1677622389
transform 1 0 1268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9791
timestamp 1677622389
transform 1 0 1204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9792
timestamp 1677622389
transform 1 0 1220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9793
timestamp 1677622389
transform 1 0 1236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9794
timestamp 1677622389
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9795
timestamp 1677622389
transform 1 0 1260 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8556
timestamp 1677622389
transform 1 0 1204 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8601
timestamp 1677622389
transform 1 0 1236 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8382
timestamp 1677622389
transform 1 0 1308 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8414
timestamp 1677622389
transform 1 0 1316 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8383
timestamp 1677622389
transform 1 0 1372 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8415
timestamp 1677622389
transform 1 0 1340 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9641
timestamp 1677622389
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9796
timestamp 1677622389
transform 1 0 1324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8557
timestamp 1677622389
transform 1 0 1324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8451
timestamp 1677622389
transform 1 0 1364 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9642
timestamp 1677622389
transform 1 0 1340 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8502
timestamp 1677622389
transform 1 0 1356 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9643
timestamp 1677622389
transform 1 0 1364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9644
timestamp 1677622389
transform 1 0 1380 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8503
timestamp 1677622389
transform 1 0 1388 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9797
timestamp 1677622389
transform 1 0 1348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9798
timestamp 1677622389
transform 1 0 1356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9799
timestamp 1677622389
transform 1 0 1372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9800
timestamp 1677622389
transform 1 0 1380 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8558
timestamp 1677622389
transform 1 0 1380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8452
timestamp 1677622389
transform 1 0 1404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8416
timestamp 1677622389
transform 1 0 1436 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8453
timestamp 1677622389
transform 1 0 1444 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9645
timestamp 1677622389
transform 1 0 1404 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8504
timestamp 1677622389
transform 1 0 1412 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9646
timestamp 1677622389
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8505
timestamp 1677622389
transform 1 0 1428 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8376
timestamp 1677622389
transform 1 0 1468 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8392
timestamp 1677622389
transform 1 0 1468 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8417
timestamp 1677622389
transform 1 0 1460 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9647
timestamp 1677622389
transform 1 0 1436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9648
timestamp 1677622389
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9649
timestamp 1677622389
transform 1 0 1460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9801
timestamp 1677622389
transform 1 0 1404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9802
timestamp 1677622389
transform 1 0 1428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9803
timestamp 1677622389
transform 1 0 1436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9804
timestamp 1677622389
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8418
timestamp 1677622389
transform 1 0 1492 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8454
timestamp 1677622389
transform 1 0 1516 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9650
timestamp 1677622389
transform 1 0 1500 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8506
timestamp 1677622389
transform 1 0 1508 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9651
timestamp 1677622389
transform 1 0 1516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9805
timestamp 1677622389
transform 1 0 1508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9806
timestamp 1677622389
transform 1 0 1516 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8559
timestamp 1677622389
transform 1 0 1500 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8560
timestamp 1677622389
transform 1 0 1516 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8602
timestamp 1677622389
transform 1 0 1508 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9652
timestamp 1677622389
transform 1 0 1572 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8507
timestamp 1677622389
transform 1 0 1580 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9807
timestamp 1677622389
transform 1 0 1580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9653
timestamp 1677622389
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9808
timestamp 1677622389
transform 1 0 1636 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8561
timestamp 1677622389
transform 1 0 1636 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8455
timestamp 1677622389
transform 1 0 1668 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9654
timestamp 1677622389
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8532
timestamp 1677622389
transform 1 0 1652 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9655
timestamp 1677622389
transform 1 0 1684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9809
timestamp 1677622389
transform 1 0 1660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9810
timestamp 1677622389
transform 1 0 1676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9811
timestamp 1677622389
transform 1 0 1684 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8562
timestamp 1677622389
transform 1 0 1684 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8603
timestamp 1677622389
transform 1 0 1676 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9656
timestamp 1677622389
transform 1 0 1716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9657
timestamp 1677622389
transform 1 0 1732 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8533
timestamp 1677622389
transform 1 0 1716 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8456
timestamp 1677622389
transform 1 0 1756 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8508
timestamp 1677622389
transform 1 0 1764 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8419
timestamp 1677622389
transform 1 0 1780 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9658
timestamp 1677622389
transform 1 0 1772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9812
timestamp 1677622389
transform 1 0 1748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9813
timestamp 1677622389
transform 1 0 1756 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8563
timestamp 1677622389
transform 1 0 1748 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8534
timestamp 1677622389
transform 1 0 1772 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9583
timestamp 1677622389
transform 1 0 1780 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8393
timestamp 1677622389
transform 1 0 1820 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9659
timestamp 1677622389
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9660
timestamp 1677622389
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9814
timestamp 1677622389
transform 1 0 1788 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8535
timestamp 1677622389
transform 1 0 1804 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9815
timestamp 1677622389
transform 1 0 1812 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8564
timestamp 1677622389
transform 1 0 1812 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8509
timestamp 1677622389
transform 1 0 1828 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9816
timestamp 1677622389
transform 1 0 1828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9661
timestamp 1677622389
transform 1 0 1860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9817
timestamp 1677622389
transform 1 0 1868 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8604
timestamp 1677622389
transform 1 0 1868 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8536
timestamp 1677622389
transform 1 0 1884 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8457
timestamp 1677622389
transform 1 0 1924 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8420
timestamp 1677622389
transform 1 0 1956 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9662
timestamp 1677622389
transform 1 0 1924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9663
timestamp 1677622389
transform 1 0 1940 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8510
timestamp 1677622389
transform 1 0 1948 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9664
timestamp 1677622389
transform 1 0 1956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9818
timestamp 1677622389
transform 1 0 1932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9819
timestamp 1677622389
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9820
timestamp 1677622389
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9665
timestamp 1677622389
transform 1 0 1988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8458
timestamp 1677622389
transform 1 0 2012 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9821
timestamp 1677622389
transform 1 0 2004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9666
timestamp 1677622389
transform 1 0 2012 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8394
timestamp 1677622389
transform 1 0 2068 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9667
timestamp 1677622389
transform 1 0 2052 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8511
timestamp 1677622389
transform 1 0 2060 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9668
timestamp 1677622389
transform 1 0 2068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9822
timestamp 1677622389
transform 1 0 2044 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8537
timestamp 1677622389
transform 1 0 2052 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9823
timestamp 1677622389
transform 1 0 2060 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8512
timestamp 1677622389
transform 1 0 2076 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9824
timestamp 1677622389
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8605
timestamp 1677622389
transform 1 0 2068 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9669
timestamp 1677622389
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9670
timestamp 1677622389
transform 1 0 2116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9671
timestamp 1677622389
transform 1 0 2172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9825
timestamp 1677622389
transform 1 0 2212 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8565
timestamp 1677622389
transform 1 0 2212 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9672
timestamp 1677622389
transform 1 0 2236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9673
timestamp 1677622389
transform 1 0 2300 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8538
timestamp 1677622389
transform 1 0 2276 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9826
timestamp 1677622389
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8566
timestamp 1677622389
transform 1 0 2244 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8567
timestamp 1677622389
transform 1 0 2324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8459
timestamp 1677622389
transform 1 0 2412 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9674
timestamp 1677622389
transform 1 0 2364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9675
timestamp 1677622389
transform 1 0 2412 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8539
timestamp 1677622389
transform 1 0 2364 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9827
timestamp 1677622389
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8568
timestamp 1677622389
transform 1 0 2444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8606
timestamp 1677622389
transform 1 0 2372 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8569
timestamp 1677622389
transform 1 0 2468 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8460
timestamp 1677622389
transform 1 0 2516 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9676
timestamp 1677622389
transform 1 0 2516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9828
timestamp 1677622389
transform 1 0 2492 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8570
timestamp 1677622389
transform 1 0 2492 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9677
timestamp 1677622389
transform 1 0 2580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9678
timestamp 1677622389
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9829
timestamp 1677622389
transform 1 0 2580 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8421
timestamp 1677622389
transform 1 0 2620 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9679
timestamp 1677622389
transform 1 0 2620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9830
timestamp 1677622389
transform 1 0 2604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9831
timestamp 1677622389
transform 1 0 2628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9832
timestamp 1677622389
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9898
timestamp 1677622389
transform 1 0 2620 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_9680
timestamp 1677622389
transform 1 0 2652 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8540
timestamp 1677622389
transform 1 0 2652 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8422
timestamp 1677622389
transform 1 0 2700 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8423
timestamp 1677622389
transform 1 0 2716 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8461
timestamp 1677622389
transform 1 0 2684 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9584
timestamp 1677622389
transform 1 0 2700 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9681
timestamp 1677622389
transform 1 0 2676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9682
timestamp 1677622389
transform 1 0 2684 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8462
timestamp 1677622389
transform 1 0 2724 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9683
timestamp 1677622389
transform 1 0 2716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9684
timestamp 1677622389
transform 1 0 2724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9833
timestamp 1677622389
transform 1 0 2708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9834
timestamp 1677622389
transform 1 0 2724 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8607
timestamp 1677622389
transform 1 0 2724 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8463
timestamp 1677622389
transform 1 0 2780 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9685
timestamp 1677622389
transform 1 0 2748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9686
timestamp 1677622389
transform 1 0 2772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9835
timestamp 1677622389
transform 1 0 2764 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8541
timestamp 1677622389
transform 1 0 2772 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9836
timestamp 1677622389
transform 1 0 2780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8571
timestamp 1677622389
transform 1 0 2764 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9687
timestamp 1677622389
transform 1 0 2796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9688
timestamp 1677622389
transform 1 0 2804 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8542
timestamp 1677622389
transform 1 0 2796 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8572
timestamp 1677622389
transform 1 0 2804 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9689
timestamp 1677622389
transform 1 0 2820 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8608
timestamp 1677622389
transform 1 0 2820 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8513
timestamp 1677622389
transform 1 0 2836 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8424
timestamp 1677622389
transform 1 0 2868 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9690
timestamp 1677622389
transform 1 0 2868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9691
timestamp 1677622389
transform 1 0 2884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9837
timestamp 1677622389
transform 1 0 2836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9838
timestamp 1677622389
transform 1 0 2844 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8543
timestamp 1677622389
transform 1 0 2852 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9839
timestamp 1677622389
transform 1 0 2860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9840
timestamp 1677622389
transform 1 0 2876 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8573
timestamp 1677622389
transform 1 0 2844 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9692
timestamp 1677622389
transform 1 0 2892 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8574
timestamp 1677622389
transform 1 0 2884 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8609
timestamp 1677622389
transform 1 0 2860 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9841
timestamp 1677622389
transform 1 0 2900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8610
timestamp 1677622389
transform 1 0 2908 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8464
timestamp 1677622389
transform 1 0 2916 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9842
timestamp 1677622389
transform 1 0 2916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9843
timestamp 1677622389
transform 1 0 2924 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8575
timestamp 1677622389
transform 1 0 2924 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8465
timestamp 1677622389
transform 1 0 2940 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9693
timestamp 1677622389
transform 1 0 2932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9694
timestamp 1677622389
transform 1 0 2940 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8576
timestamp 1677622389
transform 1 0 2948 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8514
timestamp 1677622389
transform 1 0 2980 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9695
timestamp 1677622389
transform 1 0 2988 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9696
timestamp 1677622389
transform 1 0 3004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9844
timestamp 1677622389
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9845
timestamp 1677622389
transform 1 0 2996 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8577
timestamp 1677622389
transform 1 0 3004 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8611
timestamp 1677622389
transform 1 0 2980 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9846
timestamp 1677622389
transform 1 0 3028 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8395
timestamp 1677622389
transform 1 0 3068 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9697
timestamp 1677622389
transform 1 0 3068 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8425
timestamp 1677622389
transform 1 0 3156 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9698
timestamp 1677622389
transform 1 0 3092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9699
timestamp 1677622389
transform 1 0 3132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9847
timestamp 1677622389
transform 1 0 3108 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8578
timestamp 1677622389
transform 1 0 3108 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8579
timestamp 1677622389
transform 1 0 3172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8466
timestamp 1677622389
transform 1 0 3196 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9700
timestamp 1677622389
transform 1 0 3196 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8426
timestamp 1677622389
transform 1 0 3236 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9701
timestamp 1677622389
transform 1 0 3236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9848
timestamp 1677622389
transform 1 0 3212 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8580
timestamp 1677622389
transform 1 0 3212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8581
timestamp 1677622389
transform 1 0 3284 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9702
timestamp 1677622389
transform 1 0 3308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9703
timestamp 1677622389
transform 1 0 3316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9704
timestamp 1677622389
transform 1 0 3372 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8582
timestamp 1677622389
transform 1 0 3308 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9849
timestamp 1677622389
transform 1 0 3396 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8612
timestamp 1677622389
transform 1 0 3316 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8467
timestamp 1677622389
transform 1 0 3412 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9850
timestamp 1677622389
transform 1 0 3412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8427
timestamp 1677622389
transform 1 0 3476 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9585
timestamp 1677622389
transform 1 0 3468 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8396
timestamp 1677622389
transform 1 0 3508 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9586
timestamp 1677622389
transform 1 0 3484 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9587
timestamp 1677622389
transform 1 0 3500 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9705
timestamp 1677622389
transform 1 0 3476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9851
timestamp 1677622389
transform 1 0 3468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8583
timestamp 1677622389
transform 1 0 3468 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9706
timestamp 1677622389
transform 1 0 3492 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8515
timestamp 1677622389
transform 1 0 3500 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9707
timestamp 1677622389
transform 1 0 3508 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8544
timestamp 1677622389
transform 1 0 3492 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8397
timestamp 1677622389
transform 1 0 3532 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8516
timestamp 1677622389
transform 1 0 3524 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9708
timestamp 1677622389
transform 1 0 3532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9852
timestamp 1677622389
transform 1 0 3524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8517
timestamp 1677622389
transform 1 0 3572 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9853
timestamp 1677622389
transform 1 0 3572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9854
timestamp 1677622389
transform 1 0 3580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9709
timestamp 1677622389
transform 1 0 3596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9855
timestamp 1677622389
transform 1 0 3604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9710
timestamp 1677622389
transform 1 0 3620 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8468
timestamp 1677622389
transform 1 0 3652 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9711
timestamp 1677622389
transform 1 0 3652 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8518
timestamp 1677622389
transform 1 0 3660 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9856
timestamp 1677622389
transform 1 0 3628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9857
timestamp 1677622389
transform 1 0 3644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8545
timestamp 1677622389
transform 1 0 3652 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8584
timestamp 1677622389
transform 1 0 3628 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8469
timestamp 1677622389
transform 1 0 3692 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8519
timestamp 1677622389
transform 1 0 3676 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9712
timestamp 1677622389
transform 1 0 3684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9858
timestamp 1677622389
transform 1 0 3676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9859
timestamp 1677622389
transform 1 0 3692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9860
timestamp 1677622389
transform 1 0 3708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9713
timestamp 1677622389
transform 1 0 3724 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8585
timestamp 1677622389
transform 1 0 3708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8520
timestamp 1677622389
transform 1 0 3740 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9861
timestamp 1677622389
transform 1 0 3732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9862
timestamp 1677622389
transform 1 0 3740 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8470
timestamp 1677622389
transform 1 0 3756 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9714
timestamp 1677622389
transform 1 0 3756 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8471
timestamp 1677622389
transform 1 0 3788 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9863
timestamp 1677622389
transform 1 0 3764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9864
timestamp 1677622389
transform 1 0 3780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8586
timestamp 1677622389
transform 1 0 3780 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9715
timestamp 1677622389
transform 1 0 3804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9865
timestamp 1677622389
transform 1 0 3820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9866
timestamp 1677622389
transform 1 0 3828 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8587
timestamp 1677622389
transform 1 0 3828 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8472
timestamp 1677622389
transform 1 0 3844 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8473
timestamp 1677622389
transform 1 0 3876 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9716
timestamp 1677622389
transform 1 0 3844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9717
timestamp 1677622389
transform 1 0 3860 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8521
timestamp 1677622389
transform 1 0 3868 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9718
timestamp 1677622389
transform 1 0 3876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9867
timestamp 1677622389
transform 1 0 3852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9868
timestamp 1677622389
transform 1 0 3868 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9869
timestamp 1677622389
transform 1 0 3916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9870
timestamp 1677622389
transform 1 0 3932 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8588
timestamp 1677622389
transform 1 0 3932 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8428
timestamp 1677622389
transform 1 0 3972 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8474
timestamp 1677622389
transform 1 0 3956 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8475
timestamp 1677622389
transform 1 0 3988 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9719
timestamp 1677622389
transform 1 0 3956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9720
timestamp 1677622389
transform 1 0 3972 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8522
timestamp 1677622389
transform 1 0 3980 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9721
timestamp 1677622389
transform 1 0 3988 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9871
timestamp 1677622389
transform 1 0 3964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9872
timestamp 1677622389
transform 1 0 3980 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8398
timestamp 1677622389
transform 1 0 4012 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8399
timestamp 1677622389
transform 1 0 4044 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9873
timestamp 1677622389
transform 1 0 4004 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8476
timestamp 1677622389
transform 1 0 4092 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9722
timestamp 1677622389
transform 1 0 4044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9723
timestamp 1677622389
transform 1 0 4100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9874
timestamp 1677622389
transform 1 0 4020 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8546
timestamp 1677622389
transform 1 0 4108 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8400
timestamp 1677622389
transform 1 0 4124 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8401
timestamp 1677622389
transform 1 0 4156 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8402
timestamp 1677622389
transform 1 0 4180 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8477
timestamp 1677622389
transform 1 0 4164 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9724
timestamp 1677622389
transform 1 0 4140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9725
timestamp 1677622389
transform 1 0 4148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9726
timestamp 1677622389
transform 1 0 4164 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8523
timestamp 1677622389
transform 1 0 4172 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9727
timestamp 1677622389
transform 1 0 4180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9875
timestamp 1677622389
transform 1 0 4132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9876
timestamp 1677622389
transform 1 0 4140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9877
timestamp 1677622389
transform 1 0 4156 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8547
timestamp 1677622389
transform 1 0 4164 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9878
timestamp 1677622389
transform 1 0 4172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8589
timestamp 1677622389
transform 1 0 4148 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8478
timestamp 1677622389
transform 1 0 4252 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8524
timestamp 1677622389
transform 1 0 4204 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8429
timestamp 1677622389
transform 1 0 4300 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8430
timestamp 1677622389
transform 1 0 4332 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9728
timestamp 1677622389
transform 1 0 4252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9729
timestamp 1677622389
transform 1 0 4292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9730
timestamp 1677622389
transform 1 0 4300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9731
timestamp 1677622389
transform 1 0 4316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9732
timestamp 1677622389
transform 1 0 4332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9879
timestamp 1677622389
transform 1 0 4188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9880
timestamp 1677622389
transform 1 0 4204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9881
timestamp 1677622389
transform 1 0 4292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9882
timestamp 1677622389
transform 1 0 4308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9883
timestamp 1677622389
transform 1 0 4324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8590
timestamp 1677622389
transform 1 0 4188 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8591
timestamp 1677622389
transform 1 0 4244 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8613
timestamp 1677622389
transform 1 0 4292 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8592
timestamp 1677622389
transform 1 0 4324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8479
timestamp 1677622389
transform 1 0 4364 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9884
timestamp 1677622389
transform 1 0 4356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9885
timestamp 1677622389
transform 1 0 4364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8614
timestamp 1677622389
transform 1 0 4364 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9733
timestamp 1677622389
transform 1 0 4396 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8480
timestamp 1677622389
transform 1 0 4412 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8481
timestamp 1677622389
transform 1 0 4444 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9734
timestamp 1677622389
transform 1 0 4412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9735
timestamp 1677622389
transform 1 0 4428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9736
timestamp 1677622389
transform 1 0 4444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9886
timestamp 1677622389
transform 1 0 4420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9887
timestamp 1677622389
transform 1 0 4436 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8593
timestamp 1677622389
transform 1 0 4436 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8482
timestamp 1677622389
transform 1 0 4468 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8483
timestamp 1677622389
transform 1 0 4492 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8525
timestamp 1677622389
transform 1 0 4468 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8484
timestamp 1677622389
transform 1 0 4604 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8485
timestamp 1677622389
transform 1 0 4628 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9737
timestamp 1677622389
transform 1 0 4492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9738
timestamp 1677622389
transform 1 0 4548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9739
timestamp 1677622389
transform 1 0 4564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9740
timestamp 1677622389
transform 1 0 4580 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8526
timestamp 1677622389
transform 1 0 4596 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9741
timestamp 1677622389
transform 1 0 4604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9742
timestamp 1677622389
transform 1 0 4620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9888
timestamp 1677622389
transform 1 0 4452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9889
timestamp 1677622389
transform 1 0 4468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9890
timestamp 1677622389
transform 1 0 4556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9891
timestamp 1677622389
transform 1 0 4572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9892
timestamp 1677622389
transform 1 0 4596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9893
timestamp 1677622389
transform 1 0 4612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9894
timestamp 1677622389
transform 1 0 4628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8594
timestamp 1677622389
transform 1 0 4556 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8615
timestamp 1677622389
transform 1 0 4468 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8616
timestamp 1677622389
transform 1 0 4492 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8595
timestamp 1677622389
transform 1 0 4596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8596
timestamp 1677622389
transform 1 0 4612 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8527
timestamp 1677622389
transform 1 0 4660 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9743
timestamp 1677622389
transform 1 0 4700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9895
timestamp 1677622389
transform 1 0 4676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8597
timestamp 1677622389
transform 1 0 4700 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8617
timestamp 1677622389
transform 1 0 4676 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8486
timestamp 1677622389
transform 1 0 4772 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9744
timestamp 1677622389
transform 1 0 4764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9745
timestamp 1677622389
transform 1 0 4772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9896
timestamp 1677622389
transform 1 0 4780 0 1 205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_90
timestamp 1677622389
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_10559
timestamp 1677622389
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_10560
timestamp 1677622389
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_10561
timestamp 1677622389
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_10562
timestamp 1677622389
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_10563
timestamp 1677622389
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_10564
timestamp 1677622389
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_10565
timestamp 1677622389
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_10566
timestamp 1677622389
transform 1 0 128 0 1 170
box -8 -3 16 105
use INVX2  INVX2_683
timestamp 1677622389
transform -1 0 152 0 1 170
box -9 -3 26 105
use FILL  FILL_10567
timestamp 1677622389
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_10568
timestamp 1677622389
transform 1 0 160 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_398
timestamp 1677622389
transform -1 0 208 0 1 170
box -8 -3 46 105
use FILL  FILL_10569
timestamp 1677622389
transform 1 0 208 0 1 170
box -8 -3 16 105
use INVX2  INVX2_684
timestamp 1677622389
transform -1 0 232 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_399
timestamp 1677622389
transform 1 0 232 0 1 170
box -8 -3 46 105
use FILL  FILL_10570
timestamp 1677622389
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_10573
timestamp 1677622389
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_10575
timestamp 1677622389
transform 1 0 288 0 1 170
box -8 -3 16 105
use INVX2  INVX2_685
timestamp 1677622389
transform 1 0 296 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_400
timestamp 1677622389
transform 1 0 312 0 1 170
box -8 -3 46 105
use FILL  FILL_10576
timestamp 1677622389
transform 1 0 352 0 1 170
box -8 -3 16 105
use FILL  FILL_10577
timestamp 1677622389
transform 1 0 360 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_401
timestamp 1677622389
transform 1 0 368 0 1 170
box -8 -3 46 105
use INVX2  INVX2_686
timestamp 1677622389
transform 1 0 408 0 1 170
box -9 -3 26 105
use FILL  FILL_10578
timestamp 1677622389
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_10579
timestamp 1677622389
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_10580
timestamp 1677622389
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_10581
timestamp 1677622389
transform 1 0 448 0 1 170
box -8 -3 16 105
use INVX2  INVX2_687
timestamp 1677622389
transform 1 0 456 0 1 170
box -9 -3 26 105
use FILL  FILL_10582
timestamp 1677622389
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_10583
timestamp 1677622389
transform 1 0 480 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8618
timestamp 1677622389
transform 1 0 516 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_402
timestamp 1677622389
transform 1 0 488 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_432
timestamp 1677622389
transform 1 0 528 0 1 170
box -8 -3 46 105
use FILL  FILL_10584
timestamp 1677622389
transform 1 0 568 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8619
timestamp 1677622389
transform 1 0 612 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_403
timestamp 1677622389
transform 1 0 576 0 1 170
box -8 -3 46 105
use FILL  FILL_10585
timestamp 1677622389
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_10592
timestamp 1677622389
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_10594
timestamp 1677622389
transform 1 0 632 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_404
timestamp 1677622389
transform 1 0 640 0 1 170
box -8 -3 46 105
use INVX2  INVX2_688
timestamp 1677622389
transform 1 0 680 0 1 170
box -9 -3 26 105
use FILL  FILL_10595
timestamp 1677622389
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_10596
timestamp 1677622389
transform 1 0 704 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_433
timestamp 1677622389
transform 1 0 712 0 1 170
box -8 -3 46 105
use FILL  FILL_10597
timestamp 1677622389
transform 1 0 752 0 1 170
box -8 -3 16 105
use FILL  FILL_10598
timestamp 1677622389
transform 1 0 760 0 1 170
box -8 -3 16 105
use FILL  FILL_10599
timestamp 1677622389
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_10600
timestamp 1677622389
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_10601
timestamp 1677622389
transform 1 0 784 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_434
timestamp 1677622389
transform 1 0 792 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_435
timestamp 1677622389
transform 1 0 832 0 1 170
box -8 -3 46 105
use FILL  FILL_10602
timestamp 1677622389
transform 1 0 872 0 1 170
box -8 -3 16 105
use INVX2  INVX2_689
timestamp 1677622389
transform -1 0 896 0 1 170
box -9 -3 26 105
use FILL  FILL_10603
timestamp 1677622389
transform 1 0 896 0 1 170
box -8 -3 16 105
use FILL  FILL_10604
timestamp 1677622389
transform 1 0 904 0 1 170
box -8 -3 16 105
use FILL  FILL_10605
timestamp 1677622389
transform 1 0 912 0 1 170
box -8 -3 16 105
use FILL  FILL_10613
timestamp 1677622389
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_10614
timestamp 1677622389
transform 1 0 928 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_406
timestamp 1677622389
transform -1 0 976 0 1 170
box -8 -3 46 105
use FILL  FILL_10615
timestamp 1677622389
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_10616
timestamp 1677622389
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_10617
timestamp 1677622389
transform 1 0 992 0 1 170
box -8 -3 16 105
use INVX2  INVX2_690
timestamp 1677622389
transform 1 0 1000 0 1 170
box -9 -3 26 105
use FILL  FILL_10618
timestamp 1677622389
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_10619
timestamp 1677622389
transform 1 0 1024 0 1 170
box -8 -3 16 105
use FILL  FILL_10622
timestamp 1677622389
transform 1 0 1032 0 1 170
box -8 -3 16 105
use FILL  FILL_10624
timestamp 1677622389
transform 1 0 1040 0 1 170
box -8 -3 16 105
use FILL  FILL_10626
timestamp 1677622389
transform 1 0 1048 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_119
timestamp 1677622389
transform 1 0 1056 0 1 170
box -8 -3 32 105
use FILL  FILL_10627
timestamp 1677622389
transform 1 0 1080 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_407
timestamp 1677622389
transform 1 0 1088 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_8620
timestamp 1677622389
transform 1 0 1140 0 1 175
box -3 -3 3 3
use FILL  FILL_10628
timestamp 1677622389
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_10629
timestamp 1677622389
transform 1 0 1136 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_408
timestamp 1677622389
transform 1 0 1144 0 1 170
box -8 -3 46 105
use INVX2  INVX2_691
timestamp 1677622389
transform 1 0 1184 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_436
timestamp 1677622389
transform -1 0 1240 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_437
timestamp 1677622389
transform -1 0 1280 0 1 170
box -8 -3 46 105
use FILL  FILL_10630
timestamp 1677622389
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_10635
timestamp 1677622389
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_10636
timestamp 1677622389
transform 1 0 1296 0 1 170
box -8 -3 16 105
use FILL  FILL_10637
timestamp 1677622389
transform 1 0 1304 0 1 170
box -8 -3 16 105
use FILL  FILL_10638
timestamp 1677622389
transform 1 0 1312 0 1 170
box -8 -3 16 105
use FILL  FILL_10639
timestamp 1677622389
transform 1 0 1320 0 1 170
box -8 -3 16 105
use INVX2  INVX2_693
timestamp 1677622389
transform -1 0 1344 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_409
timestamp 1677622389
transform -1 0 1384 0 1 170
box -8 -3 46 105
use FILL  FILL_10640
timestamp 1677622389
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_10642
timestamp 1677622389
transform 1 0 1392 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8621
timestamp 1677622389
transform 1 0 1412 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_410
timestamp 1677622389
transform -1 0 1440 0 1 170
box -8 -3 46 105
use INVX2  INVX2_694
timestamp 1677622389
transform 1 0 1440 0 1 170
box -9 -3 26 105
use FILL  FILL_10643
timestamp 1677622389
transform 1 0 1456 0 1 170
box -8 -3 16 105
use FILL  FILL_10644
timestamp 1677622389
transform 1 0 1464 0 1 170
box -8 -3 16 105
use FILL  FILL_10645
timestamp 1677622389
transform 1 0 1472 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_411
timestamp 1677622389
transform 1 0 1480 0 1 170
box -8 -3 46 105
use FILL  FILL_10646
timestamp 1677622389
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_10647
timestamp 1677622389
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_10648
timestamp 1677622389
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_10649
timestamp 1677622389
transform 1 0 1544 0 1 170
box -8 -3 16 105
use INVX2  INVX2_695
timestamp 1677622389
transform 1 0 1552 0 1 170
box -9 -3 26 105
use FILL  FILL_10650
timestamp 1677622389
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_10651
timestamp 1677622389
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_10652
timestamp 1677622389
transform 1 0 1584 0 1 170
box -8 -3 16 105
use INVX2  INVX2_696
timestamp 1677622389
transform 1 0 1592 0 1 170
box -9 -3 26 105
use FILL  FILL_10653
timestamp 1677622389
transform 1 0 1608 0 1 170
box -8 -3 16 105
use FILL  FILL_10654
timestamp 1677622389
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_10660
timestamp 1677622389
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_10661
timestamp 1677622389
transform 1 0 1632 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_438
timestamp 1677622389
transform -1 0 1680 0 1 170
box -8 -3 46 105
use FILL  FILL_10662
timestamp 1677622389
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_10663
timestamp 1677622389
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_10664
timestamp 1677622389
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_10665
timestamp 1677622389
transform 1 0 1704 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_412
timestamp 1677622389
transform -1 0 1752 0 1 170
box -8 -3 46 105
use FILL  FILL_10666
timestamp 1677622389
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_10670
timestamp 1677622389
transform 1 0 1760 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8622
timestamp 1677622389
transform 1 0 1780 0 1 175
box -3 -3 3 3
use FILL  FILL_10672
timestamp 1677622389
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_10674
timestamp 1677622389
transform 1 0 1776 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_413
timestamp 1677622389
transform -1 0 1824 0 1 170
box -8 -3 46 105
use FILL  FILL_10675
timestamp 1677622389
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_10676
timestamp 1677622389
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_10677
timestamp 1677622389
transform 1 0 1840 0 1 170
box -8 -3 16 105
use INVX2  INVX2_698
timestamp 1677622389
transform 1 0 1848 0 1 170
box -9 -3 26 105
use FILL  FILL_10678
timestamp 1677622389
transform 1 0 1864 0 1 170
box -8 -3 16 105
use FILL  FILL_10679
timestamp 1677622389
transform 1 0 1872 0 1 170
box -8 -3 16 105
use FILL  FILL_10680
timestamp 1677622389
transform 1 0 1880 0 1 170
box -8 -3 16 105
use FILL  FILL_10681
timestamp 1677622389
transform 1 0 1888 0 1 170
box -8 -3 16 105
use FILL  FILL_10682
timestamp 1677622389
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_10685
timestamp 1677622389
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_10687
timestamp 1677622389
transform 1 0 1912 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_414
timestamp 1677622389
transform -1 0 1960 0 1 170
box -8 -3 46 105
use FILL  FILL_10688
timestamp 1677622389
transform 1 0 1960 0 1 170
box -8 -3 16 105
use FILL  FILL_10689
timestamp 1677622389
transform 1 0 1968 0 1 170
box -8 -3 16 105
use FILL  FILL_10690
timestamp 1677622389
transform 1 0 1976 0 1 170
box -8 -3 16 105
use INVX2  INVX2_700
timestamp 1677622389
transform 1 0 1984 0 1 170
box -9 -3 26 105
use FILL  FILL_10691
timestamp 1677622389
transform 1 0 2000 0 1 170
box -8 -3 16 105
use FILL  FILL_10692
timestamp 1677622389
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_10693
timestamp 1677622389
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_10694
timestamp 1677622389
transform 1 0 2024 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_415
timestamp 1677622389
transform -1 0 2072 0 1 170
box -8 -3 46 105
use FILL  FILL_10695
timestamp 1677622389
transform 1 0 2072 0 1 170
box -8 -3 16 105
use FILL  FILL_10696
timestamp 1677622389
transform 1 0 2080 0 1 170
box -8 -3 16 105
use FILL  FILL_10697
timestamp 1677622389
transform 1 0 2088 0 1 170
box -8 -3 16 105
use INVX2  INVX2_701
timestamp 1677622389
transform 1 0 2096 0 1 170
box -9 -3 26 105
use FILL  FILL_10698
timestamp 1677622389
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_10699
timestamp 1677622389
transform 1 0 2120 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_614
timestamp 1677622389
transform -1 0 2224 0 1 170
box -8 -3 104 105
use FILL  FILL_10700
timestamp 1677622389
transform 1 0 2224 0 1 170
box -8 -3 16 105
use FILL  FILL_10701
timestamp 1677622389
transform 1 0 2232 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8623
timestamp 1677622389
transform 1 0 2300 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_8624
timestamp 1677622389
transform 1 0 2332 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_615
timestamp 1677622389
transform -1 0 2336 0 1 170
box -8 -3 104 105
use FILL  FILL_10702
timestamp 1677622389
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_10703
timestamp 1677622389
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_10704
timestamp 1677622389
transform 1 0 2352 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_616
timestamp 1677622389
transform -1 0 2456 0 1 170
box -8 -3 104 105
use FILL  FILL_10705
timestamp 1677622389
transform 1 0 2456 0 1 170
box -8 -3 16 105
use FILL  FILL_10706
timestamp 1677622389
transform 1 0 2464 0 1 170
box -8 -3 16 105
use FILL  FILL_10707
timestamp 1677622389
transform 1 0 2472 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_617
timestamp 1677622389
transform 1 0 2480 0 1 170
box -8 -3 104 105
use FILL  FILL_10708
timestamp 1677622389
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_10733
timestamp 1677622389
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_10735
timestamp 1677622389
transform 1 0 2592 0 1 170
box -8 -3 16 105
use INVX2  INVX2_702
timestamp 1677622389
transform 1 0 2600 0 1 170
box -9 -3 26 105
use NOR2X1  NOR2X1_120
timestamp 1677622389
transform 1 0 2616 0 1 170
box -8 -3 32 105
use FILL  FILL_10736
timestamp 1677622389
transform 1 0 2640 0 1 170
box -8 -3 16 105
use INVX2  INVX2_703
timestamp 1677622389
transform 1 0 2648 0 1 170
box -9 -3 26 105
use FILL  FILL_10737
timestamp 1677622389
transform 1 0 2664 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_185
timestamp 1677622389
transform 1 0 2672 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_8625
timestamp 1677622389
transform 1 0 2724 0 1 175
box -3 -3 3 3
use NAND2X1  NAND2X1_57
timestamp 1677622389
transform -1 0 2728 0 1 170
box -8 -3 32 105
use FILL  FILL_10738
timestamp 1677622389
transform 1 0 2728 0 1 170
box -8 -3 16 105
use INVX2  INVX2_704
timestamp 1677622389
transform -1 0 2752 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_416
timestamp 1677622389
transform -1 0 2792 0 1 170
box -8 -3 46 105
use FILL  FILL_10739
timestamp 1677622389
transform 1 0 2792 0 1 170
box -8 -3 16 105
use FILL  FILL_10740
timestamp 1677622389
transform 1 0 2800 0 1 170
box -8 -3 16 105
use INVX2  INVX2_705
timestamp 1677622389
transform -1 0 2824 0 1 170
box -9 -3 26 105
use FILL  FILL_10741
timestamp 1677622389
transform 1 0 2824 0 1 170
box -8 -3 16 105
use FILL  FILL_10743
timestamp 1677622389
transform 1 0 2832 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_439
timestamp 1677622389
transform 1 0 2840 0 1 170
box -8 -3 46 105
use INVX2  INVX2_707
timestamp 1677622389
transform -1 0 2896 0 1 170
box -9 -3 26 105
use FILL  FILL_10744
timestamp 1677622389
transform 1 0 2896 0 1 170
box -8 -3 16 105
use INVX2  INVX2_708
timestamp 1677622389
transform -1 0 2920 0 1 170
box -9 -3 26 105
use INVX2  INVX2_709
timestamp 1677622389
transform 1 0 2920 0 1 170
box -9 -3 26 105
use FILL  FILL_10745
timestamp 1677622389
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_10746
timestamp 1677622389
transform 1 0 2944 0 1 170
box -8 -3 16 105
use FILL  FILL_10747
timestamp 1677622389
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_10748
timestamp 1677622389
transform 1 0 2960 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_417
timestamp 1677622389
transform 1 0 2968 0 1 170
box -8 -3 46 105
use FILL  FILL_10752
timestamp 1677622389
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_10754
timestamp 1677622389
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_10756
timestamp 1677622389
transform 1 0 3024 0 1 170
box -8 -3 16 105
use BUFX2  BUFX2_113
timestamp 1677622389
transform -1 0 3056 0 1 170
box -5 -3 28 105
use FILL  FILL_10757
timestamp 1677622389
transform 1 0 3056 0 1 170
box -8 -3 16 105
use FILL  FILL_10758
timestamp 1677622389
transform 1 0 3064 0 1 170
box -8 -3 16 105
use BUFX2  BUFX2_114
timestamp 1677622389
transform -1 0 3096 0 1 170
box -5 -3 28 105
use M3_M2  M3_M2_8626
timestamp 1677622389
transform 1 0 3132 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_625
timestamp 1677622389
transform 1 0 3096 0 1 170
box -8 -3 104 105
use FILL  FILL_10759
timestamp 1677622389
transform 1 0 3192 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_626
timestamp 1677622389
transform 1 0 3200 0 1 170
box -8 -3 104 105
use FILL  FILL_10760
timestamp 1677622389
transform 1 0 3296 0 1 170
box -8 -3 16 105
use FILL  FILL_10761
timestamp 1677622389
transform 1 0 3304 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_627
timestamp 1677622389
transform -1 0 3408 0 1 170
box -8 -3 104 105
use FILL  FILL_10762
timestamp 1677622389
transform 1 0 3408 0 1 170
box -8 -3 16 105
use FILL  FILL_10763
timestamp 1677622389
transform 1 0 3416 0 1 170
box -8 -3 16 105
use FILL  FILL_10764
timestamp 1677622389
transform 1 0 3424 0 1 170
box -8 -3 16 105
use FILL  FILL_10765
timestamp 1677622389
transform 1 0 3432 0 1 170
box -8 -3 16 105
use FILL  FILL_10766
timestamp 1677622389
transform 1 0 3440 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_59
timestamp 1677622389
transform 1 0 3448 0 1 170
box -8 -3 32 105
use FILL  FILL_10767
timestamp 1677622389
transform 1 0 3472 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_60
timestamp 1677622389
transform 1 0 3480 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_8627
timestamp 1677622389
transform 1 0 3524 0 1 175
box -3 -3 3 3
use BUFX2  BUFX2_115
timestamp 1677622389
transform 1 0 3504 0 1 170
box -5 -3 28 105
use FILL  FILL_10768
timestamp 1677622389
transform 1 0 3528 0 1 170
box -8 -3 16 105
use FILL  FILL_10769
timestamp 1677622389
transform 1 0 3536 0 1 170
box -8 -3 16 105
use FILL  FILL_10770
timestamp 1677622389
transform 1 0 3544 0 1 170
box -8 -3 16 105
use BUFX2  BUFX2_116
timestamp 1677622389
transform 1 0 3552 0 1 170
box -5 -3 28 105
use INVX2  INVX2_711
timestamp 1677622389
transform 1 0 3576 0 1 170
box -9 -3 26 105
use FILL  FILL_10771
timestamp 1677622389
transform 1 0 3592 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8628
timestamp 1677622389
transform 1 0 3628 0 1 175
box -3 -3 3 3
use INVX2  INVX2_712
timestamp 1677622389
transform 1 0 3600 0 1 170
box -9 -3 26 105
use FILL  FILL_10772
timestamp 1677622389
transform 1 0 3616 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_441
timestamp 1677622389
transform 1 0 3624 0 1 170
box -8 -3 46 105
use FILL  FILL_10773
timestamp 1677622389
transform 1 0 3664 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_442
timestamp 1677622389
transform -1 0 3712 0 1 170
box -8 -3 46 105
use FILL  FILL_10774
timestamp 1677622389
transform 1 0 3712 0 1 170
box -8 -3 16 105
use INVX2  INVX2_713
timestamp 1677622389
transform -1 0 3736 0 1 170
box -9 -3 26 105
use FILL  FILL_10775
timestamp 1677622389
transform 1 0 3736 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_443
timestamp 1677622389
transform -1 0 3784 0 1 170
box -8 -3 46 105
use FILL  FILL_10776
timestamp 1677622389
transform 1 0 3784 0 1 170
box -8 -3 16 105
use FILL  FILL_10777
timestamp 1677622389
transform 1 0 3792 0 1 170
box -8 -3 16 105
use FILL  FILL_10778
timestamp 1677622389
transform 1 0 3800 0 1 170
box -8 -3 16 105
use INVX2  INVX2_714
timestamp 1677622389
transform -1 0 3824 0 1 170
box -9 -3 26 105
use FILL  FILL_10779
timestamp 1677622389
transform 1 0 3824 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_444
timestamp 1677622389
transform 1 0 3832 0 1 170
box -8 -3 46 105
use INVX2  INVX2_715
timestamp 1677622389
transform -1 0 3888 0 1 170
box -9 -3 26 105
use FILL  FILL_10780
timestamp 1677622389
transform 1 0 3888 0 1 170
box -8 -3 16 105
use FILL  FILL_10781
timestamp 1677622389
transform 1 0 3896 0 1 170
box -8 -3 16 105
use FILL  FILL_10782
timestamp 1677622389
transform 1 0 3904 0 1 170
box -8 -3 16 105
use FILL  FILL_10783
timestamp 1677622389
transform 1 0 3912 0 1 170
box -8 -3 16 105
use FILL  FILL_10784
timestamp 1677622389
transform 1 0 3920 0 1 170
box -8 -3 16 105
use FILL  FILL_10800
timestamp 1677622389
transform 1 0 3928 0 1 170
box -8 -3 16 105
use FILL  FILL_10802
timestamp 1677622389
transform 1 0 3936 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_445
timestamp 1677622389
transform 1 0 3944 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_8629
timestamp 1677622389
transform 1 0 4004 0 1 175
box -3 -3 3 3
use INVX2  INVX2_717
timestamp 1677622389
transform -1 0 4000 0 1 170
box -9 -3 26 105
use FILL  FILL_10803
timestamp 1677622389
transform 1 0 4000 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8630
timestamp 1677622389
transform 1 0 4028 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_636
timestamp 1677622389
transform 1 0 4008 0 1 170
box -8 -3 104 105
use INVX2  INVX2_718
timestamp 1677622389
transform -1 0 4120 0 1 170
box -9 -3 26 105
use FILL  FILL_10804
timestamp 1677622389
transform 1 0 4120 0 1 170
box -8 -3 16 105
use FILL  FILL_10805
timestamp 1677622389
transform 1 0 4128 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_446
timestamp 1677622389
transform 1 0 4136 0 1 170
box -8 -3 46 105
use INVX2  INVX2_719
timestamp 1677622389
transform -1 0 4192 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_637
timestamp 1677622389
transform 1 0 4192 0 1 170
box -8 -3 104 105
use OAI22X1  OAI22X1_447
timestamp 1677622389
transform 1 0 4288 0 1 170
box -8 -3 46 105
use INVX2  INVX2_720
timestamp 1677622389
transform -1 0 4344 0 1 170
box -9 -3 26 105
use FILL  FILL_10806
timestamp 1677622389
transform 1 0 4344 0 1 170
box -8 -3 16 105
use FILL  FILL_10807
timestamp 1677622389
transform 1 0 4352 0 1 170
box -8 -3 16 105
use FILL  FILL_10808
timestamp 1677622389
transform 1 0 4360 0 1 170
box -8 -3 16 105
use FILL  FILL_10815
timestamp 1677622389
transform 1 0 4368 0 1 170
box -8 -3 16 105
use FILL  FILL_10817
timestamp 1677622389
transform 1 0 4376 0 1 170
box -8 -3 16 105
use FILL  FILL_10818
timestamp 1677622389
transform 1 0 4384 0 1 170
box -8 -3 16 105
use FILL  FILL_10819
timestamp 1677622389
transform 1 0 4392 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_448
timestamp 1677622389
transform 1 0 4400 0 1 170
box -8 -3 46 105
use INVX2  INVX2_721
timestamp 1677622389
transform -1 0 4456 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_642
timestamp 1677622389
transform 1 0 4456 0 1 170
box -8 -3 104 105
use OAI22X1  OAI22X1_449
timestamp 1677622389
transform -1 0 4592 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_450
timestamp 1677622389
transform 1 0 4592 0 1 170
box -8 -3 46 105
use FILL  FILL_10820
timestamp 1677622389
transform 1 0 4632 0 1 170
box -8 -3 16 105
use FILL  FILL_10821
timestamp 1677622389
transform 1 0 4640 0 1 170
box -8 -3 16 105
use FILL  FILL_10822
timestamp 1677622389
transform 1 0 4648 0 1 170
box -8 -3 16 105
use FILL  FILL_10823
timestamp 1677622389
transform 1 0 4656 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_643
timestamp 1677622389
transform 1 0 4664 0 1 170
box -8 -3 104 105
use FILL  FILL_10824
timestamp 1677622389
transform 1 0 4760 0 1 170
box -8 -3 16 105
use INVX2  INVX2_722
timestamp 1677622389
transform -1 0 4784 0 1 170
box -9 -3 26 105
use FILL  FILL_10825
timestamp 1677622389
transform 1 0 4784 0 1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_91
timestamp 1677622389
transform 1 0 4819 0 1 170
box -10 -3 10 3
use M3_M2  M3_M2_8659
timestamp 1677622389
transform 1 0 84 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9900
timestamp 1677622389
transform 1 0 84 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8660
timestamp 1677622389
transform 1 0 180 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9901
timestamp 1677622389
transform 1 0 180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9958
timestamp 1677622389
transform 1 0 116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9959
timestamp 1677622389
transform 1 0 164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9960
timestamp 1677622389
transform 1 0 220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9961
timestamp 1677622389
transform 1 0 260 0 1 125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_92
timestamp 1677622389
transform 1 0 24 0 1 70
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_599
timestamp 1677622389
transform 1 0 72 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_600
timestamp 1677622389
transform 1 0 168 0 -1 170
box -8 -3 104 105
use FILL  FILL_10571
timestamp 1677622389
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_10572
timestamp 1677622389
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_10574
timestamp 1677622389
transform 1 0 280 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8661
timestamp 1677622389
transform 1 0 300 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8662
timestamp 1677622389
transform 1 0 364 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9902
timestamp 1677622389
transform 1 0 300 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9962
timestamp 1677622389
transform 1 0 324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9963
timestamp 1677622389
transform 1 0 380 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_601
timestamp 1677622389
transform 1 0 288 0 -1 170
box -8 -3 104 105
use FILL  FILL_10586
timestamp 1677622389
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_10587
timestamp 1677622389
transform 1 0 392 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8663
timestamp 1677622389
transform 1 0 412 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9903
timestamp 1677622389
transform 1 0 412 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8631
timestamp 1677622389
transform 1 0 500 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9964
timestamp 1677622389
transform 1 0 436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9965
timestamp 1677622389
transform 1 0 492 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_602
timestamp 1677622389
transform 1 0 400 0 -1 170
box -8 -3 104 105
use FILL  FILL_10588
timestamp 1677622389
transform 1 0 496 0 -1 170
box -8 -3 16 105
use FILL  FILL_10589
timestamp 1677622389
transform 1 0 504 0 -1 170
box -8 -3 16 105
use FILL  FILL_10590
timestamp 1677622389
transform 1 0 512 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8632
timestamp 1677622389
transform 1 0 572 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8664
timestamp 1677622389
transform 1 0 532 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9904
timestamp 1677622389
transform 1 0 532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9966
timestamp 1677622389
transform 1 0 556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9967
timestamp 1677622389
transform 1 0 612 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8707
timestamp 1677622389
transform 1 0 620 0 1 125
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_603
timestamp 1677622389
transform 1 0 520 0 -1 170
box -8 -3 104 105
use FILL  FILL_10591
timestamp 1677622389
transform 1 0 616 0 -1 170
box -8 -3 16 105
use FILL  FILL_10593
timestamp 1677622389
transform 1 0 624 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8633
timestamp 1677622389
transform 1 0 652 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8665
timestamp 1677622389
transform 1 0 644 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8666
timestamp 1677622389
transform 1 0 692 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9905
timestamp 1677622389
transform 1 0 644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9968
timestamp 1677622389
transform 1 0 684 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9969
timestamp 1677622389
transform 1 0 724 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_604
timestamp 1677622389
transform 1 0 632 0 -1 170
box -8 -3 104 105
use FILL  FILL_10606
timestamp 1677622389
transform 1 0 728 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8667
timestamp 1677622389
transform 1 0 748 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9970
timestamp 1677622389
transform 1 0 748 0 1 125
box -2 -2 2 2
use FILL  FILL_10607
timestamp 1677622389
transform 1 0 736 0 -1 170
box -8 -3 16 105
use FILL  FILL_10608
timestamp 1677622389
transform 1 0 744 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8634
timestamp 1677622389
transform 1 0 812 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8643
timestamp 1677622389
transform 1 0 836 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9906
timestamp 1677622389
transform 1 0 836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9971
timestamp 1677622389
transform 1 0 812 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8668
timestamp 1677622389
transform 1 0 852 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9907
timestamp 1677622389
transform 1 0 852 0 1 135
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_605
timestamp 1677622389
transform -1 0 848 0 -1 170
box -8 -3 104 105
use FILL  FILL_10609
timestamp 1677622389
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_10610
timestamp 1677622389
transform 1 0 856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8635
timestamp 1677622389
transform 1 0 884 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8701
timestamp 1677622389
transform 1 0 876 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8644
timestamp 1677622389
transform 1 0 908 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9972
timestamp 1677622389
transform 1 0 876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9973
timestamp 1677622389
transform 1 0 892 0 1 125
box -2 -2 2 2
use FILL  FILL_10611
timestamp 1677622389
transform 1 0 864 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8708
timestamp 1677622389
transform 1 0 900 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8702
timestamp 1677622389
transform 1 0 916 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9908
timestamp 1677622389
transform 1 0 924 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9974
timestamp 1677622389
transform 1 0 908 0 1 125
box -2 -2 2 2
use AOI22X1  AOI22X1_405
timestamp 1677622389
transform -1 0 912 0 -1 170
box -8 -3 46 105
use FILL  FILL_10612
timestamp 1677622389
transform 1 0 912 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8645
timestamp 1677622389
transform 1 0 1012 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9909
timestamp 1677622389
transform 1 0 1012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9975
timestamp 1677622389
transform 1 0 932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9976
timestamp 1677622389
transform 1 0 988 0 1 125
box -2 -2 2 2
use FILL  FILL_10620
timestamp 1677622389
transform 1 0 920 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_606
timestamp 1677622389
transform -1 0 1024 0 -1 170
box -8 -3 104 105
use FILL  FILL_10621
timestamp 1677622389
transform 1 0 1024 0 -1 170
box -8 -3 16 105
use FILL  FILL_10623
timestamp 1677622389
transform 1 0 1032 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8646
timestamp 1677622389
transform 1 0 1076 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8669
timestamp 1677622389
transform 1 0 1052 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9910
timestamp 1677622389
transform 1 0 1052 0 1 135
box -2 -2 2 2
use FILL  FILL_10625
timestamp 1677622389
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8670
timestamp 1677622389
transform 1 0 1108 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9911
timestamp 1677622389
transform 1 0 1076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9977
timestamp 1677622389
transform 1 0 1060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9978
timestamp 1677622389
transform 1 0 1100 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8709
timestamp 1677622389
transform 1 0 1140 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9979
timestamp 1677622389
transform 1 0 1156 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8723
timestamp 1677622389
transform 1 0 1060 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8724
timestamp 1677622389
transform 1 0 1100 0 1 115
box -3 -3 3 3
use INVX2  INVX2_692
timestamp 1677622389
transform 1 0 1048 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_607
timestamp 1677622389
transform 1 0 1064 0 -1 170
box -8 -3 104 105
use FILL  FILL_10631
timestamp 1677622389
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use FILL  FILL_10632
timestamp 1677622389
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8636
timestamp 1677622389
transform 1 0 1244 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8637
timestamp 1677622389
transform 1 0 1268 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8647
timestamp 1677622389
transform 1 0 1188 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9912
timestamp 1677622389
transform 1 0 1188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9980
timestamp 1677622389
transform 1 0 1212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9981
timestamp 1677622389
transform 1 0 1268 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_608
timestamp 1677622389
transform 1 0 1176 0 -1 170
box -8 -3 104 105
use FILL  FILL_10633
timestamp 1677622389
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use FILL  FILL_10634
timestamp 1677622389
transform 1 0 1280 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8648
timestamp 1677622389
transform 1 0 1300 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9913
timestamp 1677622389
transform 1 0 1300 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9982
timestamp 1677622389
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9983
timestamp 1677622389
transform 1 0 1388 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_609
timestamp 1677622389
transform 1 0 1288 0 -1 170
box -8 -3 104 105
use FILL  FILL_10641
timestamp 1677622389
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8671
timestamp 1677622389
transform 1 0 1484 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9914
timestamp 1677622389
transform 1 0 1484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9984
timestamp 1677622389
transform 1 0 1404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9985
timestamp 1677622389
transform 1 0 1452 0 1 125
box -2 -2 2 2
use FILL  FILL_10655
timestamp 1677622389
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_610
timestamp 1677622389
transform -1 0 1496 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_9986
timestamp 1677622389
transform 1 0 1508 0 1 125
box -2 -2 2 2
use FILL  FILL_10656
timestamp 1677622389
transform 1 0 1496 0 -1 170
box -8 -3 16 105
use FILL  FILL_10657
timestamp 1677622389
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use FILL  FILL_10658
timestamp 1677622389
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8672
timestamp 1677622389
transform 1 0 1604 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9915
timestamp 1677622389
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9987
timestamp 1677622389
transform 1 0 1572 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_611
timestamp 1677622389
transform -1 0 1616 0 -1 170
box -8 -3 104 105
use FILL  FILL_10659
timestamp 1677622389
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8673
timestamp 1677622389
transform 1 0 1716 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9916
timestamp 1677622389
transform 1 0 1716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9917
timestamp 1677622389
transform 1 0 1732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9988
timestamp 1677622389
transform 1 0 1636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9989
timestamp 1677622389
transform 1 0 1692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9990
timestamp 1677622389
transform 1 0 1732 0 1 125
box -2 -2 2 2
use FILL  FILL_10667
timestamp 1677622389
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8725
timestamp 1677622389
transform 1 0 1692 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8726
timestamp 1677622389
transform 1 0 1732 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_612
timestamp 1677622389
transform -1 0 1728 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_697
timestamp 1677622389
transform 1 0 1728 0 -1 170
box -9 -3 26 105
use FILL  FILL_10668
timestamp 1677622389
transform 1 0 1744 0 -1 170
box -8 -3 16 105
use FILL  FILL_10669
timestamp 1677622389
transform 1 0 1752 0 -1 170
box -8 -3 16 105
use FILL  FILL_10671
timestamp 1677622389
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use FILL  FILL_10673
timestamp 1677622389
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8674
timestamp 1677622389
transform 1 0 1868 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9918
timestamp 1677622389
transform 1 0 1868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9919
timestamp 1677622389
transform 1 0 1884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9991
timestamp 1677622389
transform 1 0 1788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9992
timestamp 1677622389
transform 1 0 1844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9993
timestamp 1677622389
transform 1 0 1884 0 1 125
box -2 -2 2 2
use FILL  FILL_10683
timestamp 1677622389
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8727
timestamp 1677622389
transform 1 0 1844 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8728
timestamp 1677622389
transform 1 0 1884 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_613
timestamp 1677622389
transform -1 0 1880 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_699
timestamp 1677622389
transform 1 0 1880 0 -1 170
box -9 -3 26 105
use FILL  FILL_10684
timestamp 1677622389
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use FILL  FILL_10686
timestamp 1677622389
transform 1 0 1904 0 -1 170
box -8 -3 16 105
use FILL  FILL_10709
timestamp 1677622389
transform 1 0 1912 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8649
timestamp 1677622389
transform 1 0 1964 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8675
timestamp 1677622389
transform 1 0 2012 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9920
timestamp 1677622389
transform 1 0 2012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9994
timestamp 1677622389
transform 1 0 1932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9995
timestamp 1677622389
transform 1 0 1988 0 1 125
box -2 -2 2 2
use FILL  FILL_10710
timestamp 1677622389
transform 1 0 1920 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8751
timestamp 1677622389
transform 1 0 2028 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_618
timestamp 1677622389
transform -1 0 2024 0 -1 170
box -8 -3 104 105
use FILL  FILL_10711
timestamp 1677622389
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9996
timestamp 1677622389
transform 1 0 2044 0 1 125
box -2 -2 2 2
use FILL  FILL_10712
timestamp 1677622389
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_10713
timestamp 1677622389
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8676
timestamp 1677622389
transform 1 0 2132 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9921
timestamp 1677622389
transform 1 0 2132 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9997
timestamp 1677622389
transform 1 0 2108 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8745
timestamp 1677622389
transform 1 0 2092 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_8746
timestamp 1677622389
transform 1 0 2116 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_8752
timestamp 1677622389
transform 1 0 2092 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_619
timestamp 1677622389
transform -1 0 2144 0 -1 170
box -8 -3 104 105
use FILL  FILL_10714
timestamp 1677622389
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8650
timestamp 1677622389
transform 1 0 2164 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8677
timestamp 1677622389
transform 1 0 2228 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8678
timestamp 1677622389
transform 1 0 2244 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9922
timestamp 1677622389
transform 1 0 2244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9998
timestamp 1677622389
transform 1 0 2164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9999
timestamp 1677622389
transform 1 0 2220 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8710
timestamp 1677622389
transform 1 0 2244 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8747
timestamp 1677622389
transform 1 0 2164 0 1 95
box -3 -3 3 3
use FILL  FILL_10715
timestamp 1677622389
transform 1 0 2152 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_620
timestamp 1677622389
transform -1 0 2256 0 -1 170
box -8 -3 104 105
use FILL  FILL_10716
timestamp 1677622389
transform 1 0 2256 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8729
timestamp 1677622389
transform 1 0 2276 0 1 115
box -3 -3 3 3
use FILL  FILL_10717
timestamp 1677622389
transform 1 0 2264 0 -1 170
box -8 -3 16 105
use FILL  FILL_10718
timestamp 1677622389
transform 1 0 2272 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8679
timestamp 1677622389
transform 1 0 2292 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8680
timestamp 1677622389
transform 1 0 2324 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9923
timestamp 1677622389
transform 1 0 2292 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8711
timestamp 1677622389
transform 1 0 2292 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10000
timestamp 1677622389
transform 1 0 2316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10001
timestamp 1677622389
transform 1 0 2372 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8730
timestamp 1677622389
transform 1 0 2316 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_621
timestamp 1677622389
transform 1 0 2280 0 -1 170
box -8 -3 104 105
use FILL  FILL_10719
timestamp 1677622389
transform 1 0 2376 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8731
timestamp 1677622389
transform 1 0 2396 0 1 115
box -3 -3 3 3
use FILL  FILL_10720
timestamp 1677622389
transform 1 0 2384 0 -1 170
box -8 -3 16 105
use FILL  FILL_10721
timestamp 1677622389
transform 1 0 2392 0 -1 170
box -8 -3 16 105
use FILL  FILL_10722
timestamp 1677622389
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8748
timestamp 1677622389
transform 1 0 2420 0 1 95
box -3 -3 3 3
use FILL  FILL_10723
timestamp 1677622389
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_10724
timestamp 1677622389
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_10725
timestamp 1677622389
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_10726
timestamp 1677622389
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_10727
timestamp 1677622389
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_10728
timestamp 1677622389
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9924
timestamp 1677622389
transform 1 0 2468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10002
timestamp 1677622389
transform 1 0 2492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10003
timestamp 1677622389
transform 1 0 2516 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8732
timestamp 1677622389
transform 1 0 2516 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_622
timestamp 1677622389
transform 1 0 2456 0 -1 170
box -8 -3 104 105
use FILL  FILL_10729
timestamp 1677622389
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_10730
timestamp 1677622389
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8651
timestamp 1677622389
transform 1 0 2588 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8681
timestamp 1677622389
transform 1 0 2588 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9925
timestamp 1677622389
transform 1 0 2588 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10004
timestamp 1677622389
transform 1 0 2580 0 1 125
box -2 -2 2 2
use FILL  FILL_10731
timestamp 1677622389
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_10732
timestamp 1677622389
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_10734
timestamp 1677622389
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8652
timestamp 1677622389
transform 1 0 2620 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8682
timestamp 1677622389
transform 1 0 2612 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8683
timestamp 1677622389
transform 1 0 2636 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8684
timestamp 1677622389
transform 1 0 2700 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9926
timestamp 1677622389
transform 1 0 2700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10005
timestamp 1677622389
transform 1 0 2604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10006
timestamp 1677622389
transform 1 0 2612 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10007
timestamp 1677622389
transform 1 0 2652 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8733
timestamp 1677622389
transform 1 0 2604 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_10051
timestamp 1677622389
transform 1 0 2612 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_58
timestamp 1677622389
transform 1 0 2592 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_8734
timestamp 1677622389
transform 1 0 2652 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_623
timestamp 1677622389
transform -1 0 2712 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8685
timestamp 1677622389
transform 1 0 2724 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8686
timestamp 1677622389
transform 1 0 2772 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9927
timestamp 1677622389
transform 1 0 2724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10008
timestamp 1677622389
transform 1 0 2772 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_624
timestamp 1677622389
transform 1 0 2712 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8687
timestamp 1677622389
transform 1 0 2828 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9899
timestamp 1677622389
transform 1 0 2836 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_9928
timestamp 1677622389
transform 1 0 2828 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8703
timestamp 1677622389
transform 1 0 2836 0 1 135
box -3 -3 3 3
use INVX2  INVX2_706
timestamp 1677622389
transform 1 0 2808 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_10009
timestamp 1677622389
transform 1 0 2836 0 1 125
box -2 -2 2 2
use FILL  FILL_10742
timestamp 1677622389
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9929
timestamp 1677622389
transform 1 0 2852 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10010
timestamp 1677622389
transform 1 0 2860 0 1 125
box -2 -2 2 2
use NOR2X1  NOR2X1_121
timestamp 1677622389
transform 1 0 2832 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_8653
timestamp 1677622389
transform 1 0 2900 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8688
timestamp 1677622389
transform 1 0 2900 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8704
timestamp 1677622389
transform 1 0 2884 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9930
timestamp 1677622389
transform 1 0 2892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9931
timestamp 1677622389
transform 1 0 2900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9932
timestamp 1677622389
transform 1 0 2916 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8712
timestamp 1677622389
transform 1 0 2868 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10011
timestamp 1677622389
transform 1 0 2884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10052
timestamp 1677622389
transform 1 0 2868 0 1 115
box -2 -2 2 2
use FILL  FILL_10749
timestamp 1677622389
transform 1 0 2856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8735
timestamp 1677622389
transform 1 0 2876 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8705
timestamp 1677622389
transform 1 0 2924 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8654
timestamp 1677622389
transform 1 0 2956 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8689
timestamp 1677622389
transform 1 0 2940 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9933
timestamp 1677622389
transform 1 0 2932 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10012
timestamp 1677622389
transform 1 0 2908 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8713
timestamp 1677622389
transform 1 0 2916 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10013
timestamp 1677622389
transform 1 0 2924 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8743
timestamp 1677622389
transform 1 0 2892 0 1 105
box -3 -3 3 3
use OAI21X1  OAI21X1_186
timestamp 1677622389
transform -1 0 2896 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_10014
timestamp 1677622389
transform 1 0 2940 0 1 125
box -2 -2 2 2
use OAI22X1  OAI22X1_440
timestamp 1677622389
transform 1 0 2896 0 -1 170
box -8 -3 46 105
use FILL  FILL_10750
timestamp 1677622389
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10015
timestamp 1677622389
transform 1 0 2956 0 1 125
box -2 -2 2 2
use INVX2  INVX2_710
timestamp 1677622389
transform -1 0 2960 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_8638
timestamp 1677622389
transform 1 0 2996 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8690
timestamp 1677622389
transform 1 0 2972 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8691
timestamp 1677622389
transform 1 0 3004 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9934
timestamp 1677622389
transform 1 0 2972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9935
timestamp 1677622389
transform 1 0 2980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9936
timestamp 1677622389
transform 1 0 2996 0 1 135
box -2 -2 2 2
use FILL  FILL_10751
timestamp 1677622389
transform 1 0 2960 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10016
timestamp 1677622389
transform 1 0 2988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10017
timestamp 1677622389
transform 1 0 3004 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8736
timestamp 1677622389
transform 1 0 2988 0 1 115
box -3 -3 3 3
use AOI22X1  AOI22X1_418
timestamp 1677622389
transform 1 0 2968 0 -1 170
box -8 -3 46 105
use FILL  FILL_10753
timestamp 1677622389
transform 1 0 3008 0 -1 170
box -8 -3 16 105
use FILL  FILL_10755
timestamp 1677622389
transform 1 0 3016 0 -1 170
box -8 -3 16 105
use FILL  FILL_10785
timestamp 1677622389
transform 1 0 3024 0 -1 170
box -8 -3 16 105
use FILL  FILL_10786
timestamp 1677622389
transform 1 0 3032 0 -1 170
box -8 -3 16 105
use FILL  FILL_10787
timestamp 1677622389
transform 1 0 3040 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8706
timestamp 1677622389
transform 1 0 3084 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9937
timestamp 1677622389
transform 1 0 3132 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10018
timestamp 1677622389
transform 1 0 3084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10019
timestamp 1677622389
transform 1 0 3148 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8744
timestamp 1677622389
transform 1 0 3148 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_628
timestamp 1677622389
transform -1 0 3144 0 -1 170
box -8 -3 104 105
use FILL  FILL_10788
timestamp 1677622389
transform 1 0 3144 0 -1 170
box -8 -3 16 105
use FILL  FILL_10789
timestamp 1677622389
transform 1 0 3152 0 -1 170
box -8 -3 16 105
use FILL  FILL_10790
timestamp 1677622389
transform 1 0 3160 0 -1 170
box -8 -3 16 105
use FILL  FILL_10791
timestamp 1677622389
transform 1 0 3168 0 -1 170
box -8 -3 16 105
use FILL  FILL_10792
timestamp 1677622389
transform 1 0 3176 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_716
timestamp 1677622389
transform -1 0 3200 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_8692
timestamp 1677622389
transform 1 0 3284 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9938
timestamp 1677622389
transform 1 0 3284 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10020
timestamp 1677622389
transform 1 0 3260 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8737
timestamp 1677622389
transform 1 0 3260 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8639
timestamp 1677622389
transform 1 0 3300 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_10021
timestamp 1677622389
transform 1 0 3300 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_629
timestamp 1677622389
transform -1 0 3296 0 -1 170
box -8 -3 104 105
use FILL  FILL_10793
timestamp 1677622389
transform 1 0 3296 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8693
timestamp 1677622389
transform 1 0 3388 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9939
timestamp 1677622389
transform 1 0 3388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10022
timestamp 1677622389
transform 1 0 3364 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_630
timestamp 1677622389
transform -1 0 3400 0 -1 170
box -8 -3 104 105
use FILL  FILL_10794
timestamp 1677622389
transform 1 0 3400 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8694
timestamp 1677622389
transform 1 0 3420 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9940
timestamp 1677622389
transform 1 0 3420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10023
timestamp 1677622389
transform 1 0 3444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10024
timestamp 1677622389
transform 1 0 3500 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8738
timestamp 1677622389
transform 1 0 3444 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_631
timestamp 1677622389
transform 1 0 3408 0 -1 170
box -8 -3 104 105
use FILL  FILL_10795
timestamp 1677622389
transform 1 0 3504 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8695
timestamp 1677622389
transform 1 0 3572 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9941
timestamp 1677622389
transform 1 0 3524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10025
timestamp 1677622389
transform 1 0 3572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10026
timestamp 1677622389
transform 1 0 3604 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8749
timestamp 1677622389
transform 1 0 3604 0 1 95
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_632
timestamp 1677622389
transform 1 0 3512 0 -1 170
box -8 -3 104 105
use FILL  FILL_10796
timestamp 1677622389
transform 1 0 3608 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8640
timestamp 1677622389
transform 1 0 3652 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8696
timestamp 1677622389
transform 1 0 3644 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9942
timestamp 1677622389
transform 1 0 3628 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8714
timestamp 1677622389
transform 1 0 3628 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10027
timestamp 1677622389
transform 1 0 3676 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8750
timestamp 1677622389
transform 1 0 3644 0 1 95
box -3 -3 3 3
use M2_M1  M2_M1_10028
timestamp 1677622389
transform 1 0 3716 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_633
timestamp 1677622389
transform 1 0 3616 0 -1 170
box -8 -3 104 105
use FILL  FILL_10797
timestamp 1677622389
transform 1 0 3712 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9943
timestamp 1677622389
transform 1 0 3732 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8715
timestamp 1677622389
transform 1 0 3732 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10029
timestamp 1677622389
transform 1 0 3764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10030
timestamp 1677622389
transform 1 0 3820 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8739
timestamp 1677622389
transform 1 0 3820 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_634
timestamp 1677622389
transform 1 0 3720 0 -1 170
box -8 -3 104 105
use FILL  FILL_10798
timestamp 1677622389
transform 1 0 3816 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9944
timestamp 1677622389
transform 1 0 3836 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8716
timestamp 1677622389
transform 1 0 3836 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10031
timestamp 1677622389
transform 1 0 3860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10032
timestamp 1677622389
transform 1 0 3916 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8740
timestamp 1677622389
transform 1 0 3868 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_635
timestamp 1677622389
transform 1 0 3824 0 -1 170
box -8 -3 104 105
use FILL  FILL_10799
timestamp 1677622389
transform 1 0 3920 0 -1 170
box -8 -3 16 105
use FILL  FILL_10801
timestamp 1677622389
transform 1 0 3928 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9945
timestamp 1677622389
transform 1 0 3948 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8717
timestamp 1677622389
transform 1 0 3948 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10033
timestamp 1677622389
transform 1 0 3972 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8718
timestamp 1677622389
transform 1 0 4020 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10034
timestamp 1677622389
transform 1 0 4028 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_638
timestamp 1677622389
transform 1 0 3936 0 -1 170
box -8 -3 104 105
use FILL  FILL_10809
timestamp 1677622389
transform 1 0 4032 0 -1 170
box -8 -3 16 105
use FILL  FILL_10810
timestamp 1677622389
transform 1 0 4040 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9946
timestamp 1677622389
transform 1 0 4060 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8719
timestamp 1677622389
transform 1 0 4060 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10035
timestamp 1677622389
transform 1 0 4092 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10036
timestamp 1677622389
transform 1 0 4140 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8753
timestamp 1677622389
transform 1 0 4116 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_8754
timestamp 1677622389
transform 1 0 4140 0 1 75
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_639
timestamp 1677622389
transform 1 0 4048 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8655
timestamp 1677622389
transform 1 0 4156 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8656
timestamp 1677622389
transform 1 0 4188 0 1 155
box -3 -3 3 3
use FILL  FILL_10811
timestamp 1677622389
transform 1 0 4144 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9947
timestamp 1677622389
transform 1 0 4164 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8720
timestamp 1677622389
transform 1 0 4164 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10037
timestamp 1677622389
transform 1 0 4188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10038
timestamp 1677622389
transform 1 0 4244 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_640
timestamp 1677622389
transform 1 0 4152 0 -1 170
box -8 -3 104 105
use FILL  FILL_10812
timestamp 1677622389
transform 1 0 4248 0 -1 170
box -8 -3 16 105
use FILL  FILL_10813
timestamp 1677622389
transform 1 0 4256 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9948
timestamp 1677622389
transform 1 0 4276 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8721
timestamp 1677622389
transform 1 0 4276 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10039
timestamp 1677622389
transform 1 0 4308 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10040
timestamp 1677622389
transform 1 0 4356 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_641
timestamp 1677622389
transform 1 0 4264 0 -1 170
box -8 -3 104 105
use FILL  FILL_10814
timestamp 1677622389
transform 1 0 4360 0 -1 170
box -8 -3 16 105
use FILL  FILL_10816
timestamp 1677622389
transform 1 0 4368 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9949
timestamp 1677622389
transform 1 0 4388 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8722
timestamp 1677622389
transform 1 0 4388 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10041
timestamp 1677622389
transform 1 0 4420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10042
timestamp 1677622389
transform 1 0 4468 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_644
timestamp 1677622389
transform 1 0 4376 0 -1 170
box -8 -3 104 105
use FILL  FILL_10826
timestamp 1677622389
transform 1 0 4472 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8657
timestamp 1677622389
transform 1 0 4580 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8697
timestamp 1677622389
transform 1 0 4540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8698
timestamp 1677622389
transform 1 0 4572 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9950
timestamp 1677622389
transform 1 0 4492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9951
timestamp 1677622389
transform 1 0 4588 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9952
timestamp 1677622389
transform 1 0 4596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10043
timestamp 1677622389
transform 1 0 4540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10044
timestamp 1677622389
transform 1 0 4572 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_645
timestamp 1677622389
transform 1 0 4480 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_723
timestamp 1677622389
transform -1 0 4592 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_8658
timestamp 1677622389
transform 1 0 4604 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10045
timestamp 1677622389
transform 1 0 4604 0 1 125
box -2 -2 2 2
use FILL  FILL_10827
timestamp 1677622389
transform 1 0 4592 0 -1 170
box -8 -3 16 105
use FILL  FILL_10828
timestamp 1677622389
transform 1 0 4600 0 -1 170
box -8 -3 16 105
use FILL  FILL_10829
timestamp 1677622389
transform 1 0 4608 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8641
timestamp 1677622389
transform 1 0 4636 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8699
timestamp 1677622389
transform 1 0 4644 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9953
timestamp 1677622389
transform 1 0 4628 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9954
timestamp 1677622389
transform 1 0 4644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9955
timestamp 1677622389
transform 1 0 4660 0 1 135
box -2 -2 2 2
use FILL  FILL_10830
timestamp 1677622389
transform 1 0 4616 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10046
timestamp 1677622389
transform 1 0 4636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10047
timestamp 1677622389
transform 1 0 4652 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8741
timestamp 1677622389
transform 1 0 4652 0 1 115
box -3 -3 3 3
use OAI22X1  OAI22X1_451
timestamp 1677622389
transform -1 0 4664 0 -1 170
box -8 -3 46 105
use FILL  FILL_10831
timestamp 1677622389
transform 1 0 4664 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8642
timestamp 1677622389
transform 1 0 4724 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8700
timestamp 1677622389
transform 1 0 4708 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9956
timestamp 1677622389
transform 1 0 4684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9957
timestamp 1677622389
transform 1 0 4780 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10048
timestamp 1677622389
transform 1 0 4708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10049
timestamp 1677622389
transform 1 0 4764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10050
timestamp 1677622389
transform 1 0 4772 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8742
timestamp 1677622389
transform 1 0 4772 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_646
timestamp 1677622389
transform 1 0 4672 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_724
timestamp 1677622389
transform -1 0 4784 0 -1 170
box -9 -3 26 105
use FILL  FILL_10832
timestamp 1677622389
transform 1 0 4784 0 -1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_93
timestamp 1677622389
transform 1 0 4843 0 1 70
box -10 -3 10 3
use M3_M2  M3_M2_8755
timestamp 1677622389
transform 1 0 3716 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_8756
timestamp 1677622389
transform 1 0 3748 0 1 65
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_4
timestamp 1677622389
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_6
timestamp 1677622389
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_8757
timestamp 1677622389
transform 1 0 2172 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_8758
timestamp 1677622389
transform 1 0 2228 0 1 35
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_5
timestamp 1677622389
transform 1 0 4819 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_8759
timestamp 1677622389
transform 1 0 2468 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8760
timestamp 1677622389
transform 1 0 2724 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8761
timestamp 1677622389
transform 1 0 3892 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8762
timestamp 1677622389
transform 1 0 3916 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8763
timestamp 1677622389
transform 1 0 3964 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8764
timestamp 1677622389
transform 1 0 4028 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8765
timestamp 1677622389
transform 1 0 4068 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8766
timestamp 1677622389
transform 1 0 4100 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8767
timestamp 1677622389
transform 1 0 4212 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8768
timestamp 1677622389
transform 1 0 4244 0 1 15
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_7
timestamp 1677622389
transform 1 0 4843 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal2 2724 1 2724 1 4 clka
rlabel metal3 2 2075 2 2075 4 clkb
rlabel metal2 2492 1 2492 1 4 reset
rlabel metal2 2516 1 2516 1 4 we_ins
rlabel metal2 2116 1 2116 1 4 load[15]
rlabel metal2 2132 1 2132 1 4 load[14]
rlabel metal2 2156 1 2156 1 4 load[13]
rlabel metal2 2364 1 2364 1 4 load[12]
rlabel metal2 2092 1 2092 1 4 load[11]
rlabel metal2 2172 1 2172 1 4 load[10]
rlabel metal2 2196 1 2196 1 4 load[9]
rlabel metal2 2212 1 2212 1 4 load[8]
rlabel metal2 2332 1 2332 1 4 load[7]
rlabel metal2 2276 1 2276 1 4 load[6]
rlabel metal2 2316 1 2316 1 4 load[5]
rlabel metal2 2348 1 2348 1 4 load[4]
rlabel metal2 2228 1 2228 1 4 load[3]
rlabel metal2 2244 1 2244 1 4 load[2]
rlabel metal2 2260 1 2260 1 4 load[1]
rlabel metal2 2076 1 2076 1 4 load[0]
rlabel metal2 4212 1 4212 1 4 reg_0_out[7]
rlabel metal2 3868 1 3868 1 4 reg_0_out[6]
rlabel metal2 4068 1 4068 1 4 reg_0_out[5]
rlabel metal2 3892 1 3892 1 4 reg_0_out[4]
rlabel metal2 3748 1 3748 1 4 reg_0_out[3]
rlabel metal2 3644 1 3644 1 4 reg_0_out[2]
rlabel metal2 4116 1 4116 1 4 reg_0_out[1]
rlabel metal2 3964 1 3964 1 4 reg_0_out[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>

magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 104 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 16
rect 21 6 23 16
rect 29 6 31 16
rect 34 6 36 16
rect 43 6 45 16
rect 59 6 61 16
rect 64 6 66 16
rect 74 6 76 16
rect 79 6 81 16
rect 87 6 89 26
<< ptransistor >>
rect 7 54 9 94
rect 15 74 17 94
rect 21 74 23 94
rect 29 74 31 94
rect 35 74 37 94
rect 43 74 45 94
rect 59 74 61 94
rect 64 74 66 94
rect 74 84 76 94
rect 79 84 81 94
rect 87 54 89 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 16 14 26
rect 82 16 87 26
rect 9 6 15 16
rect 17 6 21 16
rect 23 6 29 16
rect 31 6 34 16
rect 36 6 43 16
rect 45 6 50 16
rect 54 6 59 16
rect 61 6 64 16
rect 66 6 74 16
rect 76 6 79 16
rect 81 6 87 16
rect 89 6 94 26
<< pdiffusion >>
rect 2 54 7 94
rect 9 74 15 94
rect 17 74 21 94
rect 23 74 29 94
rect 31 74 35 94
rect 37 74 43 94
rect 45 74 50 94
rect 54 74 59 94
rect 61 74 64 94
rect 66 84 74 94
rect 76 84 79 94
rect 81 84 87 94
rect 66 74 73 84
rect 9 54 14 74
rect 82 54 87 84
rect 89 54 94 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 21 94 23 96
rect 29 94 31 96
rect 35 94 37 96
rect 43 94 45 96
rect 59 94 61 96
rect 64 94 66 96
rect 74 94 76 96
rect 79 94 81 96
rect 87 94 89 96
rect 7 37 9 54
rect 15 46 17 74
rect 21 54 23 74
rect 29 71 31 74
rect 27 67 31 71
rect 35 71 37 74
rect 35 67 39 71
rect 21 52 25 54
rect 21 50 31 52
rect 14 42 18 46
rect 6 33 10 37
rect 7 26 9 33
rect 15 16 17 42
rect 21 23 25 27
rect 21 16 23 23
rect 29 16 31 50
rect 35 23 37 67
rect 43 61 45 74
rect 59 73 61 74
rect 50 71 61 73
rect 41 57 45 61
rect 34 19 39 23
rect 34 16 36 19
rect 43 16 45 57
rect 49 67 53 71
rect 64 67 66 74
rect 49 19 51 67
rect 63 65 66 67
rect 55 60 59 61
rect 54 57 59 60
rect 54 24 56 57
rect 63 37 65 65
rect 74 61 76 84
rect 69 57 76 61
rect 79 53 81 84
rect 75 51 81 53
rect 73 47 77 51
rect 60 33 65 37
rect 60 29 62 33
rect 74 31 76 47
rect 87 45 89 54
rect 81 41 89 45
rect 60 27 71 29
rect 74 27 81 31
rect 54 22 66 24
rect 49 17 61 19
rect 59 16 61 17
rect 64 16 66 22
rect 69 19 71 27
rect 69 17 76 19
rect 74 16 76 17
rect 79 16 81 27
rect 87 26 89 41
rect 7 4 9 6
rect 15 4 17 6
rect 21 4 23 6
rect 29 4 31 6
rect 34 4 36 6
rect 43 4 45 6
rect 59 4 61 6
rect 64 4 66 6
rect 74 4 76 6
rect 79 4 81 6
rect 87 4 89 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 31 99 33 101
rect 47 99 49 101
rect 63 99 65 101
rect 79 99 81 101
rect 3 90 5 92
rect 11 91 13 93
rect 25 90 27 92
rect 39 90 41 92
rect 47 90 49 92
rect 55 90 57 92
rect 69 90 71 92
rect 83 90 85 92
rect 91 90 93 92
rect 3 85 5 87
rect 11 86 13 88
rect 25 85 27 87
rect 39 85 41 87
rect 47 85 49 87
rect 55 85 57 87
rect 69 85 71 87
rect 83 85 85 87
rect 91 85 93 87
rect 3 80 5 82
rect 11 81 13 83
rect 25 80 27 82
rect 39 80 41 82
rect 47 80 49 82
rect 55 80 57 82
rect 69 80 71 82
rect 83 80 85 82
rect 91 80 93 82
rect 3 75 5 77
rect 11 76 13 78
rect 25 75 27 77
rect 39 75 41 77
rect 47 75 49 77
rect 55 75 57 77
rect 69 75 71 77
rect 83 75 85 77
rect 91 75 93 77
rect 3 70 5 72
rect 11 71 13 73
rect 83 70 85 72
rect 91 70 93 72
rect 28 68 30 70
rect 36 68 38 70
rect 50 68 52 70
rect 3 65 5 67
rect 11 66 13 68
rect 83 65 85 67
rect 91 65 93 67
rect 3 60 5 62
rect 11 61 13 63
rect 83 60 85 62
rect 91 60 93 62
rect 42 58 44 60
rect 56 58 58 60
rect 70 58 72 60
rect 3 55 5 57
rect 11 56 13 58
rect 83 55 85 57
rect 91 55 93 57
rect 22 51 24 53
rect 74 48 76 50
rect 15 43 17 45
rect 82 42 84 44
rect 7 34 9 36
rect 61 34 63 36
rect 76 28 78 30
rect 22 24 24 26
rect 3 22 5 24
rect 11 22 13 24
rect 83 22 85 24
rect 91 22 93 24
rect 36 20 38 22
rect 3 17 5 19
rect 11 17 13 19
rect 83 17 85 19
rect 91 17 93 19
rect 3 12 5 14
rect 11 12 13 14
rect 25 12 27 14
rect 38 12 40 14
rect 47 12 49 14
rect 55 12 57 14
rect 69 12 71 14
rect 83 12 85 14
rect 91 12 93 14
rect 3 7 5 9
rect 11 7 13 9
rect 25 7 27 9
rect 38 7 40 9
rect 47 7 49 9
rect 55 7 57 9
rect 69 7 71 9
rect 83 7 85 9
rect 91 7 93 9
rect -1 -1 1 1
rect 15 -1 17 1
rect 31 -1 33 1
rect 47 -1 49 1
rect 63 -1 65 1
rect 79 -1 81 1
<< metal1 >>
rect -2 97 98 103
rect 2 52 6 94
rect 10 55 14 97
rect 24 77 28 94
rect 18 74 28 77
rect 38 74 42 97
rect 46 74 50 94
rect 54 74 58 97
rect 67 74 73 94
rect 18 70 22 74
rect 46 71 49 74
rect 27 67 31 71
rect 35 68 53 71
rect 66 70 70 74
rect 35 67 39 68
rect 49 67 53 68
rect 26 63 30 67
rect 18 60 22 61
rect 41 60 45 61
rect 18 57 45 60
rect 54 60 59 61
rect 69 60 73 61
rect 54 57 73 60
rect 54 54 57 57
rect 82 54 86 97
rect 21 52 57 54
rect 2 51 57 52
rect 90 51 94 94
rect 2 49 25 51
rect 73 48 94 51
rect 73 47 77 48
rect 34 46 38 47
rect 14 43 38 46
rect 81 44 85 45
rect 14 42 18 43
rect 66 41 85 44
rect 66 40 70 41
rect 26 37 30 38
rect 6 34 64 37
rect 6 33 14 34
rect 2 6 6 30
rect 20 27 24 34
rect 60 33 64 34
rect 90 31 94 48
rect 75 28 94 31
rect 75 27 79 28
rect 10 3 14 26
rect 21 23 25 27
rect 35 22 39 23
rect 18 16 22 20
rect 35 19 49 22
rect 46 16 49 19
rect 66 16 70 20
rect 18 13 28 16
rect 24 6 28 13
rect 37 3 42 16
rect 46 6 50 16
rect 54 3 58 16
rect 66 13 73 16
rect 67 6 73 13
rect 82 3 86 25
rect 90 6 94 28
rect -2 -3 98 3
<< metal2 >>
rect 18 54 22 74
rect 2 26 6 54
rect 18 50 21 54
rect 18 16 22 50
rect 26 34 30 67
rect 66 61 70 74
rect 66 57 69 61
rect 66 16 70 57
<< gv1 >>
rect 19 71 21 73
rect 67 71 69 73
rect 27 64 29 66
rect 19 58 21 60
rect 3 51 5 53
rect 67 41 69 43
rect 27 35 29 37
rect 3 27 5 29
rect 19 17 21 19
rect 67 17 69 19
<< m1p >>
rect 34 43 38 47
rect 90 43 94 47
rect 10 33 14 37
<< labels >>
rlabel metal1 12 35 12 35 6 CLK
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 36 45 36 45 6 D
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 92 45 92 45 6 Q
<< end >>

`timescale 1ns/100ps
module alu_fsm_tb();

reg     in_clka,
        in_clkb,
        reset_in,
        n_dec_in,
        z_dec_in,
        p_dec_in,
        n_alu_in,
        z_alu_in,
        p_alu_in,
        we_reg_in,
        br_in;

wire [3:0] state_out;
wire pc_ctl_0_out;
wire pc_latch_clkedge;

//create an FSM instance.
ALU_FSM fsm (
        .clka (in_clka),
        .clkb (in_clkb),
        .reset_in (reset_in),
        .n_dec_in (n_dec_in),
        .z_dec_in (z_dec_in),
        .p_dec_in (p_dec_in),
        .n_alu_in (n_alu_in),
        .z_alu_in (z_alu_in),
        .p_alu_in (p_alu_in),
        .we_reg_in (we_reg_in),
        .br_in (br_in),
        .pc_ctl_0_out (pc_ctl_0_out),
        .pc_latch_clkedge(pc_latch_clkedge)
        .state_out (state_out)
);

initial begin

reset_in = 0;
n_dec_in = 0;
z_dec_in = 0;
p_dec_in = 0;
n_alu_in = 0;
z_alu_in = 0;
p_alu_in = 0;
we_reg_in = 0;
br_in = 0;
in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

reset_in = 1; //reset fsm - turns to a PC Cycle

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// do for two cycles to verify that reset always holds in a PC Cycle

reset_in = 0; // the PC should latch on this clka, output on clkb

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
 // PC Output here

/**
The following blocks test that the state is not updated when the we signal is 
not asserted 
**/ 

n_alu_in = 1; // PC Should be static this cycle, FSM Should latch update here

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM Output Here


in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC Output here

n_alu_in = 0;
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM Output HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
//PC Output Here

z_alu_in = 0;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
//FSM Output HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC Output HERE

p_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM Output HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC Output HERE

/**
The following tests verify that the FSM moves between states properly
**/
we_reg_in = 1;
n_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
//FSM OUTPUT HERE

n_alu_in = 0;
we_reg_in = 0; // make sure alu not latched on wrong clk

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
n_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

n_alu_in = 0;
we_reg_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

we_reg_in = 0;
z_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

z_alu_in = 0;
we_reg_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

we_reg_in = 0;
p_alu_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

p_alu_in = 1;
we_reg_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

p_alu_in = 0;
we_reg_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

/**
The following test check that the ALU Properly asserts the 
branch out bit when it should
**/

reset_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

reset_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
n_alu_in = 1; //set state to n

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 0;
n_alu_in = 0;
n_dec_in = 1;
br_in = 1; //should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
z_alu_in = 1;
n_dec_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 0;
z_alu_in = 0;
z_dec_in = 1;
br_in = 1; // should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 1;
p_alu_in = 1;
z_dec_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

we_reg_in = 0;
p_alu_in = 0;
p_dec_in = 1;
br_in = 1; //should cause branch

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE


/**
The following tests verify that the FSM does not assert branch at the wrong time
**/

//cases when br is not asserted
we_reg_in = 1;
n_dec_in = 1;
n_alu_in = 1;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

p_dec_in = 1;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

z_dec_in = 1; // branch should not be asserted here
z_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
//FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE

//cases when wrong dec asserted
we_reg_in = 1;
br_in = 1;
n_alu_in = 1;
p_dec_in = 1;
z_dec_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM OUTPUT HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC OUTPUT HERE


n_alu_in = 0;
p_dec_in = 0;
n_dec_in = 1;
p_alu_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE
in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

p_alu_in = 0;
p_dec_in = 1;
z_alu_in = 1;
z_dec_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE
in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

//clear all signals
reset_in = 0;
n_dec_in = 0;
z_dec_in = 0;
p_dec_in = 0;
n_alu_in = 0;
z_alu_in = 0;
p_alu_in = 0;
we_reg_in = 0;
br_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

//assert reset

reset_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE

reset_in = 0;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

//verify no branches taken in idle

br_in = 1;
n_dec_in = 1;
p_dec_in = 1;
z_dec_in = 1;

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// FSM HERE

in_clka = 0; in_clkb = 0; #10;
in_clka = 1; in_clkb = 0; #10;
in_clka = 0; in_clkb = 0; #10;
in_clka = 0; in_clkb = 1; #10;
// PC HERE


end

endmodule
magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 34 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
rect 20 74 22 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 15 26
rect 17 6 23 26
rect 25 6 30 26
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 12 94
rect 14 74 20 94
rect 22 74 27 94
rect 14 54 19 74
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 20 94 22 96
rect 20 67 22 74
rect 20 65 26 67
rect 22 63 26 65
rect 7 49 9 54
rect 12 53 14 54
rect 12 51 17 53
rect 4 47 9 49
rect 4 35 6 47
rect 15 43 17 51
rect 10 39 17 43
rect 4 33 10 35
rect 6 31 10 33
rect 7 26 9 31
rect 15 26 17 39
rect 23 26 25 63
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 16 90 18 92
rect 24 90 26 92
rect 3 85 5 87
rect 16 85 18 87
rect 24 85 26 87
rect 3 80 5 82
rect 16 80 18 82
rect 24 80 26 82
rect 3 75 5 77
rect 16 75 18 77
rect 24 75 26 77
rect 3 70 5 72
rect 16 70 18 72
rect 3 65 5 67
rect 16 65 18 67
rect 23 64 25 66
rect 3 60 5 62
rect 16 60 18 62
rect 3 55 5 57
rect 16 55 18 57
rect 11 40 13 42
rect 7 32 9 34
rect 3 22 5 24
rect 19 22 21 24
rect 27 22 29 24
rect 3 17 5 19
rect 11 18 13 20
rect 19 17 21 19
rect 27 17 29 19
rect 3 12 5 14
rect 11 13 13 15
rect 19 12 21 14
rect 27 12 29 14
rect 3 7 5 9
rect 11 8 13 10
rect 19 7 21 9
rect 27 7 29 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 34 103
rect 2 54 6 97
rect 15 57 19 94
rect 23 74 27 97
rect 22 63 26 67
rect 23 57 26 63
rect 15 54 20 57
rect 23 54 30 57
rect 10 39 14 47
rect 17 37 20 54
rect 26 53 30 54
rect 2 36 6 37
rect 2 33 10 36
rect 17 33 30 37
rect 6 31 10 33
rect 3 26 21 28
rect 26 26 29 33
rect 2 25 22 26
rect 2 6 6 25
rect 10 3 14 22
rect 18 6 22 25
rect 26 6 30 26
rect -2 -3 34 3
<< m1p >>
rect 26 53 30 57
rect 10 43 14 47
rect 2 33 6 37
rect 26 33 30 37
<< labels >>
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 35 4 35 6 A
rlabel metal1 12 45 12 45 6 B
rlabel metal1 28 35 28 35 6 Y
rlabel metal1 28 55 28 55 6 C
<< end >>

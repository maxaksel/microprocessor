magic
tech scmos
timestamp 1682046639
<< metal1 >>
rect -1368 4094 -1336 4124
rect -1064 4091 -1026 4122
rect -768 4093 -734 4123
rect -468 4097 -431 4123
rect -173 4089 -116 4133
rect 128 4093 180 4132
rect 422 4091 473 4124
rect 731 4090 780 4127
rect 1034 4095 1080 4129
rect 1329 4097 1378 4128
rect 1638 4094 1679 4129
rect 1925 4098 1982 4132
rect 1931 4096 1972 4098
rect 2227 4097 2273 4132
rect 2525 4095 2583 4127
rect 2838 4101 2869 4125
rect 3130 4093 3181 4131
rect -1481 3357 -1398 3366
rect -2223 3227 -2201 3273
rect -1414 3135 -1398 3357
rect -1243 3151 -1234 3381
rect -943 3168 -934 3381
rect -643 3184 -634 3381
rect -343 3199 -334 3381
rect -43 3214 -34 3381
rect 257 3229 266 3381
rect 402 3379 498 3391
rect 857 3372 866 3381
rect 747 3362 866 3372
rect 257 3218 730 3229
rect -43 3203 714 3214
rect -343 3188 698 3199
rect -643 3173 682 3184
rect -943 3157 658 3168
rect -1243 3140 642 3151
rect -1414 3124 621 3135
rect 637 3128 642 3140
rect 653 3128 658 3157
rect 677 3128 682 3173
rect 693 3128 698 3188
rect 709 3128 714 3203
rect 725 3128 730 3218
rect 747 2932 756 3362
rect 1157 3358 1166 3381
rect 763 3347 1166 3358
rect 763 2932 772 3347
rect 1457 3337 1466 3381
rect 779 3329 1466 3337
rect 779 2932 788 3329
rect 1757 3317 1766 3377
rect 795 3309 1766 3317
rect 795 2932 804 3309
rect 2057 3301 2066 3376
rect 811 3293 2068 3301
rect 811 2932 820 3293
rect 2357 3286 2366 3375
rect 827 3275 2366 3286
rect 2502 3379 2598 3392
rect 827 2932 836 3275
rect 2957 3268 2966 3376
rect 3257 3375 3266 3376
rect 843 3259 2966 3268
rect 3178 3367 3266 3375
rect 843 2932 852 3259
rect 3178 3254 3187 3367
rect 859 3246 3187 3254
rect 3204 3349 3290 3357
rect 859 2932 868 3246
rect 3204 3241 3213 3349
rect 875 3233 3213 3241
rect 875 2932 884 3233
rect 3993 3231 4023 3271
rect 891 3218 3262 3226
rect 891 2931 900 3218
rect 1461 3206 3228 3213
rect 1461 2928 1466 3206
rect 1517 3194 3207 3201
rect 1517 2928 1522 3194
rect 1533 3182 3191 3189
rect 1533 2928 1538 3182
rect 1597 3172 3158 3179
rect 1597 2928 1602 3172
rect 1725 3162 3146 3169
rect 1725 2928 1730 3162
rect 1893 3151 3134 3158
rect 1893 2928 1898 3151
rect 2085 3140 3122 3147
rect 2085 2928 2090 3140
rect 3014 2149 3110 2156
rect 3014 2119 3098 2126
rect 3014 2099 3087 2106
rect -2224 2022 -2190 2076
rect -1481 1257 -1228 1266
rect -2225 1132 -2200 1171
rect -1235 1109 -1228 1257
rect -2218 233 -2192 265
rect 3080 -747 3087 2099
rect 3091 -447 3098 2119
rect 3103 153 3110 2149
rect 3115 453 3122 3140
rect 3127 753 3134 3151
rect 3139 1053 3146 3162
rect 3151 1353 3158 3172
rect 3184 2166 3191 3182
rect 3200 2466 3207 3194
rect 3221 2553 3228 3206
rect 3254 3066 3262 3218
rect 3254 3057 3281 3066
rect 3990 2929 4022 2979
rect 3992 2631 4025 2673
rect 3221 2544 3265 2553
rect 3200 2457 3261 2466
rect 3995 2316 4024 2367
rect 3184 2157 3264 2166
rect 4001 2020 4024 2076
rect 3989 1784 4021 1785
rect 3989 1724 4022 1784
rect 3993 1722 4022 1724
rect 3995 1428 4028 1476
rect 3151 1344 3265 1353
rect 3995 1123 4028 1180
rect 3139 1044 3265 1053
rect 3992 820 4022 876
rect 3127 744 3265 753
rect 3995 521 4026 576
rect 3115 444 3264 453
rect 3985 233 4026 272
rect 3103 144 3265 153
rect 3987 -70 4024 -20
rect 3995 -376 4026 -319
rect 3091 -456 3265 -447
rect 3995 -676 4029 -614
rect 3080 -756 3265 -747
<< m2contact >>
rect -1389 3388 -1380 3392
rect -1243 3381 -1234 3389
rect -1089 3388 -1085 3392
rect -1489 3357 -1481 3366
rect -1492 3211 -1488 3215
rect -943 3381 -934 3390
rect -789 3388 -785 3392
rect -643 3381 -634 3390
rect -489 3388 -485 3392
rect -343 3381 -334 3390
rect -189 3388 -185 3393
rect -43 3381 -34 3390
rect 111 3388 115 3392
rect 257 3381 266 3390
rect 711 3388 715 3392
rect 402 3277 498 3379
rect 857 3381 866 3389
rect 1011 3388 1015 3392
rect 1157 3381 1166 3389
rect 1311 3388 1315 3392
rect -621 2895 -372 2993
rect 621 2921 626 3135
rect 637 2921 642 3128
rect 653 2921 658 3128
rect 677 2921 682 3128
rect 693 2921 698 3128
rect 709 2921 714 3128
rect 725 2921 730 3128
rect 747 2920 756 2932
rect 1457 3381 1466 3390
rect 1611 3388 1615 3392
rect 1911 3388 1915 3392
rect 2211 3388 2215 3392
rect 763 2920 772 2932
rect 1757 3377 1766 3386
rect 779 2920 788 2932
rect 2057 3376 2066 3386
rect 2357 3375 2366 3385
rect 795 2920 804 2932
rect 811 2920 820 2932
rect 2811 3388 2815 3392
rect 3111 3388 3115 3392
rect 2502 3276 2598 3379
rect 2957 3376 2966 3385
rect 3257 3376 3266 3384
rect 827 2920 836 2932
rect 3281 3357 3290 3366
rect 843 2920 852 2932
rect 859 2920 868 2932
rect 875 2920 884 2932
rect 891 2920 900 2931
rect 1461 2924 1466 2928
rect 1517 2924 1522 2928
rect 1533 2924 1538 2928
rect 1597 2924 1602 2928
rect 1725 2924 1730 2928
rect 1893 2924 1898 2928
rect 2085 2924 2090 2928
rect 2619 2895 2889 2982
rect 3007 2149 3014 2156
rect 3007 2119 3014 2126
rect 3007 2099 3014 2106
rect -1489 2002 -1478 2098
rect -1489 1257 -1481 1266
rect -1492 1111 -1488 1115
rect -1228 1109 -1221 1116
rect -1489 202 -1480 298
rect 3288 3211 3292 3215
rect 3281 3057 3290 3066
rect 3288 2911 3292 2915
rect 3288 2611 3292 2615
rect 3265 2544 3284 2553
rect 3261 2457 3285 2466
rect 3288 2311 3292 2315
rect 3264 2157 3282 2166
rect 3288 2011 3292 2015
rect 3276 1702 3289 1798
rect 3288 1411 3292 1415
rect 3265 1344 3282 1353
rect 3288 1111 3292 1115
rect 3265 1044 3283 1053
rect 3288 811 3292 815
rect 3265 744 3282 753
rect 3288 511 3292 515
rect 3264 444 3282 453
rect 3288 211 3292 215
rect 3265 144 3282 153
rect 3283 -98 3289 -2
rect 3288 -389 3292 -385
rect 3265 -456 3283 -447
rect 3288 -689 3292 -685
rect 3265 -756 3282 -747
rect -198 -1390 -102 -1367
rect 1602 -1390 1698 -1374
<< metal2 >>
rect -1389 3344 -1380 3388
rect -1089 3379 -1085 3388
rect -1092 3344 -1082 3379
rect -789 3379 -785 3388
rect -792 3344 -783 3379
rect -489 3379 -485 3388
rect 111 3392 115 3393
rect -491 3344 -483 3379
rect -189 3379 -185 3388
rect -191 3344 -183 3379
rect 111 3379 115 3388
rect 109 3344 117 3379
rect -1460 3277 402 3344
rect 711 3344 715 3388
rect 1011 3344 1015 3388
rect 1311 3344 1315 3388
rect 1595 3382 1599 3388
rect 1611 3344 1615 3388
rect 1911 3344 1915 3388
rect 2211 3344 2215 3388
rect 498 3277 2502 3344
rect -1460 3215 -1399 3277
rect -1488 3211 -1399 3215
rect -1460 1115 -1399 3211
rect -620 2993 -373 3277
rect 2811 3344 2815 3388
rect 3111 3344 3115 3388
rect 3290 3357 3297 3366
rect 3281 3344 3297 3353
rect 2598 3277 3250 3344
rect 2619 2982 2888 3277
rect 3180 3215 3250 3277
rect 3180 3211 3288 3215
rect 3180 2915 3250 3211
rect 3180 2911 3288 2915
rect 3180 2615 3250 2911
rect 3180 2611 3288 2615
rect 3180 2529 3250 2611
rect 3180 2523 3283 2529
rect 3180 2315 3250 2523
rect 3180 2311 3288 2315
rect 3000 2155 3007 2156
rect 3000 2150 3001 2155
rect 3006 2150 3007 2155
rect 3000 2149 3007 2150
rect 3000 2125 3007 2126
rect 3000 2120 3001 2125
rect 3006 2120 3007 2125
rect 3000 2119 3007 2120
rect 3000 2105 3007 2106
rect 3000 2100 3001 2105
rect 3006 2100 3007 2105
rect 3000 2099 3007 2100
rect 3180 2015 3250 2311
rect 3180 2011 3288 2015
rect 3180 1415 3250 2011
rect 3180 1411 3288 1415
rect 3180 1329 3250 1411
rect 3180 1323 3283 1329
rect -1488 1111 -1399 1115
rect -1460 -1305 -1399 1111
rect -1221 1115 -1214 1116
rect -1221 1110 -1220 1115
rect -1215 1110 -1214 1115
rect -1221 1109 -1214 1110
rect 3180 1115 3250 1323
rect 3180 1111 3288 1115
rect 3180 1029 3250 1111
rect 3180 1023 3283 1029
rect 3180 815 3250 1023
rect 3180 811 3288 815
rect 3180 729 3250 811
rect 3180 723 3283 729
rect 3180 515 3250 723
rect 3180 511 3288 515
rect 3180 429 3250 511
rect 3180 423 3284 429
rect 3180 215 3250 423
rect 3180 211 3288 215
rect 3180 129 3250 211
rect 3180 123 3286 129
rect 3180 -385 3250 123
rect 3180 -389 3288 -385
rect 3180 -471 3250 -389
rect 3180 -477 3286 -471
rect 3180 -685 3250 -477
rect 3180 -689 3288 -685
rect 3180 -771 3250 -689
rect 3180 -777 3283 -771
rect 3180 -1271 3250 -777
rect 3179 -1305 3250 -1271
rect -1460 -1345 3250 -1305
rect -1461 -1356 3250 -1345
rect -198 -1367 -102 -1356
rect 1602 -1374 1698 -1356
<< m3contact >>
rect -1405 3388 -1401 3392
rect -1477 3378 -1471 3384
rect -1105 3388 -1101 3392
rect -1177 3378 -1171 3383
rect -805 3388 -801 3392
rect -877 3377 -871 3383
rect -505 3387 -501 3392
rect -577 3378 -571 3384
rect -205 3388 -201 3392
rect -277 3377 -271 3383
rect 95 3388 99 3392
rect 23 3378 29 3383
rect 695 3388 699 3393
rect 623 3378 629 3383
rect 995 3388 999 3392
rect 923 3377 929 3383
rect 1295 3388 1299 3392
rect 1223 3378 1229 3384
rect 2195 3388 2199 3392
rect 1523 3377 1529 3383
rect 1595 3377 1599 3382
rect 1895 3384 1899 3388
rect 1823 3378 1829 3384
rect 2123 3377 2129 3383
rect 2795 3386 2799 3390
rect -1492 3195 -1488 3199
rect -1483 3123 -1478 3129
rect -1482 2823 -1476 2829
rect -1482 2523 -1476 2529
rect -1482 2223 -1476 2229
rect -1478 2002 -1467 2098
rect 2723 3378 2729 3383
rect 3095 3386 3099 3390
rect 3023 3378 3029 3383
rect 3288 3195 3292 3199
rect 3277 3123 3283 3129
rect 3288 2895 3292 2899
rect 3276 2823 3282 2829
rect 3288 2595 3292 2599
rect 3001 2150 3006 2155
rect 3001 2120 3006 2125
rect 3001 2100 3006 2105
rect 3288 2295 3292 2299
rect 3276 2223 3282 2229
rect 2949 1666 2965 1751
rect 3288 1995 3292 1999
rect 3276 1923 3282 1929
rect 3256 1702 3276 1798
rect 3288 1395 3292 1399
rect -1492 1095 -1488 1099
rect -1483 1023 -1478 1029
rect -1483 723 -1478 729
rect -1483 423 -1478 429
rect -1480 202 -1471 298
rect -1482 71 -1476 77
rect -1482 -477 -1476 -471
rect -1483 -777 -1477 -771
rect -1483 -1077 -1477 -1071
rect -1220 1110 -1215 1115
rect 3288 1095 3292 1099
rect 3288 795 3292 799
rect 3288 495 3292 499
rect 3288 195 3292 199
rect 2948 -136 2966 -50
rect 3277 -98 3283 -2
rect 3288 -405 3292 -401
rect 3288 -705 3292 -701
rect 3276 -1077 3282 -1071
rect -1482 -1382 -1471 -1371
rect -1177 -1382 -1171 -1376
rect -877 -1382 -871 -1376
rect -577 -1382 -571 -1376
rect 23 -1382 29 -1376
rect 323 -1382 329 -1376
rect 623 -1382 629 -1376
rect 923 -1382 929 -1376
rect 1223 -1382 1229 -1376
rect 1823 -1382 1829 -1376
rect 2123 -1382 2129 -1376
rect 2423 -1382 2429 -1376
rect 2723 -1382 2729 -1376
rect 3023 -1382 3029 -1376
rect 3277 -1377 3283 -1371
<< metal3 >>
rect 694 3393 700 3395
rect -1407 3392 -1399 3393
rect -1407 3388 -1405 3392
rect -1401 3388 -1399 3392
rect -1478 3384 -1470 3385
rect -1478 3378 -1477 3384
rect -1471 3378 -1470 3384
rect -1478 3341 -1470 3378
rect -1407 3341 -1399 3388
rect -1106 3392 -1100 3393
rect -1106 3388 -1105 3392
rect -1101 3388 -1100 3392
rect -1178 3383 -1170 3384
rect -1178 3378 -1177 3383
rect -1171 3378 -1170 3383
rect -1178 3341 -1170 3378
rect -1106 3341 -1100 3388
rect -806 3392 -800 3393
rect -806 3388 -805 3392
rect -801 3388 -800 3392
rect -878 3383 -870 3384
rect -878 3377 -877 3383
rect -871 3377 -870 3383
rect -878 3341 -870 3377
rect -806 3341 -800 3388
rect -506 3392 -500 3393
rect -506 3387 -505 3392
rect -501 3387 -500 3392
rect -578 3384 -570 3385
rect -578 3378 -577 3384
rect -571 3378 -570 3384
rect -578 3341 -570 3378
rect -506 3341 -500 3387
rect -206 3392 -200 3393
rect -206 3388 -205 3392
rect -201 3388 -200 3392
rect -278 3383 -270 3384
rect -278 3377 -277 3383
rect -271 3377 -270 3383
rect -278 3341 -270 3377
rect -206 3341 -200 3388
rect 94 3392 100 3393
rect 94 3388 95 3392
rect 99 3388 100 3392
rect 22 3383 30 3384
rect 22 3378 23 3383
rect 29 3378 30 3383
rect 22 3341 30 3378
rect 94 3341 100 3388
rect 694 3388 695 3393
rect 699 3388 700 3393
rect 622 3383 630 3384
rect 622 3378 623 3383
rect 629 3378 630 3383
rect 622 3341 630 3378
rect 694 3341 700 3388
rect 994 3392 1000 3393
rect 994 3388 995 3392
rect 999 3388 1000 3392
rect 922 3383 930 3384
rect 922 3377 923 3383
rect 929 3377 930 3383
rect 922 3341 930 3377
rect 994 3341 1000 3388
rect 1294 3392 1300 3393
rect 1294 3388 1295 3392
rect 1299 3388 1300 3392
rect 2194 3392 2200 3393
rect 1222 3384 1230 3385
rect 1222 3378 1223 3384
rect 1229 3378 1230 3384
rect 1222 3341 1230 3378
rect 1294 3341 1300 3388
rect 1894 3388 1900 3389
rect 1522 3383 1530 3385
rect 1822 3384 1830 3385
rect 1522 3377 1523 3383
rect 1529 3377 1530 3383
rect 1522 3341 1530 3377
rect 1594 3382 1600 3383
rect 1594 3377 1595 3382
rect 1599 3377 1600 3382
rect 1594 3341 1600 3377
rect 1822 3378 1823 3384
rect 1829 3378 1830 3384
rect 1822 3341 1830 3378
rect 1894 3384 1895 3388
rect 1899 3384 1900 3388
rect 2194 3388 2195 3392
rect 2199 3388 2200 3392
rect 1894 3341 1900 3384
rect 2122 3383 2130 3384
rect 2122 3377 2123 3383
rect 2129 3377 2130 3383
rect 2122 3341 2130 3377
rect 2194 3341 2200 3388
rect 2794 3390 2800 3391
rect 2794 3386 2795 3390
rect 2799 3386 2800 3390
rect 2722 3383 2730 3385
rect 2722 3378 2723 3383
rect 2729 3378 2730 3383
rect 2722 3341 2730 3378
rect 2794 3341 2800 3386
rect 3094 3390 3100 3391
rect 3094 3386 3095 3390
rect 3099 3386 3100 3390
rect 3022 3383 3030 3384
rect 3022 3378 3023 3383
rect 3029 3378 3030 3383
rect 3022 3341 3030 3378
rect 3094 3341 3100 3386
rect -1478 3334 3246 3341
rect -1454 3289 3246 3334
rect -1454 3288 -1293 3289
rect -1454 3201 -1396 3288
rect -1313 3201 -1299 3288
rect -1493 3199 -1299 3201
rect -1493 3195 -1492 3199
rect -1488 3195 -1299 3199
rect -1493 3193 -1299 3195
rect 3175 3200 3246 3289
rect 3175 3199 3293 3200
rect 3175 3195 3288 3199
rect 3292 3195 3293 3199
rect 3175 3194 3293 3195
rect -1454 3130 -1396 3193
rect -1484 3129 -1396 3130
rect -1484 3123 -1483 3129
rect -1478 3123 -1396 3129
rect -1484 3122 -1396 3123
rect -1454 2830 -1396 3122
rect -1483 2829 -1396 2830
rect -1483 2823 -1482 2829
rect -1476 2823 -1396 2829
rect -1483 2822 -1396 2823
rect -1454 2530 -1396 2822
rect -1483 2529 -1396 2530
rect -1483 2523 -1482 2529
rect -1476 2523 -1396 2529
rect -1483 2522 -1396 2523
rect -1454 2230 -1396 2522
rect -1483 2229 -1396 2230
rect -1483 2223 -1482 2229
rect -1476 2223 -1396 2229
rect -1483 2222 -1396 2223
rect -1454 2099 -1396 2222
rect 3175 3130 3246 3194
rect 3175 3129 3284 3130
rect 3175 3123 3277 3129
rect 3283 3123 3284 3129
rect 3175 3122 3284 3123
rect 3175 2900 3246 3122
rect 3175 2899 3293 2900
rect 3175 2895 3288 2899
rect 3292 2895 3293 2899
rect 3175 2894 3293 2895
rect 3175 2830 3246 2894
rect 3175 2829 3283 2830
rect 3175 2823 3276 2829
rect 3282 2823 3283 2829
rect 3175 2822 3283 2823
rect 3175 2600 3246 2822
rect 3175 2599 3293 2600
rect 3175 2595 3288 2599
rect 3292 2595 3293 2599
rect 3175 2594 3293 2595
rect 3175 2300 3246 2594
rect 3175 2299 3293 2300
rect 3175 2295 3288 2299
rect 3292 2295 3293 2299
rect 3175 2294 3293 2295
rect 3175 2230 3246 2294
rect 3175 2229 3283 2230
rect 3175 2223 3276 2229
rect 3282 2223 3283 2229
rect 3175 2222 3283 2223
rect 3000 2155 3007 2156
rect 3000 2150 3001 2155
rect 3006 2150 3007 2155
rect 3000 2149 3007 2150
rect 3000 2125 3007 2126
rect 3000 2120 3001 2125
rect 3006 2120 3007 2125
rect 3000 2119 3007 2120
rect 3000 2105 3007 2106
rect 3000 2100 3001 2105
rect 3006 2100 3007 2105
rect 3000 2099 3007 2100
rect -1479 2098 -1396 2099
rect -1479 2002 -1478 2098
rect -1467 2002 -1396 2098
rect -1479 2001 -1396 2002
rect -1454 1100 -1396 2001
rect 3175 2000 3246 2222
rect 3175 1999 3293 2000
rect 3175 1995 3288 1999
rect 3292 1995 3293 1999
rect 3175 1994 3293 1995
rect 3175 1930 3246 1994
rect 3175 1929 3283 1930
rect 3175 1923 3276 1929
rect 3282 1923 3283 1929
rect 3175 1922 3283 1923
rect 3175 1799 3246 1922
rect 3175 1798 3277 1799
rect 3175 1752 3256 1798
rect 2948 1751 3256 1752
rect 2948 1666 2949 1751
rect 2965 1702 3256 1751
rect 3276 1702 3277 1798
rect 2965 1701 3277 1702
rect 2965 1666 3246 1701
rect 2948 1665 3246 1666
rect 3175 1400 3246 1665
rect 3175 1399 3293 1400
rect 3175 1395 3288 1399
rect 3292 1395 3293 1399
rect 3175 1394 3293 1395
rect -1221 1115 -1214 1116
rect -1221 1110 -1220 1115
rect -1215 1110 -1214 1115
rect -1221 1109 -1214 1110
rect -1493 1099 -1396 1100
rect -1493 1095 -1492 1099
rect -1488 1095 -1396 1099
rect -1493 1094 -1396 1095
rect -1454 1030 -1396 1094
rect -1484 1029 -1396 1030
rect -1484 1023 -1483 1029
rect -1478 1023 -1396 1029
rect -1484 1022 -1396 1023
rect -1454 730 -1396 1022
rect -1484 729 -1396 730
rect -1484 723 -1483 729
rect -1478 723 -1396 729
rect -1484 722 -1396 723
rect -1454 430 -1396 722
rect -1484 429 -1396 430
rect -1484 423 -1483 429
rect -1478 423 -1396 429
rect -1484 422 -1396 423
rect -1454 299 -1396 422
rect -1481 298 -1396 299
rect -1481 202 -1480 298
rect -1471 202 -1396 298
rect -1481 201 -1396 202
rect -1454 78 -1396 201
rect -1483 77 -1396 78
rect -1483 71 -1482 77
rect -1476 71 -1396 77
rect -1483 70 -1396 71
rect -1454 -470 -1396 70
rect 3175 1100 3246 1394
rect 3175 1099 3293 1100
rect 3175 1095 3288 1099
rect 3292 1095 3293 1099
rect 3175 1094 3293 1095
rect 3175 800 3246 1094
rect 3175 799 3293 800
rect 3175 795 3288 799
rect 3292 795 3293 799
rect 3175 794 3293 795
rect 3175 500 3246 794
rect 3175 499 3293 500
rect 3175 495 3288 499
rect 3292 495 3293 499
rect 3175 494 3293 495
rect 3175 200 3246 494
rect 3175 199 3293 200
rect 3175 195 3288 199
rect 3292 195 3293 199
rect 3175 194 3293 195
rect 3175 -1 3246 194
rect 3175 -2 3284 -1
rect 3175 -49 3277 -2
rect 2947 -50 3277 -49
rect 2947 -136 2948 -50
rect 2966 -98 3277 -50
rect 3283 -98 3284 -2
rect 2966 -99 3284 -98
rect 2966 -136 3246 -99
rect 2947 -137 3246 -136
rect -1483 -471 -1396 -470
rect -1483 -477 -1482 -471
rect -1476 -477 -1396 -471
rect -1483 -478 -1396 -477
rect -1454 -770 -1396 -478
rect -1484 -771 -1396 -770
rect -1484 -777 -1483 -771
rect -1477 -777 -1396 -771
rect -1484 -778 -1396 -777
rect -1454 -1070 -1396 -778
rect -1484 -1071 -1396 -1070
rect -1484 -1077 -1483 -1071
rect -1477 -1077 -1396 -1071
rect -1484 -1078 -1396 -1077
rect -1454 -1294 -1396 -1078
rect 3175 -400 3246 -137
rect 3175 -401 3293 -400
rect 3175 -405 3288 -401
rect 3292 -405 3293 -401
rect 3175 -406 3293 -405
rect 3175 -700 3246 -406
rect 3175 -701 3293 -700
rect 3175 -705 3288 -701
rect 3292 -705 3293 -701
rect 3175 -706 3293 -705
rect 3175 -1070 3246 -706
rect 3175 -1071 3283 -1070
rect 3175 -1077 3276 -1071
rect 3282 -1077 3283 -1071
rect 3175 -1078 3283 -1077
rect 3175 -1294 3246 -1078
rect -1454 -1351 3246 -1294
rect -1444 -1370 -1439 -1351
rect -1483 -1371 -1439 -1370
rect -1483 -1382 -1482 -1371
rect -1471 -1375 -1439 -1371
rect -1471 -1382 -1470 -1375
rect -1483 -1383 -1470 -1382
rect -1178 -1376 -1170 -1351
rect -1178 -1382 -1177 -1376
rect -1171 -1382 -1170 -1376
rect -1178 -1383 -1170 -1382
rect -878 -1376 -870 -1351
rect -878 -1382 -877 -1376
rect -871 -1382 -870 -1376
rect -878 -1383 -870 -1382
rect -578 -1376 -570 -1351
rect -578 -1382 -577 -1376
rect -571 -1382 -570 -1376
rect -578 -1383 -570 -1382
rect 22 -1376 30 -1351
rect 22 -1382 23 -1376
rect 29 -1382 30 -1376
rect 22 -1383 30 -1382
rect 322 -1376 330 -1351
rect 322 -1382 323 -1376
rect 329 -1382 330 -1376
rect 322 -1383 330 -1382
rect 622 -1376 630 -1351
rect 622 -1382 623 -1376
rect 629 -1382 630 -1376
rect 622 -1383 630 -1382
rect 922 -1376 930 -1351
rect 922 -1382 923 -1376
rect 929 -1382 930 -1376
rect 922 -1383 930 -1382
rect 1222 -1376 1230 -1351
rect 1222 -1382 1223 -1376
rect 1229 -1382 1230 -1376
rect 1222 -1383 1230 -1382
rect 1822 -1376 1830 -1351
rect 1822 -1382 1823 -1376
rect 1829 -1382 1830 -1376
rect 1822 -1383 1830 -1382
rect 2122 -1376 2130 -1351
rect 2122 -1382 2123 -1376
rect 2129 -1382 2130 -1376
rect 2122 -1383 2130 -1382
rect 2422 -1376 2430 -1351
rect 2422 -1382 2423 -1376
rect 2429 -1382 2430 -1376
rect 2422 -1383 2430 -1382
rect 2722 -1376 2730 -1351
rect 2722 -1382 2723 -1376
rect 2729 -1382 2730 -1376
rect 2722 -1383 2730 -1382
rect 3022 -1376 3030 -1351
rect 3022 -1382 3023 -1376
rect 3029 -1382 3030 -1376
rect 3237 -1370 3246 -1351
rect 3237 -1371 3284 -1370
rect 3237 -1377 3277 -1371
rect 3283 -1377 3284 -1371
rect 3237 -1378 3284 -1377
rect 3022 -1383 3030 -1382
use top_level  top_level_0
timestamp 1680464795
transform 1 0 -1220 0 1 -1212
box 0 12 4226 4140
use PadFrame64  PadFrame64_0
timestamp 1681001061
transform 1 0 0 0 1 0
box -2500 -2400 4300 4400
<< labels >>
rlabel m2contact 3282 3361 3282 3361 3 17_17_DI
rlabel metal2 3282 3348 3282 3348 3 17_17_DIB
rlabel metal1 -2206 249 -2206 249 1 Gnd!
rlabel metal1 447 4108 447 4108 1 Vdd!
rlabel metal1 -2207 2051 -2207 2051 1 Gnd!
rlabel metal1 -2212 1154 -2212 1154 1 p_clkb
rlabel metal1 -2212 3250 -2212 3250 1 p_load[8]
rlabel metal1 -1352 4113 -1352 4113 1 p_load[0]
rlabel metal1 -1047 4106 -1047 4106 1 p_load[14]
rlabel metal1 -753 4109 -753 4109 1 p_load[12]
rlabel metal1 -448 4112 -448 4112 1 p_load[13]
rlabel metal1 -145 4112 -145 4112 1 p_load[9]
rlabel metal1 153 4115 153 4115 1 p_load[7]
rlabel metal1 754 4109 754 4109 1 p_load[3]
rlabel metal1 1055 4112 1055 4112 1 p_load[10]
rlabel metal1 1353 4109 1353 4109 1 p_load[5]
rlabel metal1 1660 4112 1660 4112 1 p_load[11]
rlabel metal1 1952 4114 1952 4114 1 p_load[6]
rlabel metal1 2254 4113 2254 4113 1 p_load[15]
rlabel metal1 2549 4110 2549 4110 1 Vdd!
rlabel metal1 2846 4106 2846 4106 1 p_load[2]
rlabel metal1 3145 4106 3145 4106 1 p_load[1]
rlabel metal1 4006 3244 4006 3244 1 p_we_ins
rlabel metal1 4001 2946 4001 2946 1 p_load[4]
rlabel metal1 4010 2655 4010 2655 1 p_reg_0_out[7]
rlabel metal1 4011 2345 4011 2345 1 p_clka
rlabel metal1 4015 2053 4015 2053 1 p_reset
rlabel metal1 4013 1453 4013 1453 1 p_reg_0_out[1]
rlabel metal1 4007 1757 4007 1757 1 Gnd!
rlabel metal1 4013 1151 4013 1151 1 p_reg_0_out[0]
rlabel metal1 4008 848 4008 848 1 p_reg_0_out[6]
rlabel metal1 4008 557 4008 557 1 p_reg_0_out[2]
rlabel metal1 4007 253 4007 253 1 p_reg_0_out[3]
rlabel metal1 4008 -350 4008 -350 1 p_reg_0_out[5]
rlabel metal1 4009 -645 4009 -645 1 p_reg_0_out[4]
rlabel metal1 4002 -48 4002 -48 1 Gnd!
<< end >>

magic
tech scmos
timestamp 1682952543
<< nwell >>
rect 671 246 1003 330
rect 670 -3 1003 246
<< psubstratepdiff >>
rect 330 344 1000 670
rect 330 0 655 344
<< nsubstratendiff >>
rect 674 89 1000 327
rect 673 0 1000 89
<< genericcontact >>
rect 331 667 333 669
rect 336 667 338 669
rect 341 667 343 669
rect 346 667 348 669
rect 351 667 353 669
rect 356 667 358 669
rect 361 667 363 669
rect 366 667 368 669
rect 371 667 373 669
rect 376 667 378 669
rect 381 667 383 669
rect 386 667 388 669
rect 391 667 393 669
rect 396 667 398 669
rect 401 667 403 669
rect 406 667 408 669
rect 411 667 413 669
rect 416 667 418 669
rect 421 667 423 669
rect 426 667 428 669
rect 431 667 433 669
rect 436 667 438 669
rect 441 667 443 669
rect 446 667 448 669
rect 451 667 453 669
rect 456 667 458 669
rect 461 667 463 669
rect 466 667 468 669
rect 471 667 473 669
rect 476 667 478 669
rect 481 667 483 669
rect 486 667 488 669
rect 491 667 493 669
rect 496 667 498 669
rect 501 667 503 669
rect 506 667 508 669
rect 511 667 513 669
rect 516 667 518 669
rect 521 667 523 669
rect 526 667 528 669
rect 531 667 533 669
rect 536 667 538 669
rect 541 667 543 669
rect 546 667 548 669
rect 551 667 553 669
rect 556 667 558 669
rect 561 667 563 669
rect 566 667 568 669
rect 571 667 573 669
rect 576 667 578 669
rect 581 667 583 669
rect 586 667 588 669
rect 591 667 593 669
rect 596 667 598 669
rect 601 667 603 669
rect 606 667 608 669
rect 611 667 613 669
rect 616 667 618 669
rect 621 667 623 669
rect 626 667 628 669
rect 631 667 633 669
rect 636 667 638 669
rect 641 667 643 669
rect 646 667 648 669
rect 651 667 653 669
rect 656 667 658 669
rect 661 667 663 669
rect 666 667 668 669
rect 671 667 673 669
rect 676 667 678 669
rect 681 667 683 669
rect 686 667 688 669
rect 691 667 693 669
rect 696 667 698 669
rect 701 667 703 669
rect 706 667 708 669
rect 711 667 713 669
rect 716 667 718 669
rect 721 667 723 669
rect 726 667 728 669
rect 731 667 733 669
rect 736 667 738 669
rect 741 667 743 669
rect 746 667 748 669
rect 751 667 753 669
rect 756 667 758 669
rect 761 667 763 669
rect 766 667 768 669
rect 771 667 773 669
rect 776 667 778 669
rect 781 667 783 669
rect 786 667 788 669
rect 791 667 793 669
rect 796 667 798 669
rect 801 667 803 669
rect 806 667 808 669
rect 811 667 813 669
rect 816 667 818 669
rect 821 667 823 669
rect 826 667 828 669
rect 831 667 833 669
rect 836 667 838 669
rect 841 667 843 669
rect 846 667 848 669
rect 851 667 853 669
rect 856 667 858 669
rect 861 667 863 669
rect 866 667 868 669
rect 871 667 873 669
rect 876 667 878 669
rect 881 667 883 669
rect 886 667 888 669
rect 891 667 893 669
rect 896 667 898 669
rect 901 667 903 669
rect 906 667 908 669
rect 911 667 913 669
rect 916 667 918 669
rect 921 667 923 669
rect 926 667 928 669
rect 931 667 933 669
rect 936 667 938 669
rect 941 667 943 669
rect 946 667 948 669
rect 951 667 953 669
rect 956 667 958 669
rect 961 667 963 669
rect 966 667 968 669
rect 971 667 973 669
rect 976 667 978 669
rect 981 667 983 669
rect 986 667 988 669
rect 991 667 993 669
rect 996 667 998 669
rect 331 662 333 664
rect 336 662 338 664
rect 341 662 343 664
rect 346 662 348 664
rect 351 662 353 664
rect 356 662 358 664
rect 361 662 363 664
rect 366 662 368 664
rect 371 662 373 664
rect 376 662 378 664
rect 381 662 383 664
rect 386 662 388 664
rect 391 662 393 664
rect 396 662 398 664
rect 401 662 403 664
rect 406 662 408 664
rect 411 662 413 664
rect 416 662 418 664
rect 421 662 423 664
rect 426 662 428 664
rect 431 662 433 664
rect 436 662 438 664
rect 441 662 443 664
rect 446 662 448 664
rect 451 662 453 664
rect 456 662 458 664
rect 461 662 463 664
rect 466 662 468 664
rect 471 662 473 664
rect 476 662 478 664
rect 481 662 483 664
rect 486 662 488 664
rect 491 662 493 664
rect 496 662 498 664
rect 501 662 503 664
rect 506 662 508 664
rect 511 662 513 664
rect 516 662 518 664
rect 521 662 523 664
rect 526 662 528 664
rect 531 662 533 664
rect 536 662 538 664
rect 541 662 543 664
rect 546 662 548 664
rect 551 662 553 664
rect 556 662 558 664
rect 561 662 563 664
rect 566 662 568 664
rect 571 662 573 664
rect 576 662 578 664
rect 581 662 583 664
rect 586 662 588 664
rect 591 662 593 664
rect 596 662 598 664
rect 601 662 603 664
rect 606 662 608 664
rect 611 662 613 664
rect 616 662 618 664
rect 621 662 623 664
rect 626 662 628 664
rect 631 662 633 664
rect 636 662 638 664
rect 641 662 643 664
rect 646 662 648 664
rect 651 662 653 664
rect 656 662 658 664
rect 661 662 663 664
rect 666 662 668 664
rect 671 662 673 664
rect 676 662 678 664
rect 681 662 683 664
rect 686 662 688 664
rect 691 662 693 664
rect 696 662 698 664
rect 701 662 703 664
rect 706 662 708 664
rect 711 662 713 664
rect 716 662 718 664
rect 721 662 723 664
rect 726 662 728 664
rect 731 662 733 664
rect 736 662 738 664
rect 741 662 743 664
rect 746 662 748 664
rect 751 662 753 664
rect 756 662 758 664
rect 761 662 763 664
rect 766 662 768 664
rect 771 662 773 664
rect 776 662 778 664
rect 781 662 783 664
rect 786 662 788 664
rect 791 662 793 664
rect 796 662 798 664
rect 801 662 803 664
rect 806 662 808 664
rect 811 662 813 664
rect 816 662 818 664
rect 821 662 823 664
rect 826 662 828 664
rect 831 662 833 664
rect 836 662 838 664
rect 841 662 843 664
rect 846 662 848 664
rect 851 662 853 664
rect 856 662 858 664
rect 861 662 863 664
rect 866 662 868 664
rect 871 662 873 664
rect 876 662 878 664
rect 881 662 883 664
rect 886 662 888 664
rect 891 662 893 664
rect 896 662 898 664
rect 901 662 903 664
rect 906 662 908 664
rect 911 662 913 664
rect 916 662 918 664
rect 921 662 923 664
rect 926 662 928 664
rect 931 662 933 664
rect 936 662 938 664
rect 941 662 943 664
rect 946 662 948 664
rect 951 662 953 664
rect 956 662 958 664
rect 961 662 963 664
rect 966 662 968 664
rect 971 662 973 664
rect 976 662 978 664
rect 981 662 983 664
rect 986 662 988 664
rect 991 662 993 664
rect 996 662 998 664
rect 331 657 333 659
rect 336 657 338 659
rect 341 657 343 659
rect 346 657 348 659
rect 351 657 353 659
rect 356 657 358 659
rect 361 657 363 659
rect 366 657 368 659
rect 371 657 373 659
rect 376 657 378 659
rect 381 657 383 659
rect 386 657 388 659
rect 391 657 393 659
rect 396 657 398 659
rect 401 657 403 659
rect 406 657 408 659
rect 411 657 413 659
rect 416 657 418 659
rect 421 657 423 659
rect 426 657 428 659
rect 431 657 433 659
rect 436 657 438 659
rect 441 657 443 659
rect 446 657 448 659
rect 451 657 453 659
rect 456 657 458 659
rect 461 657 463 659
rect 466 657 468 659
rect 471 657 473 659
rect 476 657 478 659
rect 481 657 483 659
rect 486 657 488 659
rect 491 657 493 659
rect 496 657 498 659
rect 501 657 503 659
rect 506 657 508 659
rect 511 657 513 659
rect 516 657 518 659
rect 521 657 523 659
rect 526 657 528 659
rect 531 657 533 659
rect 536 657 538 659
rect 541 657 543 659
rect 546 657 548 659
rect 551 657 553 659
rect 556 657 558 659
rect 561 657 563 659
rect 566 657 568 659
rect 571 657 573 659
rect 576 657 578 659
rect 581 657 583 659
rect 586 657 588 659
rect 591 657 593 659
rect 596 657 598 659
rect 601 657 603 659
rect 606 657 608 659
rect 611 657 613 659
rect 616 657 618 659
rect 621 657 623 659
rect 626 657 628 659
rect 631 657 633 659
rect 636 657 638 659
rect 641 657 643 659
rect 646 657 648 659
rect 651 657 653 659
rect 656 657 658 659
rect 661 657 663 659
rect 666 657 668 659
rect 671 657 673 659
rect 676 657 678 659
rect 681 657 683 659
rect 686 657 688 659
rect 691 657 693 659
rect 696 657 698 659
rect 701 657 703 659
rect 706 657 708 659
rect 711 657 713 659
rect 716 657 718 659
rect 721 657 723 659
rect 726 657 728 659
rect 731 657 733 659
rect 736 657 738 659
rect 741 657 743 659
rect 746 657 748 659
rect 751 657 753 659
rect 756 657 758 659
rect 761 657 763 659
rect 766 657 768 659
rect 771 657 773 659
rect 776 657 778 659
rect 781 657 783 659
rect 786 657 788 659
rect 791 657 793 659
rect 796 657 798 659
rect 801 657 803 659
rect 806 657 808 659
rect 811 657 813 659
rect 816 657 818 659
rect 821 657 823 659
rect 826 657 828 659
rect 831 657 833 659
rect 836 657 838 659
rect 841 657 843 659
rect 846 657 848 659
rect 851 657 853 659
rect 856 657 858 659
rect 861 657 863 659
rect 866 657 868 659
rect 871 657 873 659
rect 876 657 878 659
rect 881 657 883 659
rect 886 657 888 659
rect 891 657 893 659
rect 896 657 898 659
rect 901 657 903 659
rect 906 657 908 659
rect 911 657 913 659
rect 916 657 918 659
rect 921 657 923 659
rect 926 657 928 659
rect 931 657 933 659
rect 936 657 938 659
rect 941 657 943 659
rect 946 657 948 659
rect 951 657 953 659
rect 956 657 958 659
rect 961 657 963 659
rect 966 657 968 659
rect 971 657 973 659
rect 976 657 978 659
rect 981 657 983 659
rect 986 657 988 659
rect 991 657 993 659
rect 996 657 998 659
rect 331 652 333 654
rect 336 652 338 654
rect 341 652 343 654
rect 346 652 348 654
rect 351 652 353 654
rect 356 652 358 654
rect 361 652 363 654
rect 366 652 368 654
rect 371 652 373 654
rect 376 652 378 654
rect 381 652 383 654
rect 386 652 388 654
rect 391 652 393 654
rect 396 652 398 654
rect 401 652 403 654
rect 406 652 408 654
rect 411 652 413 654
rect 416 652 418 654
rect 421 652 423 654
rect 426 652 428 654
rect 431 652 433 654
rect 436 652 438 654
rect 441 652 443 654
rect 446 652 448 654
rect 451 652 453 654
rect 456 652 458 654
rect 461 652 463 654
rect 466 652 468 654
rect 471 652 473 654
rect 476 652 478 654
rect 481 652 483 654
rect 486 652 488 654
rect 491 652 493 654
rect 496 652 498 654
rect 501 652 503 654
rect 506 652 508 654
rect 511 652 513 654
rect 516 652 518 654
rect 521 652 523 654
rect 526 652 528 654
rect 531 652 533 654
rect 536 652 538 654
rect 541 652 543 654
rect 546 652 548 654
rect 551 652 553 654
rect 556 652 558 654
rect 561 652 563 654
rect 566 652 568 654
rect 571 652 573 654
rect 576 652 578 654
rect 581 652 583 654
rect 586 652 588 654
rect 591 652 593 654
rect 596 652 598 654
rect 601 652 603 654
rect 606 652 608 654
rect 611 652 613 654
rect 616 652 618 654
rect 621 652 623 654
rect 626 652 628 654
rect 631 652 633 654
rect 636 652 638 654
rect 641 652 643 654
rect 646 652 648 654
rect 651 652 653 654
rect 656 652 658 654
rect 661 652 663 654
rect 666 652 668 654
rect 671 652 673 654
rect 676 652 678 654
rect 681 652 683 654
rect 686 652 688 654
rect 691 652 693 654
rect 696 652 698 654
rect 701 652 703 654
rect 706 652 708 654
rect 711 652 713 654
rect 716 652 718 654
rect 721 652 723 654
rect 726 652 728 654
rect 731 652 733 654
rect 736 652 738 654
rect 741 652 743 654
rect 746 652 748 654
rect 751 652 753 654
rect 756 652 758 654
rect 761 652 763 654
rect 766 652 768 654
rect 771 652 773 654
rect 776 652 778 654
rect 781 652 783 654
rect 786 652 788 654
rect 791 652 793 654
rect 796 652 798 654
rect 801 652 803 654
rect 806 652 808 654
rect 811 652 813 654
rect 816 652 818 654
rect 821 652 823 654
rect 826 652 828 654
rect 831 652 833 654
rect 836 652 838 654
rect 841 652 843 654
rect 846 652 848 654
rect 851 652 853 654
rect 856 652 858 654
rect 861 652 863 654
rect 866 652 868 654
rect 871 652 873 654
rect 876 652 878 654
rect 881 652 883 654
rect 886 652 888 654
rect 891 652 893 654
rect 896 652 898 654
rect 901 652 903 654
rect 906 652 908 654
rect 911 652 913 654
rect 916 652 918 654
rect 921 652 923 654
rect 926 652 928 654
rect 931 652 933 654
rect 936 652 938 654
rect 941 652 943 654
rect 946 652 948 654
rect 951 652 953 654
rect 956 652 958 654
rect 961 652 963 654
rect 966 652 968 654
rect 971 652 973 654
rect 976 652 978 654
rect 981 652 983 654
rect 986 652 988 654
rect 991 652 993 654
rect 996 652 998 654
rect 331 647 333 649
rect 336 647 338 649
rect 341 647 343 649
rect 346 647 348 649
rect 351 647 353 649
rect 356 647 358 649
rect 361 647 363 649
rect 366 647 368 649
rect 371 647 373 649
rect 376 647 378 649
rect 381 647 383 649
rect 386 647 388 649
rect 391 647 393 649
rect 396 647 398 649
rect 401 647 403 649
rect 406 647 408 649
rect 411 647 413 649
rect 416 647 418 649
rect 421 647 423 649
rect 426 647 428 649
rect 431 647 433 649
rect 436 647 438 649
rect 441 647 443 649
rect 446 647 448 649
rect 451 647 453 649
rect 456 647 458 649
rect 461 647 463 649
rect 466 647 468 649
rect 471 647 473 649
rect 476 647 478 649
rect 481 647 483 649
rect 486 647 488 649
rect 491 647 493 649
rect 496 647 498 649
rect 501 647 503 649
rect 506 647 508 649
rect 511 647 513 649
rect 516 647 518 649
rect 521 647 523 649
rect 526 647 528 649
rect 531 647 533 649
rect 536 647 538 649
rect 541 647 543 649
rect 546 647 548 649
rect 551 647 553 649
rect 556 647 558 649
rect 561 647 563 649
rect 566 647 568 649
rect 571 647 573 649
rect 576 647 578 649
rect 581 647 583 649
rect 586 647 588 649
rect 591 647 593 649
rect 596 647 598 649
rect 601 647 603 649
rect 606 647 608 649
rect 611 647 613 649
rect 616 647 618 649
rect 621 647 623 649
rect 626 647 628 649
rect 631 647 633 649
rect 636 647 638 649
rect 641 647 643 649
rect 646 647 648 649
rect 651 647 653 649
rect 656 647 658 649
rect 661 647 663 649
rect 666 647 668 649
rect 671 647 673 649
rect 676 647 678 649
rect 681 647 683 649
rect 686 647 688 649
rect 691 647 693 649
rect 696 647 698 649
rect 701 647 703 649
rect 706 647 708 649
rect 711 647 713 649
rect 716 647 718 649
rect 721 647 723 649
rect 726 647 728 649
rect 731 647 733 649
rect 736 647 738 649
rect 741 647 743 649
rect 746 647 748 649
rect 751 647 753 649
rect 756 647 758 649
rect 761 647 763 649
rect 766 647 768 649
rect 771 647 773 649
rect 776 647 778 649
rect 781 647 783 649
rect 786 647 788 649
rect 791 647 793 649
rect 796 647 798 649
rect 801 647 803 649
rect 806 647 808 649
rect 811 647 813 649
rect 816 647 818 649
rect 821 647 823 649
rect 826 647 828 649
rect 831 647 833 649
rect 836 647 838 649
rect 841 647 843 649
rect 846 647 848 649
rect 851 647 853 649
rect 856 647 858 649
rect 861 647 863 649
rect 866 647 868 649
rect 871 647 873 649
rect 876 647 878 649
rect 881 647 883 649
rect 886 647 888 649
rect 891 647 893 649
rect 896 647 898 649
rect 901 647 903 649
rect 906 647 908 649
rect 911 647 913 649
rect 916 647 918 649
rect 921 647 923 649
rect 926 647 928 649
rect 931 647 933 649
rect 936 647 938 649
rect 941 647 943 649
rect 946 647 948 649
rect 951 647 953 649
rect 956 647 958 649
rect 961 647 963 649
rect 966 647 968 649
rect 971 647 973 649
rect 976 647 978 649
rect 981 647 983 649
rect 986 647 988 649
rect 991 647 993 649
rect 996 647 998 649
rect 331 642 333 644
rect 336 642 338 644
rect 341 642 343 644
rect 346 642 348 644
rect 351 642 353 644
rect 356 642 358 644
rect 361 642 363 644
rect 366 642 368 644
rect 371 642 373 644
rect 376 642 378 644
rect 381 642 383 644
rect 386 642 388 644
rect 391 642 393 644
rect 396 642 398 644
rect 401 642 403 644
rect 406 642 408 644
rect 411 642 413 644
rect 416 642 418 644
rect 421 642 423 644
rect 426 642 428 644
rect 431 642 433 644
rect 436 642 438 644
rect 441 642 443 644
rect 446 642 448 644
rect 451 642 453 644
rect 456 642 458 644
rect 461 642 463 644
rect 466 642 468 644
rect 471 642 473 644
rect 476 642 478 644
rect 481 642 483 644
rect 486 642 488 644
rect 491 642 493 644
rect 496 642 498 644
rect 501 642 503 644
rect 506 642 508 644
rect 511 642 513 644
rect 516 642 518 644
rect 521 642 523 644
rect 526 642 528 644
rect 531 642 533 644
rect 536 642 538 644
rect 541 642 543 644
rect 546 642 548 644
rect 551 642 553 644
rect 556 642 558 644
rect 561 642 563 644
rect 566 642 568 644
rect 571 642 573 644
rect 576 642 578 644
rect 581 642 583 644
rect 586 642 588 644
rect 591 642 593 644
rect 596 642 598 644
rect 601 642 603 644
rect 606 642 608 644
rect 611 642 613 644
rect 616 642 618 644
rect 621 642 623 644
rect 626 642 628 644
rect 631 642 633 644
rect 636 642 638 644
rect 641 642 643 644
rect 646 642 648 644
rect 651 642 653 644
rect 656 642 658 644
rect 661 642 663 644
rect 666 642 668 644
rect 671 642 673 644
rect 676 642 678 644
rect 681 642 683 644
rect 686 642 688 644
rect 691 642 693 644
rect 696 642 698 644
rect 701 642 703 644
rect 706 642 708 644
rect 711 642 713 644
rect 716 642 718 644
rect 721 642 723 644
rect 726 642 728 644
rect 731 642 733 644
rect 736 642 738 644
rect 741 642 743 644
rect 746 642 748 644
rect 751 642 753 644
rect 756 642 758 644
rect 761 642 763 644
rect 766 642 768 644
rect 771 642 773 644
rect 776 642 778 644
rect 781 642 783 644
rect 786 642 788 644
rect 791 642 793 644
rect 796 642 798 644
rect 801 642 803 644
rect 806 642 808 644
rect 811 642 813 644
rect 816 642 818 644
rect 821 642 823 644
rect 826 642 828 644
rect 831 642 833 644
rect 836 642 838 644
rect 841 642 843 644
rect 846 642 848 644
rect 851 642 853 644
rect 856 642 858 644
rect 861 642 863 644
rect 866 642 868 644
rect 871 642 873 644
rect 876 642 878 644
rect 881 642 883 644
rect 886 642 888 644
rect 891 642 893 644
rect 896 642 898 644
rect 901 642 903 644
rect 906 642 908 644
rect 911 642 913 644
rect 916 642 918 644
rect 921 642 923 644
rect 926 642 928 644
rect 931 642 933 644
rect 936 642 938 644
rect 941 642 943 644
rect 946 642 948 644
rect 951 642 953 644
rect 956 642 958 644
rect 961 642 963 644
rect 966 642 968 644
rect 971 642 973 644
rect 976 642 978 644
rect 981 642 983 644
rect 986 642 988 644
rect 991 642 993 644
rect 996 642 998 644
rect 331 637 333 639
rect 336 637 338 639
rect 341 637 343 639
rect 346 637 348 639
rect 351 637 353 639
rect 356 637 358 639
rect 361 637 363 639
rect 366 637 368 639
rect 371 637 373 639
rect 376 637 378 639
rect 381 637 383 639
rect 386 637 388 639
rect 391 637 393 639
rect 396 637 398 639
rect 401 637 403 639
rect 406 637 408 639
rect 411 637 413 639
rect 416 637 418 639
rect 421 637 423 639
rect 426 637 428 639
rect 431 637 433 639
rect 436 637 438 639
rect 441 637 443 639
rect 446 637 448 639
rect 451 637 453 639
rect 456 637 458 639
rect 461 637 463 639
rect 466 637 468 639
rect 471 637 473 639
rect 476 637 478 639
rect 481 637 483 639
rect 486 637 488 639
rect 491 637 493 639
rect 496 637 498 639
rect 501 637 503 639
rect 506 637 508 639
rect 511 637 513 639
rect 516 637 518 639
rect 521 637 523 639
rect 526 637 528 639
rect 531 637 533 639
rect 536 637 538 639
rect 541 637 543 639
rect 546 637 548 639
rect 551 637 553 639
rect 556 637 558 639
rect 561 637 563 639
rect 566 637 568 639
rect 571 637 573 639
rect 576 637 578 639
rect 581 637 583 639
rect 586 637 588 639
rect 591 637 593 639
rect 596 637 598 639
rect 601 637 603 639
rect 606 637 608 639
rect 611 637 613 639
rect 616 637 618 639
rect 621 637 623 639
rect 626 637 628 639
rect 631 637 633 639
rect 636 637 638 639
rect 641 637 643 639
rect 646 637 648 639
rect 651 637 653 639
rect 656 637 658 639
rect 661 637 663 639
rect 666 637 668 639
rect 671 637 673 639
rect 676 637 678 639
rect 681 637 683 639
rect 686 637 688 639
rect 691 637 693 639
rect 696 637 698 639
rect 701 637 703 639
rect 706 637 708 639
rect 711 637 713 639
rect 716 637 718 639
rect 721 637 723 639
rect 726 637 728 639
rect 731 637 733 639
rect 736 637 738 639
rect 741 637 743 639
rect 746 637 748 639
rect 751 637 753 639
rect 756 637 758 639
rect 761 637 763 639
rect 766 637 768 639
rect 771 637 773 639
rect 776 637 778 639
rect 781 637 783 639
rect 786 637 788 639
rect 791 637 793 639
rect 796 637 798 639
rect 801 637 803 639
rect 806 637 808 639
rect 811 637 813 639
rect 816 637 818 639
rect 821 637 823 639
rect 826 637 828 639
rect 831 637 833 639
rect 836 637 838 639
rect 841 637 843 639
rect 846 637 848 639
rect 851 637 853 639
rect 856 637 858 639
rect 861 637 863 639
rect 866 637 868 639
rect 871 637 873 639
rect 876 637 878 639
rect 881 637 883 639
rect 886 637 888 639
rect 891 637 893 639
rect 896 637 898 639
rect 901 637 903 639
rect 906 637 908 639
rect 911 637 913 639
rect 916 637 918 639
rect 921 637 923 639
rect 926 637 928 639
rect 931 637 933 639
rect 936 637 938 639
rect 941 637 943 639
rect 946 637 948 639
rect 951 637 953 639
rect 956 637 958 639
rect 961 637 963 639
rect 966 637 968 639
rect 971 637 973 639
rect 976 637 978 639
rect 981 637 983 639
rect 986 637 988 639
rect 991 637 993 639
rect 996 637 998 639
rect 331 632 333 634
rect 336 632 338 634
rect 341 632 343 634
rect 346 632 348 634
rect 351 632 353 634
rect 356 632 358 634
rect 361 632 363 634
rect 366 632 368 634
rect 371 632 373 634
rect 376 632 378 634
rect 381 632 383 634
rect 386 632 388 634
rect 391 632 393 634
rect 396 632 398 634
rect 401 632 403 634
rect 406 632 408 634
rect 411 632 413 634
rect 416 632 418 634
rect 421 632 423 634
rect 426 632 428 634
rect 431 632 433 634
rect 436 632 438 634
rect 441 632 443 634
rect 446 632 448 634
rect 451 632 453 634
rect 456 632 458 634
rect 461 632 463 634
rect 466 632 468 634
rect 471 632 473 634
rect 476 632 478 634
rect 481 632 483 634
rect 486 632 488 634
rect 491 632 493 634
rect 496 632 498 634
rect 501 632 503 634
rect 506 632 508 634
rect 511 632 513 634
rect 516 632 518 634
rect 521 632 523 634
rect 526 632 528 634
rect 531 632 533 634
rect 536 632 538 634
rect 541 632 543 634
rect 546 632 548 634
rect 551 632 553 634
rect 556 632 558 634
rect 561 632 563 634
rect 566 632 568 634
rect 571 632 573 634
rect 576 632 578 634
rect 581 632 583 634
rect 586 632 588 634
rect 591 632 593 634
rect 596 632 598 634
rect 601 632 603 634
rect 606 632 608 634
rect 611 632 613 634
rect 616 632 618 634
rect 621 632 623 634
rect 626 632 628 634
rect 631 632 633 634
rect 636 632 638 634
rect 641 632 643 634
rect 646 632 648 634
rect 651 632 653 634
rect 656 632 658 634
rect 661 632 663 634
rect 666 632 668 634
rect 671 632 673 634
rect 676 632 678 634
rect 681 632 683 634
rect 686 632 688 634
rect 691 632 693 634
rect 696 632 698 634
rect 701 632 703 634
rect 706 632 708 634
rect 711 632 713 634
rect 716 632 718 634
rect 721 632 723 634
rect 726 632 728 634
rect 731 632 733 634
rect 736 632 738 634
rect 741 632 743 634
rect 746 632 748 634
rect 751 632 753 634
rect 756 632 758 634
rect 761 632 763 634
rect 766 632 768 634
rect 771 632 773 634
rect 776 632 778 634
rect 781 632 783 634
rect 786 632 788 634
rect 791 632 793 634
rect 796 632 798 634
rect 801 632 803 634
rect 806 632 808 634
rect 811 632 813 634
rect 816 632 818 634
rect 821 632 823 634
rect 826 632 828 634
rect 831 632 833 634
rect 836 632 838 634
rect 841 632 843 634
rect 846 632 848 634
rect 851 632 853 634
rect 856 632 858 634
rect 861 632 863 634
rect 866 632 868 634
rect 871 632 873 634
rect 876 632 878 634
rect 881 632 883 634
rect 886 632 888 634
rect 891 632 893 634
rect 896 632 898 634
rect 901 632 903 634
rect 906 632 908 634
rect 911 632 913 634
rect 916 632 918 634
rect 921 632 923 634
rect 926 632 928 634
rect 931 632 933 634
rect 936 632 938 634
rect 941 632 943 634
rect 946 632 948 634
rect 951 632 953 634
rect 956 632 958 634
rect 961 632 963 634
rect 966 632 968 634
rect 971 632 973 634
rect 976 632 978 634
rect 981 632 983 634
rect 986 632 988 634
rect 991 632 993 634
rect 996 632 998 634
rect 331 627 333 629
rect 336 627 338 629
rect 341 627 343 629
rect 346 627 348 629
rect 351 627 353 629
rect 356 627 358 629
rect 361 627 363 629
rect 366 627 368 629
rect 371 627 373 629
rect 376 627 378 629
rect 381 627 383 629
rect 386 627 388 629
rect 391 627 393 629
rect 396 627 398 629
rect 401 627 403 629
rect 406 627 408 629
rect 411 627 413 629
rect 416 627 418 629
rect 421 627 423 629
rect 426 627 428 629
rect 431 627 433 629
rect 436 627 438 629
rect 441 627 443 629
rect 446 627 448 629
rect 451 627 453 629
rect 456 627 458 629
rect 461 627 463 629
rect 466 627 468 629
rect 471 627 473 629
rect 476 627 478 629
rect 481 627 483 629
rect 486 627 488 629
rect 491 627 493 629
rect 496 627 498 629
rect 501 627 503 629
rect 506 627 508 629
rect 511 627 513 629
rect 516 627 518 629
rect 521 627 523 629
rect 526 627 528 629
rect 531 627 533 629
rect 536 627 538 629
rect 541 627 543 629
rect 546 627 548 629
rect 551 627 553 629
rect 556 627 558 629
rect 561 627 563 629
rect 566 627 568 629
rect 571 627 573 629
rect 576 627 578 629
rect 581 627 583 629
rect 586 627 588 629
rect 591 627 593 629
rect 596 627 598 629
rect 601 627 603 629
rect 606 627 608 629
rect 611 627 613 629
rect 616 627 618 629
rect 621 627 623 629
rect 626 627 628 629
rect 631 627 633 629
rect 636 627 638 629
rect 641 627 643 629
rect 646 627 648 629
rect 651 627 653 629
rect 656 627 658 629
rect 661 627 663 629
rect 666 627 668 629
rect 671 627 673 629
rect 676 627 678 629
rect 681 627 683 629
rect 686 627 688 629
rect 691 627 693 629
rect 696 627 698 629
rect 701 627 703 629
rect 706 627 708 629
rect 711 627 713 629
rect 716 627 718 629
rect 721 627 723 629
rect 726 627 728 629
rect 731 627 733 629
rect 736 627 738 629
rect 741 627 743 629
rect 746 627 748 629
rect 751 627 753 629
rect 756 627 758 629
rect 761 627 763 629
rect 766 627 768 629
rect 771 627 773 629
rect 776 627 778 629
rect 781 627 783 629
rect 786 627 788 629
rect 791 627 793 629
rect 796 627 798 629
rect 801 627 803 629
rect 806 627 808 629
rect 811 627 813 629
rect 816 627 818 629
rect 821 627 823 629
rect 826 627 828 629
rect 831 627 833 629
rect 836 627 838 629
rect 841 627 843 629
rect 846 627 848 629
rect 851 627 853 629
rect 856 627 858 629
rect 861 627 863 629
rect 866 627 868 629
rect 871 627 873 629
rect 876 627 878 629
rect 881 627 883 629
rect 886 627 888 629
rect 891 627 893 629
rect 896 627 898 629
rect 901 627 903 629
rect 906 627 908 629
rect 911 627 913 629
rect 916 627 918 629
rect 921 627 923 629
rect 926 627 928 629
rect 931 627 933 629
rect 936 627 938 629
rect 941 627 943 629
rect 946 627 948 629
rect 951 627 953 629
rect 956 627 958 629
rect 961 627 963 629
rect 966 627 968 629
rect 971 627 973 629
rect 976 627 978 629
rect 981 627 983 629
rect 986 627 988 629
rect 991 627 993 629
rect 996 627 998 629
rect 331 622 333 624
rect 336 622 338 624
rect 341 622 343 624
rect 346 622 348 624
rect 351 622 353 624
rect 356 622 358 624
rect 361 622 363 624
rect 366 622 368 624
rect 371 622 373 624
rect 376 622 378 624
rect 381 622 383 624
rect 386 622 388 624
rect 391 622 393 624
rect 396 622 398 624
rect 401 622 403 624
rect 406 622 408 624
rect 411 622 413 624
rect 416 622 418 624
rect 421 622 423 624
rect 426 622 428 624
rect 431 622 433 624
rect 436 622 438 624
rect 441 622 443 624
rect 446 622 448 624
rect 451 622 453 624
rect 456 622 458 624
rect 461 622 463 624
rect 466 622 468 624
rect 471 622 473 624
rect 476 622 478 624
rect 481 622 483 624
rect 486 622 488 624
rect 491 622 493 624
rect 496 622 498 624
rect 501 622 503 624
rect 506 622 508 624
rect 511 622 513 624
rect 516 622 518 624
rect 521 622 523 624
rect 526 622 528 624
rect 531 622 533 624
rect 536 622 538 624
rect 541 622 543 624
rect 546 622 548 624
rect 551 622 553 624
rect 556 622 558 624
rect 561 622 563 624
rect 566 622 568 624
rect 571 622 573 624
rect 576 622 578 624
rect 581 622 583 624
rect 586 622 588 624
rect 591 622 593 624
rect 596 622 598 624
rect 601 622 603 624
rect 606 622 608 624
rect 611 622 613 624
rect 616 622 618 624
rect 621 622 623 624
rect 626 622 628 624
rect 631 622 633 624
rect 636 622 638 624
rect 641 622 643 624
rect 646 622 648 624
rect 651 622 653 624
rect 656 622 658 624
rect 661 622 663 624
rect 666 622 668 624
rect 671 622 673 624
rect 676 622 678 624
rect 681 622 683 624
rect 686 622 688 624
rect 691 622 693 624
rect 696 622 698 624
rect 701 622 703 624
rect 706 622 708 624
rect 711 622 713 624
rect 716 622 718 624
rect 721 622 723 624
rect 726 622 728 624
rect 731 622 733 624
rect 736 622 738 624
rect 741 622 743 624
rect 746 622 748 624
rect 751 622 753 624
rect 756 622 758 624
rect 761 622 763 624
rect 766 622 768 624
rect 771 622 773 624
rect 776 622 778 624
rect 781 622 783 624
rect 786 622 788 624
rect 791 622 793 624
rect 796 622 798 624
rect 801 622 803 624
rect 806 622 808 624
rect 811 622 813 624
rect 816 622 818 624
rect 821 622 823 624
rect 826 622 828 624
rect 831 622 833 624
rect 836 622 838 624
rect 841 622 843 624
rect 846 622 848 624
rect 851 622 853 624
rect 856 622 858 624
rect 861 622 863 624
rect 866 622 868 624
rect 871 622 873 624
rect 876 622 878 624
rect 881 622 883 624
rect 886 622 888 624
rect 891 622 893 624
rect 896 622 898 624
rect 901 622 903 624
rect 906 622 908 624
rect 911 622 913 624
rect 916 622 918 624
rect 921 622 923 624
rect 926 622 928 624
rect 931 622 933 624
rect 936 622 938 624
rect 941 622 943 624
rect 946 622 948 624
rect 951 622 953 624
rect 956 622 958 624
rect 961 622 963 624
rect 966 622 968 624
rect 971 622 973 624
rect 976 622 978 624
rect 981 622 983 624
rect 986 622 988 624
rect 991 622 993 624
rect 996 622 998 624
rect 331 617 333 619
rect 336 617 338 619
rect 341 617 343 619
rect 346 617 348 619
rect 351 617 353 619
rect 356 617 358 619
rect 361 617 363 619
rect 366 617 368 619
rect 371 617 373 619
rect 376 617 378 619
rect 381 617 383 619
rect 386 617 388 619
rect 391 617 393 619
rect 396 617 398 619
rect 401 617 403 619
rect 406 617 408 619
rect 411 617 413 619
rect 416 617 418 619
rect 421 617 423 619
rect 426 617 428 619
rect 431 617 433 619
rect 436 617 438 619
rect 441 617 443 619
rect 446 617 448 619
rect 451 617 453 619
rect 456 617 458 619
rect 461 617 463 619
rect 466 617 468 619
rect 471 617 473 619
rect 476 617 478 619
rect 481 617 483 619
rect 486 617 488 619
rect 491 617 493 619
rect 496 617 498 619
rect 501 617 503 619
rect 506 617 508 619
rect 511 617 513 619
rect 516 617 518 619
rect 521 617 523 619
rect 526 617 528 619
rect 531 617 533 619
rect 536 617 538 619
rect 541 617 543 619
rect 546 617 548 619
rect 551 617 553 619
rect 556 617 558 619
rect 561 617 563 619
rect 566 617 568 619
rect 571 617 573 619
rect 576 617 578 619
rect 581 617 583 619
rect 586 617 588 619
rect 591 617 593 619
rect 596 617 598 619
rect 601 617 603 619
rect 606 617 608 619
rect 611 617 613 619
rect 616 617 618 619
rect 621 617 623 619
rect 626 617 628 619
rect 631 617 633 619
rect 636 617 638 619
rect 641 617 643 619
rect 646 617 648 619
rect 651 617 653 619
rect 656 617 658 619
rect 661 617 663 619
rect 666 617 668 619
rect 671 617 673 619
rect 676 617 678 619
rect 681 617 683 619
rect 686 617 688 619
rect 691 617 693 619
rect 696 617 698 619
rect 701 617 703 619
rect 706 617 708 619
rect 711 617 713 619
rect 716 617 718 619
rect 721 617 723 619
rect 726 617 728 619
rect 731 617 733 619
rect 736 617 738 619
rect 741 617 743 619
rect 746 617 748 619
rect 751 617 753 619
rect 756 617 758 619
rect 761 617 763 619
rect 766 617 768 619
rect 771 617 773 619
rect 776 617 778 619
rect 781 617 783 619
rect 786 617 788 619
rect 791 617 793 619
rect 796 617 798 619
rect 801 617 803 619
rect 806 617 808 619
rect 811 617 813 619
rect 816 617 818 619
rect 821 617 823 619
rect 826 617 828 619
rect 831 617 833 619
rect 836 617 838 619
rect 841 617 843 619
rect 846 617 848 619
rect 851 617 853 619
rect 856 617 858 619
rect 861 617 863 619
rect 866 617 868 619
rect 871 617 873 619
rect 876 617 878 619
rect 881 617 883 619
rect 886 617 888 619
rect 891 617 893 619
rect 896 617 898 619
rect 901 617 903 619
rect 906 617 908 619
rect 911 617 913 619
rect 916 617 918 619
rect 921 617 923 619
rect 926 617 928 619
rect 931 617 933 619
rect 936 617 938 619
rect 941 617 943 619
rect 946 617 948 619
rect 951 617 953 619
rect 956 617 958 619
rect 961 617 963 619
rect 966 617 968 619
rect 971 617 973 619
rect 976 617 978 619
rect 981 617 983 619
rect 986 617 988 619
rect 991 617 993 619
rect 996 617 998 619
rect 331 612 333 614
rect 336 612 338 614
rect 341 612 343 614
rect 346 612 348 614
rect 351 612 353 614
rect 356 612 358 614
rect 361 612 363 614
rect 366 612 368 614
rect 371 612 373 614
rect 376 612 378 614
rect 381 612 383 614
rect 386 612 388 614
rect 391 612 393 614
rect 396 612 398 614
rect 401 612 403 614
rect 406 612 408 614
rect 411 612 413 614
rect 416 612 418 614
rect 421 612 423 614
rect 426 612 428 614
rect 431 612 433 614
rect 436 612 438 614
rect 441 612 443 614
rect 446 612 448 614
rect 451 612 453 614
rect 456 612 458 614
rect 461 612 463 614
rect 466 612 468 614
rect 471 612 473 614
rect 476 612 478 614
rect 481 612 483 614
rect 486 612 488 614
rect 491 612 493 614
rect 496 612 498 614
rect 501 612 503 614
rect 506 612 508 614
rect 511 612 513 614
rect 516 612 518 614
rect 521 612 523 614
rect 526 612 528 614
rect 531 612 533 614
rect 536 612 538 614
rect 541 612 543 614
rect 546 612 548 614
rect 551 612 553 614
rect 556 612 558 614
rect 561 612 563 614
rect 566 612 568 614
rect 571 612 573 614
rect 576 612 578 614
rect 581 612 583 614
rect 586 612 588 614
rect 591 612 593 614
rect 596 612 598 614
rect 601 612 603 614
rect 606 612 608 614
rect 611 612 613 614
rect 616 612 618 614
rect 621 612 623 614
rect 626 612 628 614
rect 631 612 633 614
rect 636 612 638 614
rect 641 612 643 614
rect 646 612 648 614
rect 651 612 653 614
rect 656 612 658 614
rect 661 612 663 614
rect 666 612 668 614
rect 671 612 673 614
rect 676 612 678 614
rect 681 612 683 614
rect 686 612 688 614
rect 691 612 693 614
rect 696 612 698 614
rect 701 612 703 614
rect 706 612 708 614
rect 711 612 713 614
rect 716 612 718 614
rect 721 612 723 614
rect 726 612 728 614
rect 731 612 733 614
rect 736 612 738 614
rect 741 612 743 614
rect 746 612 748 614
rect 751 612 753 614
rect 756 612 758 614
rect 761 612 763 614
rect 766 612 768 614
rect 771 612 773 614
rect 776 612 778 614
rect 781 612 783 614
rect 786 612 788 614
rect 791 612 793 614
rect 796 612 798 614
rect 801 612 803 614
rect 806 612 808 614
rect 811 612 813 614
rect 816 612 818 614
rect 821 612 823 614
rect 826 612 828 614
rect 831 612 833 614
rect 836 612 838 614
rect 841 612 843 614
rect 846 612 848 614
rect 851 612 853 614
rect 856 612 858 614
rect 861 612 863 614
rect 866 612 868 614
rect 871 612 873 614
rect 876 612 878 614
rect 881 612 883 614
rect 886 612 888 614
rect 891 612 893 614
rect 896 612 898 614
rect 901 612 903 614
rect 906 612 908 614
rect 911 612 913 614
rect 916 612 918 614
rect 921 612 923 614
rect 926 612 928 614
rect 931 612 933 614
rect 936 612 938 614
rect 941 612 943 614
rect 946 612 948 614
rect 951 612 953 614
rect 956 612 958 614
rect 961 612 963 614
rect 966 612 968 614
rect 971 612 973 614
rect 976 612 978 614
rect 981 612 983 614
rect 986 612 988 614
rect 991 612 993 614
rect 996 612 998 614
rect 331 607 333 609
rect 336 607 338 609
rect 341 607 343 609
rect 346 607 348 609
rect 351 607 353 609
rect 356 607 358 609
rect 361 607 363 609
rect 366 607 368 609
rect 371 607 373 609
rect 376 607 378 609
rect 381 607 383 609
rect 386 607 388 609
rect 391 607 393 609
rect 396 607 398 609
rect 401 607 403 609
rect 406 607 408 609
rect 411 607 413 609
rect 416 607 418 609
rect 421 607 423 609
rect 426 607 428 609
rect 431 607 433 609
rect 436 607 438 609
rect 441 607 443 609
rect 446 607 448 609
rect 451 607 453 609
rect 456 607 458 609
rect 461 607 463 609
rect 466 607 468 609
rect 471 607 473 609
rect 476 607 478 609
rect 481 607 483 609
rect 486 607 488 609
rect 491 607 493 609
rect 496 607 498 609
rect 501 607 503 609
rect 506 607 508 609
rect 511 607 513 609
rect 516 607 518 609
rect 521 607 523 609
rect 526 607 528 609
rect 531 607 533 609
rect 536 607 538 609
rect 541 607 543 609
rect 546 607 548 609
rect 551 607 553 609
rect 556 607 558 609
rect 561 607 563 609
rect 566 607 568 609
rect 571 607 573 609
rect 576 607 578 609
rect 581 607 583 609
rect 586 607 588 609
rect 591 607 593 609
rect 596 607 598 609
rect 601 607 603 609
rect 606 607 608 609
rect 611 607 613 609
rect 616 607 618 609
rect 621 607 623 609
rect 626 607 628 609
rect 631 607 633 609
rect 636 607 638 609
rect 641 607 643 609
rect 646 607 648 609
rect 651 607 653 609
rect 656 607 658 609
rect 661 607 663 609
rect 666 607 668 609
rect 671 607 673 609
rect 676 607 678 609
rect 681 607 683 609
rect 686 607 688 609
rect 691 607 693 609
rect 696 607 698 609
rect 701 607 703 609
rect 706 607 708 609
rect 711 607 713 609
rect 716 607 718 609
rect 721 607 723 609
rect 726 607 728 609
rect 731 607 733 609
rect 736 607 738 609
rect 741 607 743 609
rect 746 607 748 609
rect 751 607 753 609
rect 756 607 758 609
rect 761 607 763 609
rect 766 607 768 609
rect 771 607 773 609
rect 776 607 778 609
rect 781 607 783 609
rect 786 607 788 609
rect 791 607 793 609
rect 796 607 798 609
rect 801 607 803 609
rect 806 607 808 609
rect 811 607 813 609
rect 816 607 818 609
rect 821 607 823 609
rect 826 607 828 609
rect 831 607 833 609
rect 836 607 838 609
rect 841 607 843 609
rect 846 607 848 609
rect 851 607 853 609
rect 856 607 858 609
rect 861 607 863 609
rect 866 607 868 609
rect 871 607 873 609
rect 876 607 878 609
rect 881 607 883 609
rect 886 607 888 609
rect 891 607 893 609
rect 896 607 898 609
rect 901 607 903 609
rect 906 607 908 609
rect 911 607 913 609
rect 916 607 918 609
rect 921 607 923 609
rect 926 607 928 609
rect 931 607 933 609
rect 936 607 938 609
rect 941 607 943 609
rect 946 607 948 609
rect 951 607 953 609
rect 956 607 958 609
rect 961 607 963 609
rect 966 607 968 609
rect 971 607 973 609
rect 976 607 978 609
rect 981 607 983 609
rect 986 607 988 609
rect 991 607 993 609
rect 996 607 998 609
rect 331 602 333 604
rect 336 602 338 604
rect 341 602 343 604
rect 346 602 348 604
rect 351 602 353 604
rect 356 602 358 604
rect 361 602 363 604
rect 366 602 368 604
rect 371 602 373 604
rect 376 602 378 604
rect 381 602 383 604
rect 386 602 388 604
rect 391 602 393 604
rect 396 602 398 604
rect 401 602 403 604
rect 406 602 408 604
rect 411 602 413 604
rect 416 602 418 604
rect 421 602 423 604
rect 426 602 428 604
rect 431 602 433 604
rect 436 602 438 604
rect 441 602 443 604
rect 446 602 448 604
rect 451 602 453 604
rect 456 602 458 604
rect 461 602 463 604
rect 466 602 468 604
rect 471 602 473 604
rect 476 602 478 604
rect 481 602 483 604
rect 486 602 488 604
rect 491 602 493 604
rect 496 602 498 604
rect 501 602 503 604
rect 506 602 508 604
rect 511 602 513 604
rect 516 602 518 604
rect 521 602 523 604
rect 526 602 528 604
rect 531 602 533 604
rect 536 602 538 604
rect 541 602 543 604
rect 546 602 548 604
rect 551 602 553 604
rect 556 602 558 604
rect 561 602 563 604
rect 566 602 568 604
rect 571 602 573 604
rect 576 602 578 604
rect 581 602 583 604
rect 586 602 588 604
rect 591 602 593 604
rect 596 602 598 604
rect 601 602 603 604
rect 606 602 608 604
rect 611 602 613 604
rect 616 602 618 604
rect 621 602 623 604
rect 626 602 628 604
rect 631 602 633 604
rect 636 602 638 604
rect 641 602 643 604
rect 646 602 648 604
rect 651 602 653 604
rect 656 602 658 604
rect 661 602 663 604
rect 666 602 668 604
rect 671 602 673 604
rect 676 602 678 604
rect 681 602 683 604
rect 686 602 688 604
rect 691 602 693 604
rect 696 602 698 604
rect 701 602 703 604
rect 706 602 708 604
rect 711 602 713 604
rect 716 602 718 604
rect 721 602 723 604
rect 726 602 728 604
rect 731 602 733 604
rect 736 602 738 604
rect 741 602 743 604
rect 746 602 748 604
rect 751 602 753 604
rect 756 602 758 604
rect 761 602 763 604
rect 766 602 768 604
rect 771 602 773 604
rect 776 602 778 604
rect 781 602 783 604
rect 786 602 788 604
rect 791 602 793 604
rect 796 602 798 604
rect 801 602 803 604
rect 806 602 808 604
rect 811 602 813 604
rect 816 602 818 604
rect 821 602 823 604
rect 826 602 828 604
rect 831 602 833 604
rect 836 602 838 604
rect 841 602 843 604
rect 846 602 848 604
rect 851 602 853 604
rect 856 602 858 604
rect 861 602 863 604
rect 866 602 868 604
rect 871 602 873 604
rect 876 602 878 604
rect 881 602 883 604
rect 886 602 888 604
rect 891 602 893 604
rect 896 602 898 604
rect 901 602 903 604
rect 906 602 908 604
rect 911 602 913 604
rect 916 602 918 604
rect 921 602 923 604
rect 926 602 928 604
rect 931 602 933 604
rect 936 602 938 604
rect 941 602 943 604
rect 946 602 948 604
rect 951 602 953 604
rect 956 602 958 604
rect 961 602 963 604
rect 966 602 968 604
rect 971 602 973 604
rect 976 602 978 604
rect 981 602 983 604
rect 986 602 988 604
rect 991 602 993 604
rect 996 602 998 604
rect 331 597 333 599
rect 336 597 338 599
rect 341 597 343 599
rect 346 597 348 599
rect 351 597 353 599
rect 356 597 358 599
rect 361 597 363 599
rect 366 597 368 599
rect 371 597 373 599
rect 376 597 378 599
rect 381 597 383 599
rect 386 597 388 599
rect 391 597 393 599
rect 396 597 398 599
rect 401 597 403 599
rect 406 597 408 599
rect 411 597 413 599
rect 416 597 418 599
rect 421 597 423 599
rect 426 597 428 599
rect 431 597 433 599
rect 436 597 438 599
rect 441 597 443 599
rect 446 597 448 599
rect 451 597 453 599
rect 456 597 458 599
rect 461 597 463 599
rect 466 597 468 599
rect 471 597 473 599
rect 476 597 478 599
rect 481 597 483 599
rect 486 597 488 599
rect 491 597 493 599
rect 496 597 498 599
rect 501 597 503 599
rect 506 597 508 599
rect 511 597 513 599
rect 516 597 518 599
rect 521 597 523 599
rect 526 597 528 599
rect 531 597 533 599
rect 536 597 538 599
rect 541 597 543 599
rect 546 597 548 599
rect 551 597 553 599
rect 556 597 558 599
rect 561 597 563 599
rect 566 597 568 599
rect 571 597 573 599
rect 576 597 578 599
rect 581 597 583 599
rect 586 597 588 599
rect 591 597 593 599
rect 596 597 598 599
rect 601 597 603 599
rect 606 597 608 599
rect 611 597 613 599
rect 616 597 618 599
rect 621 597 623 599
rect 626 597 628 599
rect 631 597 633 599
rect 636 597 638 599
rect 641 597 643 599
rect 646 597 648 599
rect 651 597 653 599
rect 656 597 658 599
rect 661 597 663 599
rect 666 597 668 599
rect 671 597 673 599
rect 676 597 678 599
rect 681 597 683 599
rect 686 597 688 599
rect 691 597 693 599
rect 696 597 698 599
rect 701 597 703 599
rect 706 597 708 599
rect 711 597 713 599
rect 716 597 718 599
rect 721 597 723 599
rect 726 597 728 599
rect 731 597 733 599
rect 736 597 738 599
rect 741 597 743 599
rect 746 597 748 599
rect 751 597 753 599
rect 756 597 758 599
rect 761 597 763 599
rect 766 597 768 599
rect 771 597 773 599
rect 776 597 778 599
rect 781 597 783 599
rect 786 597 788 599
rect 791 597 793 599
rect 796 597 798 599
rect 801 597 803 599
rect 806 597 808 599
rect 811 597 813 599
rect 816 597 818 599
rect 821 597 823 599
rect 826 597 828 599
rect 831 597 833 599
rect 836 597 838 599
rect 841 597 843 599
rect 846 597 848 599
rect 851 597 853 599
rect 856 597 858 599
rect 861 597 863 599
rect 866 597 868 599
rect 871 597 873 599
rect 876 597 878 599
rect 881 597 883 599
rect 886 597 888 599
rect 891 597 893 599
rect 896 597 898 599
rect 901 597 903 599
rect 906 597 908 599
rect 911 597 913 599
rect 916 597 918 599
rect 921 597 923 599
rect 926 597 928 599
rect 931 597 933 599
rect 936 597 938 599
rect 941 597 943 599
rect 946 597 948 599
rect 951 597 953 599
rect 956 597 958 599
rect 961 597 963 599
rect 966 597 968 599
rect 971 597 973 599
rect 976 597 978 599
rect 981 597 983 599
rect 986 597 988 599
rect 991 597 993 599
rect 996 597 998 599
rect 331 592 333 594
rect 336 592 338 594
rect 341 592 343 594
rect 346 592 348 594
rect 351 592 353 594
rect 356 592 358 594
rect 361 592 363 594
rect 366 592 368 594
rect 371 592 373 594
rect 376 592 378 594
rect 381 592 383 594
rect 386 592 388 594
rect 391 592 393 594
rect 396 592 398 594
rect 401 592 403 594
rect 406 592 408 594
rect 411 592 413 594
rect 416 592 418 594
rect 421 592 423 594
rect 426 592 428 594
rect 431 592 433 594
rect 436 592 438 594
rect 441 592 443 594
rect 446 592 448 594
rect 451 592 453 594
rect 456 592 458 594
rect 461 592 463 594
rect 466 592 468 594
rect 471 592 473 594
rect 476 592 478 594
rect 481 592 483 594
rect 486 592 488 594
rect 491 592 493 594
rect 496 592 498 594
rect 501 592 503 594
rect 506 592 508 594
rect 511 592 513 594
rect 516 592 518 594
rect 521 592 523 594
rect 526 592 528 594
rect 531 592 533 594
rect 536 592 538 594
rect 541 592 543 594
rect 546 592 548 594
rect 551 592 553 594
rect 556 592 558 594
rect 561 592 563 594
rect 566 592 568 594
rect 571 592 573 594
rect 576 592 578 594
rect 581 592 583 594
rect 586 592 588 594
rect 591 592 593 594
rect 596 592 598 594
rect 601 592 603 594
rect 606 592 608 594
rect 611 592 613 594
rect 616 592 618 594
rect 621 592 623 594
rect 626 592 628 594
rect 631 592 633 594
rect 636 592 638 594
rect 641 592 643 594
rect 646 592 648 594
rect 651 592 653 594
rect 656 592 658 594
rect 661 592 663 594
rect 666 592 668 594
rect 671 592 673 594
rect 676 592 678 594
rect 681 592 683 594
rect 686 592 688 594
rect 691 592 693 594
rect 696 592 698 594
rect 701 592 703 594
rect 706 592 708 594
rect 711 592 713 594
rect 716 592 718 594
rect 721 592 723 594
rect 726 592 728 594
rect 731 592 733 594
rect 736 592 738 594
rect 741 592 743 594
rect 746 592 748 594
rect 751 592 753 594
rect 756 592 758 594
rect 761 592 763 594
rect 766 592 768 594
rect 771 592 773 594
rect 776 592 778 594
rect 781 592 783 594
rect 786 592 788 594
rect 791 592 793 594
rect 796 592 798 594
rect 801 592 803 594
rect 806 592 808 594
rect 811 592 813 594
rect 816 592 818 594
rect 821 592 823 594
rect 826 592 828 594
rect 831 592 833 594
rect 836 592 838 594
rect 841 592 843 594
rect 846 592 848 594
rect 851 592 853 594
rect 856 592 858 594
rect 861 592 863 594
rect 866 592 868 594
rect 871 592 873 594
rect 876 592 878 594
rect 881 592 883 594
rect 886 592 888 594
rect 891 592 893 594
rect 896 592 898 594
rect 901 592 903 594
rect 906 592 908 594
rect 911 592 913 594
rect 916 592 918 594
rect 921 592 923 594
rect 926 592 928 594
rect 931 592 933 594
rect 936 592 938 594
rect 941 592 943 594
rect 946 592 948 594
rect 951 592 953 594
rect 956 592 958 594
rect 961 592 963 594
rect 966 592 968 594
rect 971 592 973 594
rect 976 592 978 594
rect 981 592 983 594
rect 986 592 988 594
rect 991 592 993 594
rect 996 592 998 594
rect 331 587 333 589
rect 336 587 338 589
rect 341 587 343 589
rect 346 587 348 589
rect 351 587 353 589
rect 356 587 358 589
rect 361 587 363 589
rect 366 587 368 589
rect 371 587 373 589
rect 376 587 378 589
rect 381 587 383 589
rect 386 587 388 589
rect 391 587 393 589
rect 396 587 398 589
rect 401 587 403 589
rect 406 587 408 589
rect 411 587 413 589
rect 416 587 418 589
rect 421 587 423 589
rect 426 587 428 589
rect 431 587 433 589
rect 436 587 438 589
rect 441 587 443 589
rect 446 587 448 589
rect 451 587 453 589
rect 456 587 458 589
rect 461 587 463 589
rect 466 587 468 589
rect 471 587 473 589
rect 476 587 478 589
rect 481 587 483 589
rect 486 587 488 589
rect 491 587 493 589
rect 496 587 498 589
rect 501 587 503 589
rect 506 587 508 589
rect 511 587 513 589
rect 516 587 518 589
rect 521 587 523 589
rect 526 587 528 589
rect 531 587 533 589
rect 536 587 538 589
rect 541 587 543 589
rect 546 587 548 589
rect 551 587 553 589
rect 556 587 558 589
rect 561 587 563 589
rect 566 587 568 589
rect 571 587 573 589
rect 576 587 578 589
rect 581 587 583 589
rect 586 587 588 589
rect 591 587 593 589
rect 596 587 598 589
rect 601 587 603 589
rect 606 587 608 589
rect 611 587 613 589
rect 616 587 618 589
rect 621 587 623 589
rect 626 587 628 589
rect 631 587 633 589
rect 636 587 638 589
rect 641 587 643 589
rect 646 587 648 589
rect 651 587 653 589
rect 656 587 658 589
rect 661 587 663 589
rect 666 587 668 589
rect 671 587 673 589
rect 676 587 678 589
rect 681 587 683 589
rect 686 587 688 589
rect 691 587 693 589
rect 696 587 698 589
rect 701 587 703 589
rect 706 587 708 589
rect 711 587 713 589
rect 716 587 718 589
rect 721 587 723 589
rect 726 587 728 589
rect 731 587 733 589
rect 736 587 738 589
rect 741 587 743 589
rect 746 587 748 589
rect 751 587 753 589
rect 756 587 758 589
rect 761 587 763 589
rect 766 587 768 589
rect 771 587 773 589
rect 776 587 778 589
rect 781 587 783 589
rect 786 587 788 589
rect 791 587 793 589
rect 796 587 798 589
rect 801 587 803 589
rect 806 587 808 589
rect 811 587 813 589
rect 816 587 818 589
rect 821 587 823 589
rect 826 587 828 589
rect 831 587 833 589
rect 836 587 838 589
rect 841 587 843 589
rect 846 587 848 589
rect 851 587 853 589
rect 856 587 858 589
rect 861 587 863 589
rect 866 587 868 589
rect 871 587 873 589
rect 876 587 878 589
rect 881 587 883 589
rect 886 587 888 589
rect 891 587 893 589
rect 896 587 898 589
rect 901 587 903 589
rect 906 587 908 589
rect 911 587 913 589
rect 916 587 918 589
rect 921 587 923 589
rect 926 587 928 589
rect 931 587 933 589
rect 936 587 938 589
rect 941 587 943 589
rect 946 587 948 589
rect 951 587 953 589
rect 956 587 958 589
rect 961 587 963 589
rect 966 587 968 589
rect 971 587 973 589
rect 976 587 978 589
rect 981 587 983 589
rect 986 587 988 589
rect 991 587 993 589
rect 996 587 998 589
rect 331 582 333 584
rect 336 582 338 584
rect 341 582 343 584
rect 346 582 348 584
rect 351 582 353 584
rect 356 582 358 584
rect 361 582 363 584
rect 366 582 368 584
rect 371 582 373 584
rect 376 582 378 584
rect 381 582 383 584
rect 386 582 388 584
rect 391 582 393 584
rect 396 582 398 584
rect 401 582 403 584
rect 406 582 408 584
rect 411 582 413 584
rect 416 582 418 584
rect 421 582 423 584
rect 426 582 428 584
rect 431 582 433 584
rect 436 582 438 584
rect 441 582 443 584
rect 446 582 448 584
rect 451 582 453 584
rect 456 582 458 584
rect 461 582 463 584
rect 466 582 468 584
rect 471 582 473 584
rect 476 582 478 584
rect 481 582 483 584
rect 486 582 488 584
rect 491 582 493 584
rect 496 582 498 584
rect 501 582 503 584
rect 506 582 508 584
rect 511 582 513 584
rect 516 582 518 584
rect 521 582 523 584
rect 526 582 528 584
rect 531 582 533 584
rect 536 582 538 584
rect 541 582 543 584
rect 546 582 548 584
rect 551 582 553 584
rect 556 582 558 584
rect 561 582 563 584
rect 566 582 568 584
rect 571 582 573 584
rect 576 582 578 584
rect 581 582 583 584
rect 586 582 588 584
rect 591 582 593 584
rect 596 582 598 584
rect 601 582 603 584
rect 606 582 608 584
rect 611 582 613 584
rect 616 582 618 584
rect 621 582 623 584
rect 626 582 628 584
rect 631 582 633 584
rect 636 582 638 584
rect 641 582 643 584
rect 646 582 648 584
rect 651 582 653 584
rect 656 582 658 584
rect 661 582 663 584
rect 666 582 668 584
rect 671 582 673 584
rect 676 582 678 584
rect 681 582 683 584
rect 686 582 688 584
rect 691 582 693 584
rect 696 582 698 584
rect 701 582 703 584
rect 706 582 708 584
rect 711 582 713 584
rect 716 582 718 584
rect 721 582 723 584
rect 726 582 728 584
rect 731 582 733 584
rect 736 582 738 584
rect 741 582 743 584
rect 746 582 748 584
rect 751 582 753 584
rect 756 582 758 584
rect 761 582 763 584
rect 766 582 768 584
rect 771 582 773 584
rect 776 582 778 584
rect 781 582 783 584
rect 786 582 788 584
rect 791 582 793 584
rect 796 582 798 584
rect 801 582 803 584
rect 806 582 808 584
rect 811 582 813 584
rect 816 582 818 584
rect 821 582 823 584
rect 826 582 828 584
rect 831 582 833 584
rect 836 582 838 584
rect 841 582 843 584
rect 846 582 848 584
rect 851 582 853 584
rect 856 582 858 584
rect 861 582 863 584
rect 866 582 868 584
rect 871 582 873 584
rect 876 582 878 584
rect 881 582 883 584
rect 886 582 888 584
rect 891 582 893 584
rect 896 582 898 584
rect 901 582 903 584
rect 906 582 908 584
rect 911 582 913 584
rect 916 582 918 584
rect 921 582 923 584
rect 926 582 928 584
rect 931 582 933 584
rect 936 582 938 584
rect 941 582 943 584
rect 946 582 948 584
rect 951 582 953 584
rect 956 582 958 584
rect 961 582 963 584
rect 966 582 968 584
rect 971 582 973 584
rect 976 582 978 584
rect 981 582 983 584
rect 986 582 988 584
rect 991 582 993 584
rect 996 582 998 584
rect 331 577 333 579
rect 336 577 338 579
rect 341 577 343 579
rect 346 577 348 579
rect 351 577 353 579
rect 356 577 358 579
rect 361 577 363 579
rect 366 577 368 579
rect 371 577 373 579
rect 376 577 378 579
rect 381 577 383 579
rect 386 577 388 579
rect 391 577 393 579
rect 396 577 398 579
rect 401 577 403 579
rect 406 577 408 579
rect 411 577 413 579
rect 416 577 418 579
rect 421 577 423 579
rect 426 577 428 579
rect 431 577 433 579
rect 436 577 438 579
rect 441 577 443 579
rect 446 577 448 579
rect 451 577 453 579
rect 456 577 458 579
rect 461 577 463 579
rect 466 577 468 579
rect 471 577 473 579
rect 476 577 478 579
rect 481 577 483 579
rect 486 577 488 579
rect 491 577 493 579
rect 496 577 498 579
rect 501 577 503 579
rect 506 577 508 579
rect 511 577 513 579
rect 516 577 518 579
rect 521 577 523 579
rect 526 577 528 579
rect 531 577 533 579
rect 536 577 538 579
rect 541 577 543 579
rect 546 577 548 579
rect 551 577 553 579
rect 556 577 558 579
rect 561 577 563 579
rect 566 577 568 579
rect 571 577 573 579
rect 576 577 578 579
rect 581 577 583 579
rect 586 577 588 579
rect 591 577 593 579
rect 596 577 598 579
rect 601 577 603 579
rect 606 577 608 579
rect 611 577 613 579
rect 616 577 618 579
rect 621 577 623 579
rect 626 577 628 579
rect 631 577 633 579
rect 636 577 638 579
rect 641 577 643 579
rect 646 577 648 579
rect 651 577 653 579
rect 656 577 658 579
rect 661 577 663 579
rect 666 577 668 579
rect 671 577 673 579
rect 676 577 678 579
rect 681 577 683 579
rect 686 577 688 579
rect 691 577 693 579
rect 696 577 698 579
rect 701 577 703 579
rect 706 577 708 579
rect 711 577 713 579
rect 716 577 718 579
rect 721 577 723 579
rect 726 577 728 579
rect 731 577 733 579
rect 736 577 738 579
rect 741 577 743 579
rect 746 577 748 579
rect 751 577 753 579
rect 756 577 758 579
rect 761 577 763 579
rect 766 577 768 579
rect 771 577 773 579
rect 776 577 778 579
rect 781 577 783 579
rect 786 577 788 579
rect 791 577 793 579
rect 796 577 798 579
rect 801 577 803 579
rect 806 577 808 579
rect 811 577 813 579
rect 816 577 818 579
rect 821 577 823 579
rect 826 577 828 579
rect 831 577 833 579
rect 836 577 838 579
rect 841 577 843 579
rect 846 577 848 579
rect 851 577 853 579
rect 856 577 858 579
rect 861 577 863 579
rect 866 577 868 579
rect 871 577 873 579
rect 876 577 878 579
rect 881 577 883 579
rect 886 577 888 579
rect 891 577 893 579
rect 896 577 898 579
rect 901 577 903 579
rect 906 577 908 579
rect 911 577 913 579
rect 916 577 918 579
rect 921 577 923 579
rect 926 577 928 579
rect 931 577 933 579
rect 936 577 938 579
rect 941 577 943 579
rect 946 577 948 579
rect 951 577 953 579
rect 956 577 958 579
rect 961 577 963 579
rect 966 577 968 579
rect 971 577 973 579
rect 976 577 978 579
rect 981 577 983 579
rect 986 577 988 579
rect 991 577 993 579
rect 996 577 998 579
rect 331 572 333 574
rect 336 572 338 574
rect 341 572 343 574
rect 346 572 348 574
rect 351 572 353 574
rect 356 572 358 574
rect 361 572 363 574
rect 366 572 368 574
rect 371 572 373 574
rect 376 572 378 574
rect 381 572 383 574
rect 386 572 388 574
rect 391 572 393 574
rect 396 572 398 574
rect 401 572 403 574
rect 406 572 408 574
rect 411 572 413 574
rect 416 572 418 574
rect 421 572 423 574
rect 426 572 428 574
rect 431 572 433 574
rect 436 572 438 574
rect 441 572 443 574
rect 446 572 448 574
rect 451 572 453 574
rect 456 572 458 574
rect 461 572 463 574
rect 466 572 468 574
rect 471 572 473 574
rect 476 572 478 574
rect 481 572 483 574
rect 486 572 488 574
rect 491 572 493 574
rect 496 572 498 574
rect 501 572 503 574
rect 506 572 508 574
rect 511 572 513 574
rect 516 572 518 574
rect 521 572 523 574
rect 526 572 528 574
rect 531 572 533 574
rect 536 572 538 574
rect 541 572 543 574
rect 546 572 548 574
rect 551 572 553 574
rect 556 572 558 574
rect 561 572 563 574
rect 566 572 568 574
rect 571 572 573 574
rect 576 572 578 574
rect 581 572 583 574
rect 586 572 588 574
rect 591 572 593 574
rect 596 572 598 574
rect 601 572 603 574
rect 606 572 608 574
rect 611 572 613 574
rect 616 572 618 574
rect 621 572 623 574
rect 626 572 628 574
rect 631 572 633 574
rect 636 572 638 574
rect 641 572 643 574
rect 646 572 648 574
rect 651 572 653 574
rect 656 572 658 574
rect 661 572 663 574
rect 666 572 668 574
rect 671 572 673 574
rect 676 572 678 574
rect 681 572 683 574
rect 686 572 688 574
rect 691 572 693 574
rect 696 572 698 574
rect 701 572 703 574
rect 706 572 708 574
rect 711 572 713 574
rect 716 572 718 574
rect 721 572 723 574
rect 726 572 728 574
rect 731 572 733 574
rect 736 572 738 574
rect 741 572 743 574
rect 746 572 748 574
rect 751 572 753 574
rect 756 572 758 574
rect 761 572 763 574
rect 766 572 768 574
rect 771 572 773 574
rect 776 572 778 574
rect 781 572 783 574
rect 786 572 788 574
rect 791 572 793 574
rect 796 572 798 574
rect 801 572 803 574
rect 806 572 808 574
rect 811 572 813 574
rect 816 572 818 574
rect 821 572 823 574
rect 826 572 828 574
rect 831 572 833 574
rect 836 572 838 574
rect 841 572 843 574
rect 846 572 848 574
rect 851 572 853 574
rect 856 572 858 574
rect 861 572 863 574
rect 866 572 868 574
rect 871 572 873 574
rect 876 572 878 574
rect 881 572 883 574
rect 886 572 888 574
rect 891 572 893 574
rect 896 572 898 574
rect 901 572 903 574
rect 906 572 908 574
rect 911 572 913 574
rect 916 572 918 574
rect 921 572 923 574
rect 926 572 928 574
rect 931 572 933 574
rect 936 572 938 574
rect 941 572 943 574
rect 946 572 948 574
rect 951 572 953 574
rect 956 572 958 574
rect 961 572 963 574
rect 966 572 968 574
rect 971 572 973 574
rect 976 572 978 574
rect 981 572 983 574
rect 986 572 988 574
rect 991 572 993 574
rect 996 572 998 574
rect 331 567 333 569
rect 336 567 338 569
rect 341 567 343 569
rect 346 567 348 569
rect 351 567 353 569
rect 356 567 358 569
rect 361 567 363 569
rect 366 567 368 569
rect 371 567 373 569
rect 376 567 378 569
rect 381 567 383 569
rect 386 567 388 569
rect 391 567 393 569
rect 396 567 398 569
rect 401 567 403 569
rect 406 567 408 569
rect 411 567 413 569
rect 416 567 418 569
rect 421 567 423 569
rect 426 567 428 569
rect 431 567 433 569
rect 436 567 438 569
rect 441 567 443 569
rect 446 567 448 569
rect 451 567 453 569
rect 456 567 458 569
rect 461 567 463 569
rect 466 567 468 569
rect 471 567 473 569
rect 476 567 478 569
rect 481 567 483 569
rect 486 567 488 569
rect 491 567 493 569
rect 496 567 498 569
rect 501 567 503 569
rect 506 567 508 569
rect 511 567 513 569
rect 516 567 518 569
rect 521 567 523 569
rect 526 567 528 569
rect 531 567 533 569
rect 536 567 538 569
rect 541 567 543 569
rect 546 567 548 569
rect 551 567 553 569
rect 556 567 558 569
rect 561 567 563 569
rect 566 567 568 569
rect 571 567 573 569
rect 576 567 578 569
rect 581 567 583 569
rect 586 567 588 569
rect 591 567 593 569
rect 596 567 598 569
rect 601 567 603 569
rect 606 567 608 569
rect 611 567 613 569
rect 616 567 618 569
rect 621 567 623 569
rect 626 567 628 569
rect 631 567 633 569
rect 636 567 638 569
rect 641 567 643 569
rect 646 567 648 569
rect 651 567 653 569
rect 656 567 658 569
rect 661 567 663 569
rect 666 567 668 569
rect 671 567 673 569
rect 676 567 678 569
rect 681 567 683 569
rect 686 567 688 569
rect 691 567 693 569
rect 696 567 698 569
rect 701 567 703 569
rect 706 567 708 569
rect 711 567 713 569
rect 716 567 718 569
rect 721 567 723 569
rect 726 567 728 569
rect 731 567 733 569
rect 736 567 738 569
rect 741 567 743 569
rect 746 567 748 569
rect 751 567 753 569
rect 756 567 758 569
rect 761 567 763 569
rect 766 567 768 569
rect 771 567 773 569
rect 776 567 778 569
rect 781 567 783 569
rect 786 567 788 569
rect 791 567 793 569
rect 796 567 798 569
rect 801 567 803 569
rect 806 567 808 569
rect 811 567 813 569
rect 816 567 818 569
rect 821 567 823 569
rect 826 567 828 569
rect 831 567 833 569
rect 836 567 838 569
rect 841 567 843 569
rect 846 567 848 569
rect 851 567 853 569
rect 856 567 858 569
rect 861 567 863 569
rect 866 567 868 569
rect 871 567 873 569
rect 876 567 878 569
rect 881 567 883 569
rect 886 567 888 569
rect 891 567 893 569
rect 896 567 898 569
rect 901 567 903 569
rect 906 567 908 569
rect 911 567 913 569
rect 916 567 918 569
rect 921 567 923 569
rect 926 567 928 569
rect 931 567 933 569
rect 936 567 938 569
rect 941 567 943 569
rect 946 567 948 569
rect 951 567 953 569
rect 956 567 958 569
rect 961 567 963 569
rect 966 567 968 569
rect 971 567 973 569
rect 976 567 978 569
rect 981 567 983 569
rect 986 567 988 569
rect 991 567 993 569
rect 996 567 998 569
rect 331 562 333 564
rect 336 562 338 564
rect 341 562 343 564
rect 346 562 348 564
rect 351 562 353 564
rect 356 562 358 564
rect 361 562 363 564
rect 366 562 368 564
rect 371 562 373 564
rect 376 562 378 564
rect 381 562 383 564
rect 386 562 388 564
rect 391 562 393 564
rect 396 562 398 564
rect 401 562 403 564
rect 406 562 408 564
rect 411 562 413 564
rect 416 562 418 564
rect 421 562 423 564
rect 426 562 428 564
rect 431 562 433 564
rect 436 562 438 564
rect 441 562 443 564
rect 446 562 448 564
rect 451 562 453 564
rect 456 562 458 564
rect 461 562 463 564
rect 466 562 468 564
rect 471 562 473 564
rect 476 562 478 564
rect 481 562 483 564
rect 486 562 488 564
rect 491 562 493 564
rect 496 562 498 564
rect 501 562 503 564
rect 506 562 508 564
rect 511 562 513 564
rect 516 562 518 564
rect 521 562 523 564
rect 526 562 528 564
rect 531 562 533 564
rect 536 562 538 564
rect 541 562 543 564
rect 546 562 548 564
rect 551 562 553 564
rect 556 562 558 564
rect 561 562 563 564
rect 566 562 568 564
rect 571 562 573 564
rect 576 562 578 564
rect 581 562 583 564
rect 586 562 588 564
rect 591 562 593 564
rect 596 562 598 564
rect 601 562 603 564
rect 606 562 608 564
rect 611 562 613 564
rect 616 562 618 564
rect 621 562 623 564
rect 626 562 628 564
rect 631 562 633 564
rect 636 562 638 564
rect 641 562 643 564
rect 646 562 648 564
rect 651 562 653 564
rect 656 562 658 564
rect 661 562 663 564
rect 666 562 668 564
rect 671 562 673 564
rect 676 562 678 564
rect 681 562 683 564
rect 686 562 688 564
rect 691 562 693 564
rect 696 562 698 564
rect 701 562 703 564
rect 706 562 708 564
rect 711 562 713 564
rect 716 562 718 564
rect 721 562 723 564
rect 726 562 728 564
rect 731 562 733 564
rect 736 562 738 564
rect 741 562 743 564
rect 746 562 748 564
rect 751 562 753 564
rect 756 562 758 564
rect 761 562 763 564
rect 766 562 768 564
rect 771 562 773 564
rect 776 562 778 564
rect 781 562 783 564
rect 786 562 788 564
rect 791 562 793 564
rect 796 562 798 564
rect 801 562 803 564
rect 806 562 808 564
rect 811 562 813 564
rect 816 562 818 564
rect 821 562 823 564
rect 826 562 828 564
rect 831 562 833 564
rect 836 562 838 564
rect 841 562 843 564
rect 846 562 848 564
rect 851 562 853 564
rect 856 562 858 564
rect 861 562 863 564
rect 866 562 868 564
rect 871 562 873 564
rect 876 562 878 564
rect 881 562 883 564
rect 886 562 888 564
rect 891 562 893 564
rect 896 562 898 564
rect 901 562 903 564
rect 906 562 908 564
rect 911 562 913 564
rect 916 562 918 564
rect 921 562 923 564
rect 926 562 928 564
rect 931 562 933 564
rect 936 562 938 564
rect 941 562 943 564
rect 946 562 948 564
rect 951 562 953 564
rect 956 562 958 564
rect 961 562 963 564
rect 966 562 968 564
rect 971 562 973 564
rect 976 562 978 564
rect 981 562 983 564
rect 986 562 988 564
rect 991 562 993 564
rect 996 562 998 564
rect 331 557 333 559
rect 336 557 338 559
rect 341 557 343 559
rect 346 557 348 559
rect 351 557 353 559
rect 356 557 358 559
rect 361 557 363 559
rect 366 557 368 559
rect 371 557 373 559
rect 376 557 378 559
rect 381 557 383 559
rect 386 557 388 559
rect 391 557 393 559
rect 396 557 398 559
rect 401 557 403 559
rect 406 557 408 559
rect 411 557 413 559
rect 416 557 418 559
rect 421 557 423 559
rect 426 557 428 559
rect 431 557 433 559
rect 436 557 438 559
rect 441 557 443 559
rect 446 557 448 559
rect 451 557 453 559
rect 456 557 458 559
rect 461 557 463 559
rect 466 557 468 559
rect 471 557 473 559
rect 476 557 478 559
rect 481 557 483 559
rect 486 557 488 559
rect 491 557 493 559
rect 496 557 498 559
rect 501 557 503 559
rect 506 557 508 559
rect 511 557 513 559
rect 516 557 518 559
rect 521 557 523 559
rect 526 557 528 559
rect 531 557 533 559
rect 536 557 538 559
rect 541 557 543 559
rect 546 557 548 559
rect 551 557 553 559
rect 556 557 558 559
rect 561 557 563 559
rect 566 557 568 559
rect 571 557 573 559
rect 576 557 578 559
rect 581 557 583 559
rect 586 557 588 559
rect 591 557 593 559
rect 596 557 598 559
rect 601 557 603 559
rect 606 557 608 559
rect 611 557 613 559
rect 616 557 618 559
rect 621 557 623 559
rect 626 557 628 559
rect 631 557 633 559
rect 636 557 638 559
rect 641 557 643 559
rect 646 557 648 559
rect 651 557 653 559
rect 656 557 658 559
rect 661 557 663 559
rect 666 557 668 559
rect 671 557 673 559
rect 676 557 678 559
rect 681 557 683 559
rect 686 557 688 559
rect 691 557 693 559
rect 696 557 698 559
rect 701 557 703 559
rect 706 557 708 559
rect 711 557 713 559
rect 716 557 718 559
rect 721 557 723 559
rect 726 557 728 559
rect 731 557 733 559
rect 736 557 738 559
rect 741 557 743 559
rect 746 557 748 559
rect 751 557 753 559
rect 756 557 758 559
rect 761 557 763 559
rect 766 557 768 559
rect 771 557 773 559
rect 776 557 778 559
rect 781 557 783 559
rect 786 557 788 559
rect 791 557 793 559
rect 796 557 798 559
rect 801 557 803 559
rect 806 557 808 559
rect 811 557 813 559
rect 816 557 818 559
rect 821 557 823 559
rect 826 557 828 559
rect 831 557 833 559
rect 836 557 838 559
rect 841 557 843 559
rect 846 557 848 559
rect 851 557 853 559
rect 856 557 858 559
rect 861 557 863 559
rect 866 557 868 559
rect 871 557 873 559
rect 876 557 878 559
rect 881 557 883 559
rect 886 557 888 559
rect 891 557 893 559
rect 896 557 898 559
rect 901 557 903 559
rect 906 557 908 559
rect 911 557 913 559
rect 916 557 918 559
rect 921 557 923 559
rect 926 557 928 559
rect 931 557 933 559
rect 936 557 938 559
rect 941 557 943 559
rect 946 557 948 559
rect 951 557 953 559
rect 956 557 958 559
rect 961 557 963 559
rect 966 557 968 559
rect 971 557 973 559
rect 976 557 978 559
rect 981 557 983 559
rect 986 557 988 559
rect 991 557 993 559
rect 996 557 998 559
rect 331 552 333 554
rect 336 552 338 554
rect 341 552 343 554
rect 346 552 348 554
rect 351 552 353 554
rect 356 552 358 554
rect 361 552 363 554
rect 366 552 368 554
rect 371 552 373 554
rect 376 552 378 554
rect 381 552 383 554
rect 386 552 388 554
rect 391 552 393 554
rect 396 552 398 554
rect 401 552 403 554
rect 406 552 408 554
rect 411 552 413 554
rect 416 552 418 554
rect 421 552 423 554
rect 426 552 428 554
rect 431 552 433 554
rect 436 552 438 554
rect 441 552 443 554
rect 446 552 448 554
rect 451 552 453 554
rect 456 552 458 554
rect 461 552 463 554
rect 466 552 468 554
rect 471 552 473 554
rect 476 552 478 554
rect 481 552 483 554
rect 486 552 488 554
rect 491 552 493 554
rect 496 552 498 554
rect 501 552 503 554
rect 506 552 508 554
rect 511 552 513 554
rect 516 552 518 554
rect 521 552 523 554
rect 526 552 528 554
rect 531 552 533 554
rect 536 552 538 554
rect 541 552 543 554
rect 546 552 548 554
rect 551 552 553 554
rect 556 552 558 554
rect 561 552 563 554
rect 566 552 568 554
rect 571 552 573 554
rect 576 552 578 554
rect 581 552 583 554
rect 586 552 588 554
rect 591 552 593 554
rect 596 552 598 554
rect 601 552 603 554
rect 606 552 608 554
rect 611 552 613 554
rect 616 552 618 554
rect 621 552 623 554
rect 626 552 628 554
rect 631 552 633 554
rect 636 552 638 554
rect 641 552 643 554
rect 646 552 648 554
rect 651 552 653 554
rect 656 552 658 554
rect 661 552 663 554
rect 666 552 668 554
rect 671 552 673 554
rect 676 552 678 554
rect 681 552 683 554
rect 686 552 688 554
rect 691 552 693 554
rect 696 552 698 554
rect 701 552 703 554
rect 706 552 708 554
rect 711 552 713 554
rect 716 552 718 554
rect 721 552 723 554
rect 726 552 728 554
rect 731 552 733 554
rect 736 552 738 554
rect 741 552 743 554
rect 746 552 748 554
rect 751 552 753 554
rect 756 552 758 554
rect 761 552 763 554
rect 766 552 768 554
rect 771 552 773 554
rect 776 552 778 554
rect 781 552 783 554
rect 786 552 788 554
rect 791 552 793 554
rect 796 552 798 554
rect 801 552 803 554
rect 806 552 808 554
rect 811 552 813 554
rect 816 552 818 554
rect 821 552 823 554
rect 826 552 828 554
rect 831 552 833 554
rect 836 552 838 554
rect 841 552 843 554
rect 846 552 848 554
rect 851 552 853 554
rect 856 552 858 554
rect 861 552 863 554
rect 866 552 868 554
rect 871 552 873 554
rect 876 552 878 554
rect 881 552 883 554
rect 886 552 888 554
rect 891 552 893 554
rect 896 552 898 554
rect 901 552 903 554
rect 906 552 908 554
rect 911 552 913 554
rect 916 552 918 554
rect 921 552 923 554
rect 926 552 928 554
rect 931 552 933 554
rect 936 552 938 554
rect 941 552 943 554
rect 946 552 948 554
rect 951 552 953 554
rect 956 552 958 554
rect 961 552 963 554
rect 966 552 968 554
rect 971 552 973 554
rect 976 552 978 554
rect 981 552 983 554
rect 986 552 988 554
rect 991 552 993 554
rect 996 552 998 554
rect 331 547 333 549
rect 336 547 338 549
rect 341 547 343 549
rect 346 547 348 549
rect 351 547 353 549
rect 356 547 358 549
rect 361 547 363 549
rect 366 547 368 549
rect 371 547 373 549
rect 376 547 378 549
rect 381 547 383 549
rect 386 547 388 549
rect 391 547 393 549
rect 396 547 398 549
rect 401 547 403 549
rect 406 547 408 549
rect 411 547 413 549
rect 416 547 418 549
rect 421 547 423 549
rect 426 547 428 549
rect 431 547 433 549
rect 436 547 438 549
rect 441 547 443 549
rect 446 547 448 549
rect 451 547 453 549
rect 456 547 458 549
rect 461 547 463 549
rect 466 547 468 549
rect 471 547 473 549
rect 476 547 478 549
rect 481 547 483 549
rect 486 547 488 549
rect 491 547 493 549
rect 496 547 498 549
rect 501 547 503 549
rect 506 547 508 549
rect 511 547 513 549
rect 516 547 518 549
rect 521 547 523 549
rect 526 547 528 549
rect 531 547 533 549
rect 536 547 538 549
rect 541 547 543 549
rect 546 547 548 549
rect 551 547 553 549
rect 556 547 558 549
rect 561 547 563 549
rect 566 547 568 549
rect 571 547 573 549
rect 576 547 578 549
rect 581 547 583 549
rect 586 547 588 549
rect 591 547 593 549
rect 596 547 598 549
rect 601 547 603 549
rect 606 547 608 549
rect 611 547 613 549
rect 616 547 618 549
rect 621 547 623 549
rect 626 547 628 549
rect 631 547 633 549
rect 636 547 638 549
rect 641 547 643 549
rect 646 547 648 549
rect 651 547 653 549
rect 656 547 658 549
rect 661 547 663 549
rect 666 547 668 549
rect 671 547 673 549
rect 676 547 678 549
rect 681 547 683 549
rect 686 547 688 549
rect 691 547 693 549
rect 696 547 698 549
rect 701 547 703 549
rect 706 547 708 549
rect 711 547 713 549
rect 716 547 718 549
rect 721 547 723 549
rect 726 547 728 549
rect 731 547 733 549
rect 736 547 738 549
rect 741 547 743 549
rect 746 547 748 549
rect 751 547 753 549
rect 756 547 758 549
rect 761 547 763 549
rect 766 547 768 549
rect 771 547 773 549
rect 776 547 778 549
rect 781 547 783 549
rect 786 547 788 549
rect 791 547 793 549
rect 796 547 798 549
rect 801 547 803 549
rect 806 547 808 549
rect 811 547 813 549
rect 816 547 818 549
rect 821 547 823 549
rect 826 547 828 549
rect 831 547 833 549
rect 836 547 838 549
rect 841 547 843 549
rect 846 547 848 549
rect 851 547 853 549
rect 856 547 858 549
rect 861 547 863 549
rect 866 547 868 549
rect 871 547 873 549
rect 876 547 878 549
rect 881 547 883 549
rect 886 547 888 549
rect 891 547 893 549
rect 896 547 898 549
rect 901 547 903 549
rect 906 547 908 549
rect 911 547 913 549
rect 916 547 918 549
rect 921 547 923 549
rect 926 547 928 549
rect 931 547 933 549
rect 936 547 938 549
rect 941 547 943 549
rect 946 547 948 549
rect 951 547 953 549
rect 956 547 958 549
rect 961 547 963 549
rect 966 547 968 549
rect 971 547 973 549
rect 976 547 978 549
rect 981 547 983 549
rect 986 547 988 549
rect 991 547 993 549
rect 996 547 998 549
rect 331 542 333 544
rect 336 542 338 544
rect 341 542 343 544
rect 346 542 348 544
rect 351 542 353 544
rect 356 542 358 544
rect 361 542 363 544
rect 366 542 368 544
rect 371 542 373 544
rect 376 542 378 544
rect 381 542 383 544
rect 386 542 388 544
rect 391 542 393 544
rect 396 542 398 544
rect 401 542 403 544
rect 406 542 408 544
rect 411 542 413 544
rect 416 542 418 544
rect 421 542 423 544
rect 426 542 428 544
rect 431 542 433 544
rect 436 542 438 544
rect 441 542 443 544
rect 446 542 448 544
rect 451 542 453 544
rect 456 542 458 544
rect 461 542 463 544
rect 466 542 468 544
rect 471 542 473 544
rect 476 542 478 544
rect 481 542 483 544
rect 486 542 488 544
rect 491 542 493 544
rect 496 542 498 544
rect 501 542 503 544
rect 506 542 508 544
rect 511 542 513 544
rect 516 542 518 544
rect 521 542 523 544
rect 526 542 528 544
rect 531 542 533 544
rect 536 542 538 544
rect 541 542 543 544
rect 546 542 548 544
rect 551 542 553 544
rect 556 542 558 544
rect 561 542 563 544
rect 566 542 568 544
rect 571 542 573 544
rect 576 542 578 544
rect 581 542 583 544
rect 586 542 588 544
rect 591 542 593 544
rect 596 542 598 544
rect 601 542 603 544
rect 606 542 608 544
rect 611 542 613 544
rect 616 542 618 544
rect 621 542 623 544
rect 626 542 628 544
rect 631 542 633 544
rect 636 542 638 544
rect 641 542 643 544
rect 646 542 648 544
rect 651 542 653 544
rect 656 542 658 544
rect 661 542 663 544
rect 666 542 668 544
rect 671 542 673 544
rect 676 542 678 544
rect 681 542 683 544
rect 686 542 688 544
rect 691 542 693 544
rect 696 542 698 544
rect 701 542 703 544
rect 706 542 708 544
rect 711 542 713 544
rect 716 542 718 544
rect 721 542 723 544
rect 726 542 728 544
rect 731 542 733 544
rect 736 542 738 544
rect 741 542 743 544
rect 746 542 748 544
rect 751 542 753 544
rect 756 542 758 544
rect 761 542 763 544
rect 766 542 768 544
rect 771 542 773 544
rect 776 542 778 544
rect 781 542 783 544
rect 786 542 788 544
rect 791 542 793 544
rect 796 542 798 544
rect 801 542 803 544
rect 806 542 808 544
rect 811 542 813 544
rect 816 542 818 544
rect 821 542 823 544
rect 826 542 828 544
rect 831 542 833 544
rect 836 542 838 544
rect 841 542 843 544
rect 846 542 848 544
rect 851 542 853 544
rect 856 542 858 544
rect 861 542 863 544
rect 866 542 868 544
rect 871 542 873 544
rect 876 542 878 544
rect 881 542 883 544
rect 886 542 888 544
rect 891 542 893 544
rect 896 542 898 544
rect 901 542 903 544
rect 906 542 908 544
rect 911 542 913 544
rect 916 542 918 544
rect 921 542 923 544
rect 926 542 928 544
rect 931 542 933 544
rect 936 542 938 544
rect 941 542 943 544
rect 946 542 948 544
rect 951 542 953 544
rect 956 542 958 544
rect 961 542 963 544
rect 966 542 968 544
rect 971 542 973 544
rect 976 542 978 544
rect 981 542 983 544
rect 986 542 988 544
rect 991 542 993 544
rect 996 542 998 544
rect 331 537 333 539
rect 336 537 338 539
rect 341 537 343 539
rect 346 537 348 539
rect 351 537 353 539
rect 356 537 358 539
rect 361 537 363 539
rect 366 537 368 539
rect 371 537 373 539
rect 376 537 378 539
rect 381 537 383 539
rect 386 537 388 539
rect 391 537 393 539
rect 396 537 398 539
rect 401 537 403 539
rect 406 537 408 539
rect 411 537 413 539
rect 416 537 418 539
rect 421 537 423 539
rect 426 537 428 539
rect 431 537 433 539
rect 436 537 438 539
rect 441 537 443 539
rect 446 537 448 539
rect 451 537 453 539
rect 456 537 458 539
rect 461 537 463 539
rect 466 537 468 539
rect 471 537 473 539
rect 476 537 478 539
rect 481 537 483 539
rect 486 537 488 539
rect 491 537 493 539
rect 496 537 498 539
rect 501 537 503 539
rect 506 537 508 539
rect 511 537 513 539
rect 516 537 518 539
rect 521 537 523 539
rect 526 537 528 539
rect 531 537 533 539
rect 536 537 538 539
rect 541 537 543 539
rect 546 537 548 539
rect 551 537 553 539
rect 556 537 558 539
rect 561 537 563 539
rect 566 537 568 539
rect 571 537 573 539
rect 576 537 578 539
rect 581 537 583 539
rect 586 537 588 539
rect 591 537 593 539
rect 596 537 598 539
rect 601 537 603 539
rect 606 537 608 539
rect 611 537 613 539
rect 616 537 618 539
rect 621 537 623 539
rect 626 537 628 539
rect 631 537 633 539
rect 636 537 638 539
rect 641 537 643 539
rect 646 537 648 539
rect 651 537 653 539
rect 656 537 658 539
rect 661 537 663 539
rect 666 537 668 539
rect 671 537 673 539
rect 676 537 678 539
rect 681 537 683 539
rect 686 537 688 539
rect 691 537 693 539
rect 696 537 698 539
rect 701 537 703 539
rect 706 537 708 539
rect 711 537 713 539
rect 716 537 718 539
rect 721 537 723 539
rect 726 537 728 539
rect 731 537 733 539
rect 736 537 738 539
rect 741 537 743 539
rect 746 537 748 539
rect 751 537 753 539
rect 756 537 758 539
rect 761 537 763 539
rect 766 537 768 539
rect 771 537 773 539
rect 776 537 778 539
rect 781 537 783 539
rect 786 537 788 539
rect 791 537 793 539
rect 796 537 798 539
rect 801 537 803 539
rect 806 537 808 539
rect 811 537 813 539
rect 816 537 818 539
rect 821 537 823 539
rect 826 537 828 539
rect 831 537 833 539
rect 836 537 838 539
rect 841 537 843 539
rect 846 537 848 539
rect 851 537 853 539
rect 856 537 858 539
rect 861 537 863 539
rect 866 537 868 539
rect 871 537 873 539
rect 876 537 878 539
rect 881 537 883 539
rect 886 537 888 539
rect 891 537 893 539
rect 896 537 898 539
rect 901 537 903 539
rect 906 537 908 539
rect 911 537 913 539
rect 916 537 918 539
rect 921 537 923 539
rect 926 537 928 539
rect 931 537 933 539
rect 936 537 938 539
rect 941 537 943 539
rect 946 537 948 539
rect 951 537 953 539
rect 956 537 958 539
rect 961 537 963 539
rect 966 537 968 539
rect 971 537 973 539
rect 976 537 978 539
rect 981 537 983 539
rect 986 537 988 539
rect 991 537 993 539
rect 996 537 998 539
rect 331 532 333 534
rect 336 532 338 534
rect 341 532 343 534
rect 346 532 348 534
rect 351 532 353 534
rect 356 532 358 534
rect 361 532 363 534
rect 366 532 368 534
rect 371 532 373 534
rect 376 532 378 534
rect 381 532 383 534
rect 386 532 388 534
rect 391 532 393 534
rect 396 532 398 534
rect 401 532 403 534
rect 406 532 408 534
rect 411 532 413 534
rect 416 532 418 534
rect 421 532 423 534
rect 426 532 428 534
rect 431 532 433 534
rect 436 532 438 534
rect 441 532 443 534
rect 446 532 448 534
rect 451 532 453 534
rect 456 532 458 534
rect 461 532 463 534
rect 466 532 468 534
rect 471 532 473 534
rect 476 532 478 534
rect 481 532 483 534
rect 486 532 488 534
rect 491 532 493 534
rect 496 532 498 534
rect 501 532 503 534
rect 506 532 508 534
rect 511 532 513 534
rect 516 532 518 534
rect 521 532 523 534
rect 526 532 528 534
rect 531 532 533 534
rect 536 532 538 534
rect 541 532 543 534
rect 546 532 548 534
rect 551 532 553 534
rect 556 532 558 534
rect 561 532 563 534
rect 566 532 568 534
rect 571 532 573 534
rect 576 532 578 534
rect 581 532 583 534
rect 586 532 588 534
rect 591 532 593 534
rect 596 532 598 534
rect 601 532 603 534
rect 606 532 608 534
rect 611 532 613 534
rect 616 532 618 534
rect 621 532 623 534
rect 626 532 628 534
rect 631 532 633 534
rect 636 532 638 534
rect 641 532 643 534
rect 646 532 648 534
rect 651 532 653 534
rect 656 532 658 534
rect 661 532 663 534
rect 666 532 668 534
rect 671 532 673 534
rect 676 532 678 534
rect 681 532 683 534
rect 686 532 688 534
rect 691 532 693 534
rect 696 532 698 534
rect 701 532 703 534
rect 706 532 708 534
rect 711 532 713 534
rect 716 532 718 534
rect 721 532 723 534
rect 726 532 728 534
rect 731 532 733 534
rect 736 532 738 534
rect 741 532 743 534
rect 746 532 748 534
rect 751 532 753 534
rect 756 532 758 534
rect 761 532 763 534
rect 766 532 768 534
rect 771 532 773 534
rect 776 532 778 534
rect 781 532 783 534
rect 786 532 788 534
rect 791 532 793 534
rect 796 532 798 534
rect 801 532 803 534
rect 806 532 808 534
rect 811 532 813 534
rect 816 532 818 534
rect 821 532 823 534
rect 826 532 828 534
rect 831 532 833 534
rect 836 532 838 534
rect 841 532 843 534
rect 846 532 848 534
rect 851 532 853 534
rect 856 532 858 534
rect 861 532 863 534
rect 866 532 868 534
rect 871 532 873 534
rect 876 532 878 534
rect 881 532 883 534
rect 886 532 888 534
rect 891 532 893 534
rect 896 532 898 534
rect 901 532 903 534
rect 906 532 908 534
rect 911 532 913 534
rect 916 532 918 534
rect 921 532 923 534
rect 926 532 928 534
rect 931 532 933 534
rect 936 532 938 534
rect 941 532 943 534
rect 946 532 948 534
rect 951 532 953 534
rect 956 532 958 534
rect 961 532 963 534
rect 966 532 968 534
rect 971 532 973 534
rect 976 532 978 534
rect 981 532 983 534
rect 986 532 988 534
rect 991 532 993 534
rect 996 532 998 534
rect 331 527 333 529
rect 336 527 338 529
rect 341 527 343 529
rect 346 527 348 529
rect 351 527 353 529
rect 356 527 358 529
rect 361 527 363 529
rect 366 527 368 529
rect 371 527 373 529
rect 376 527 378 529
rect 381 527 383 529
rect 386 527 388 529
rect 391 527 393 529
rect 396 527 398 529
rect 401 527 403 529
rect 406 527 408 529
rect 411 527 413 529
rect 416 527 418 529
rect 421 527 423 529
rect 426 527 428 529
rect 431 527 433 529
rect 436 527 438 529
rect 441 527 443 529
rect 446 527 448 529
rect 451 527 453 529
rect 456 527 458 529
rect 461 527 463 529
rect 466 527 468 529
rect 471 527 473 529
rect 476 527 478 529
rect 481 527 483 529
rect 486 527 488 529
rect 491 527 493 529
rect 496 527 498 529
rect 501 527 503 529
rect 506 527 508 529
rect 511 527 513 529
rect 516 527 518 529
rect 521 527 523 529
rect 526 527 528 529
rect 531 527 533 529
rect 536 527 538 529
rect 541 527 543 529
rect 546 527 548 529
rect 551 527 553 529
rect 556 527 558 529
rect 561 527 563 529
rect 566 527 568 529
rect 571 527 573 529
rect 576 527 578 529
rect 581 527 583 529
rect 586 527 588 529
rect 591 527 593 529
rect 596 527 598 529
rect 601 527 603 529
rect 606 527 608 529
rect 611 527 613 529
rect 616 527 618 529
rect 621 527 623 529
rect 626 527 628 529
rect 631 527 633 529
rect 636 527 638 529
rect 641 527 643 529
rect 646 527 648 529
rect 651 527 653 529
rect 656 527 658 529
rect 661 527 663 529
rect 666 527 668 529
rect 671 527 673 529
rect 676 527 678 529
rect 681 527 683 529
rect 686 527 688 529
rect 691 527 693 529
rect 696 527 698 529
rect 701 527 703 529
rect 706 527 708 529
rect 711 527 713 529
rect 716 527 718 529
rect 721 527 723 529
rect 726 527 728 529
rect 731 527 733 529
rect 736 527 738 529
rect 741 527 743 529
rect 746 527 748 529
rect 751 527 753 529
rect 756 527 758 529
rect 761 527 763 529
rect 766 527 768 529
rect 771 527 773 529
rect 776 527 778 529
rect 781 527 783 529
rect 786 527 788 529
rect 791 527 793 529
rect 796 527 798 529
rect 801 527 803 529
rect 806 527 808 529
rect 811 527 813 529
rect 816 527 818 529
rect 821 527 823 529
rect 826 527 828 529
rect 831 527 833 529
rect 836 527 838 529
rect 841 527 843 529
rect 846 527 848 529
rect 851 527 853 529
rect 856 527 858 529
rect 861 527 863 529
rect 866 527 868 529
rect 871 527 873 529
rect 876 527 878 529
rect 881 527 883 529
rect 886 527 888 529
rect 891 527 893 529
rect 896 527 898 529
rect 901 527 903 529
rect 906 527 908 529
rect 911 527 913 529
rect 916 527 918 529
rect 921 527 923 529
rect 926 527 928 529
rect 931 527 933 529
rect 936 527 938 529
rect 941 527 943 529
rect 946 527 948 529
rect 951 527 953 529
rect 956 527 958 529
rect 961 527 963 529
rect 966 527 968 529
rect 971 527 973 529
rect 976 527 978 529
rect 981 527 983 529
rect 986 527 988 529
rect 991 527 993 529
rect 996 527 998 529
rect 331 522 333 524
rect 336 522 338 524
rect 341 522 343 524
rect 346 522 348 524
rect 351 522 353 524
rect 356 522 358 524
rect 361 522 363 524
rect 366 522 368 524
rect 371 522 373 524
rect 376 522 378 524
rect 381 522 383 524
rect 386 522 388 524
rect 391 522 393 524
rect 396 522 398 524
rect 401 522 403 524
rect 406 522 408 524
rect 411 522 413 524
rect 416 522 418 524
rect 421 522 423 524
rect 426 522 428 524
rect 431 522 433 524
rect 436 522 438 524
rect 441 522 443 524
rect 446 522 448 524
rect 451 522 453 524
rect 456 522 458 524
rect 461 522 463 524
rect 466 522 468 524
rect 471 522 473 524
rect 476 522 478 524
rect 481 522 483 524
rect 486 522 488 524
rect 491 522 493 524
rect 496 522 498 524
rect 501 522 503 524
rect 506 522 508 524
rect 511 522 513 524
rect 516 522 518 524
rect 521 522 523 524
rect 526 522 528 524
rect 531 522 533 524
rect 536 522 538 524
rect 541 522 543 524
rect 546 522 548 524
rect 551 522 553 524
rect 556 522 558 524
rect 561 522 563 524
rect 566 522 568 524
rect 571 522 573 524
rect 576 522 578 524
rect 581 522 583 524
rect 586 522 588 524
rect 591 522 593 524
rect 596 522 598 524
rect 601 522 603 524
rect 606 522 608 524
rect 611 522 613 524
rect 616 522 618 524
rect 621 522 623 524
rect 626 522 628 524
rect 631 522 633 524
rect 636 522 638 524
rect 641 522 643 524
rect 646 522 648 524
rect 651 522 653 524
rect 656 522 658 524
rect 661 522 663 524
rect 666 522 668 524
rect 671 522 673 524
rect 676 522 678 524
rect 681 522 683 524
rect 686 522 688 524
rect 691 522 693 524
rect 696 522 698 524
rect 701 522 703 524
rect 706 522 708 524
rect 711 522 713 524
rect 716 522 718 524
rect 721 522 723 524
rect 726 522 728 524
rect 731 522 733 524
rect 736 522 738 524
rect 741 522 743 524
rect 746 522 748 524
rect 751 522 753 524
rect 756 522 758 524
rect 761 522 763 524
rect 766 522 768 524
rect 771 522 773 524
rect 776 522 778 524
rect 781 522 783 524
rect 786 522 788 524
rect 791 522 793 524
rect 796 522 798 524
rect 801 522 803 524
rect 806 522 808 524
rect 811 522 813 524
rect 816 522 818 524
rect 821 522 823 524
rect 826 522 828 524
rect 831 522 833 524
rect 836 522 838 524
rect 841 522 843 524
rect 846 522 848 524
rect 851 522 853 524
rect 856 522 858 524
rect 861 522 863 524
rect 866 522 868 524
rect 871 522 873 524
rect 876 522 878 524
rect 881 522 883 524
rect 886 522 888 524
rect 891 522 893 524
rect 896 522 898 524
rect 901 522 903 524
rect 906 522 908 524
rect 911 522 913 524
rect 916 522 918 524
rect 921 522 923 524
rect 926 522 928 524
rect 931 522 933 524
rect 936 522 938 524
rect 941 522 943 524
rect 946 522 948 524
rect 951 522 953 524
rect 956 522 958 524
rect 961 522 963 524
rect 966 522 968 524
rect 971 522 973 524
rect 976 522 978 524
rect 981 522 983 524
rect 986 522 988 524
rect 991 522 993 524
rect 996 522 998 524
rect 331 517 333 519
rect 336 517 338 519
rect 341 517 343 519
rect 346 517 348 519
rect 351 517 353 519
rect 356 517 358 519
rect 361 517 363 519
rect 366 517 368 519
rect 371 517 373 519
rect 376 517 378 519
rect 381 517 383 519
rect 386 517 388 519
rect 391 517 393 519
rect 396 517 398 519
rect 401 517 403 519
rect 406 517 408 519
rect 411 517 413 519
rect 416 517 418 519
rect 421 517 423 519
rect 426 517 428 519
rect 431 517 433 519
rect 436 517 438 519
rect 441 517 443 519
rect 446 517 448 519
rect 451 517 453 519
rect 456 517 458 519
rect 461 517 463 519
rect 466 517 468 519
rect 471 517 473 519
rect 476 517 478 519
rect 481 517 483 519
rect 486 517 488 519
rect 491 517 493 519
rect 496 517 498 519
rect 501 517 503 519
rect 506 517 508 519
rect 511 517 513 519
rect 516 517 518 519
rect 521 517 523 519
rect 526 517 528 519
rect 531 517 533 519
rect 536 517 538 519
rect 541 517 543 519
rect 546 517 548 519
rect 551 517 553 519
rect 556 517 558 519
rect 561 517 563 519
rect 566 517 568 519
rect 571 517 573 519
rect 576 517 578 519
rect 581 517 583 519
rect 586 517 588 519
rect 591 517 593 519
rect 596 517 598 519
rect 601 517 603 519
rect 606 517 608 519
rect 611 517 613 519
rect 616 517 618 519
rect 621 517 623 519
rect 626 517 628 519
rect 631 517 633 519
rect 636 517 638 519
rect 641 517 643 519
rect 646 517 648 519
rect 651 517 653 519
rect 656 517 658 519
rect 661 517 663 519
rect 666 517 668 519
rect 671 517 673 519
rect 676 517 678 519
rect 681 517 683 519
rect 686 517 688 519
rect 691 517 693 519
rect 696 517 698 519
rect 701 517 703 519
rect 706 517 708 519
rect 711 517 713 519
rect 716 517 718 519
rect 721 517 723 519
rect 726 517 728 519
rect 731 517 733 519
rect 736 517 738 519
rect 741 517 743 519
rect 746 517 748 519
rect 751 517 753 519
rect 756 517 758 519
rect 761 517 763 519
rect 766 517 768 519
rect 771 517 773 519
rect 776 517 778 519
rect 781 517 783 519
rect 786 517 788 519
rect 791 517 793 519
rect 796 517 798 519
rect 801 517 803 519
rect 806 517 808 519
rect 811 517 813 519
rect 816 517 818 519
rect 821 517 823 519
rect 826 517 828 519
rect 831 517 833 519
rect 836 517 838 519
rect 841 517 843 519
rect 846 517 848 519
rect 851 517 853 519
rect 856 517 858 519
rect 861 517 863 519
rect 866 517 868 519
rect 871 517 873 519
rect 876 517 878 519
rect 881 517 883 519
rect 886 517 888 519
rect 891 517 893 519
rect 896 517 898 519
rect 901 517 903 519
rect 906 517 908 519
rect 911 517 913 519
rect 916 517 918 519
rect 921 517 923 519
rect 926 517 928 519
rect 931 517 933 519
rect 936 517 938 519
rect 941 517 943 519
rect 946 517 948 519
rect 951 517 953 519
rect 956 517 958 519
rect 961 517 963 519
rect 966 517 968 519
rect 971 517 973 519
rect 976 517 978 519
rect 981 517 983 519
rect 986 517 988 519
rect 991 517 993 519
rect 996 517 998 519
rect 331 512 333 514
rect 336 512 338 514
rect 341 512 343 514
rect 346 512 348 514
rect 351 512 353 514
rect 356 512 358 514
rect 361 512 363 514
rect 366 512 368 514
rect 371 512 373 514
rect 376 512 378 514
rect 381 512 383 514
rect 386 512 388 514
rect 391 512 393 514
rect 396 512 398 514
rect 401 512 403 514
rect 406 512 408 514
rect 411 512 413 514
rect 416 512 418 514
rect 421 512 423 514
rect 426 512 428 514
rect 431 512 433 514
rect 436 512 438 514
rect 441 512 443 514
rect 446 512 448 514
rect 451 512 453 514
rect 456 512 458 514
rect 461 512 463 514
rect 466 512 468 514
rect 471 512 473 514
rect 476 512 478 514
rect 481 512 483 514
rect 486 512 488 514
rect 491 512 493 514
rect 496 512 498 514
rect 501 512 503 514
rect 506 512 508 514
rect 511 512 513 514
rect 516 512 518 514
rect 521 512 523 514
rect 526 512 528 514
rect 531 512 533 514
rect 536 512 538 514
rect 541 512 543 514
rect 546 512 548 514
rect 551 512 553 514
rect 556 512 558 514
rect 561 512 563 514
rect 566 512 568 514
rect 571 512 573 514
rect 576 512 578 514
rect 581 512 583 514
rect 586 512 588 514
rect 591 512 593 514
rect 596 512 598 514
rect 601 512 603 514
rect 606 512 608 514
rect 611 512 613 514
rect 616 512 618 514
rect 621 512 623 514
rect 626 512 628 514
rect 631 512 633 514
rect 636 512 638 514
rect 641 512 643 514
rect 646 512 648 514
rect 651 512 653 514
rect 656 512 658 514
rect 661 512 663 514
rect 666 512 668 514
rect 671 512 673 514
rect 676 512 678 514
rect 681 512 683 514
rect 686 512 688 514
rect 691 512 693 514
rect 696 512 698 514
rect 701 512 703 514
rect 706 512 708 514
rect 711 512 713 514
rect 716 512 718 514
rect 721 512 723 514
rect 726 512 728 514
rect 731 512 733 514
rect 736 512 738 514
rect 741 512 743 514
rect 746 512 748 514
rect 751 512 753 514
rect 756 512 758 514
rect 761 512 763 514
rect 766 512 768 514
rect 771 512 773 514
rect 776 512 778 514
rect 781 512 783 514
rect 786 512 788 514
rect 791 512 793 514
rect 796 512 798 514
rect 801 512 803 514
rect 806 512 808 514
rect 811 512 813 514
rect 816 512 818 514
rect 821 512 823 514
rect 826 512 828 514
rect 831 512 833 514
rect 836 512 838 514
rect 841 512 843 514
rect 846 512 848 514
rect 851 512 853 514
rect 856 512 858 514
rect 861 512 863 514
rect 866 512 868 514
rect 871 512 873 514
rect 876 512 878 514
rect 881 512 883 514
rect 886 512 888 514
rect 891 512 893 514
rect 896 512 898 514
rect 901 512 903 514
rect 906 512 908 514
rect 911 512 913 514
rect 916 512 918 514
rect 921 512 923 514
rect 926 512 928 514
rect 931 512 933 514
rect 936 512 938 514
rect 941 512 943 514
rect 946 512 948 514
rect 951 512 953 514
rect 956 512 958 514
rect 961 512 963 514
rect 966 512 968 514
rect 971 512 973 514
rect 976 512 978 514
rect 981 512 983 514
rect 986 512 988 514
rect 991 512 993 514
rect 996 512 998 514
rect 331 507 333 509
rect 336 507 338 509
rect 341 507 343 509
rect 346 507 348 509
rect 351 507 353 509
rect 356 507 358 509
rect 361 507 363 509
rect 366 507 368 509
rect 371 507 373 509
rect 376 507 378 509
rect 381 507 383 509
rect 386 507 388 509
rect 391 507 393 509
rect 396 507 398 509
rect 401 507 403 509
rect 406 507 408 509
rect 411 507 413 509
rect 416 507 418 509
rect 421 507 423 509
rect 426 507 428 509
rect 431 507 433 509
rect 436 507 438 509
rect 441 507 443 509
rect 446 507 448 509
rect 451 507 453 509
rect 456 507 458 509
rect 461 507 463 509
rect 466 507 468 509
rect 471 507 473 509
rect 476 507 478 509
rect 481 507 483 509
rect 486 507 488 509
rect 491 507 493 509
rect 496 507 498 509
rect 501 507 503 509
rect 506 507 508 509
rect 511 507 513 509
rect 516 507 518 509
rect 521 507 523 509
rect 526 507 528 509
rect 531 507 533 509
rect 536 507 538 509
rect 541 507 543 509
rect 546 507 548 509
rect 551 507 553 509
rect 556 507 558 509
rect 561 507 563 509
rect 566 507 568 509
rect 571 507 573 509
rect 576 507 578 509
rect 581 507 583 509
rect 586 507 588 509
rect 591 507 593 509
rect 596 507 598 509
rect 601 507 603 509
rect 606 507 608 509
rect 611 507 613 509
rect 616 507 618 509
rect 621 507 623 509
rect 626 507 628 509
rect 631 507 633 509
rect 636 507 638 509
rect 641 507 643 509
rect 646 507 648 509
rect 651 507 653 509
rect 656 507 658 509
rect 661 507 663 509
rect 666 507 668 509
rect 671 507 673 509
rect 676 507 678 509
rect 681 507 683 509
rect 686 507 688 509
rect 691 507 693 509
rect 696 507 698 509
rect 701 507 703 509
rect 706 507 708 509
rect 711 507 713 509
rect 716 507 718 509
rect 721 507 723 509
rect 726 507 728 509
rect 731 507 733 509
rect 736 507 738 509
rect 741 507 743 509
rect 746 507 748 509
rect 751 507 753 509
rect 756 507 758 509
rect 761 507 763 509
rect 766 507 768 509
rect 771 507 773 509
rect 776 507 778 509
rect 781 507 783 509
rect 786 507 788 509
rect 791 507 793 509
rect 796 507 798 509
rect 801 507 803 509
rect 806 507 808 509
rect 811 507 813 509
rect 816 507 818 509
rect 821 507 823 509
rect 826 507 828 509
rect 831 507 833 509
rect 836 507 838 509
rect 841 507 843 509
rect 846 507 848 509
rect 851 507 853 509
rect 856 507 858 509
rect 861 507 863 509
rect 866 507 868 509
rect 871 507 873 509
rect 876 507 878 509
rect 881 507 883 509
rect 886 507 888 509
rect 891 507 893 509
rect 896 507 898 509
rect 901 507 903 509
rect 906 507 908 509
rect 911 507 913 509
rect 916 507 918 509
rect 921 507 923 509
rect 926 507 928 509
rect 931 507 933 509
rect 936 507 938 509
rect 941 507 943 509
rect 946 507 948 509
rect 951 507 953 509
rect 956 507 958 509
rect 961 507 963 509
rect 966 507 968 509
rect 971 507 973 509
rect 976 507 978 509
rect 981 507 983 509
rect 986 507 988 509
rect 991 507 993 509
rect 996 507 998 509
rect 331 502 333 504
rect 336 502 338 504
rect 341 502 343 504
rect 346 502 348 504
rect 351 502 353 504
rect 356 502 358 504
rect 361 502 363 504
rect 366 502 368 504
rect 371 502 373 504
rect 376 502 378 504
rect 381 502 383 504
rect 386 502 388 504
rect 391 502 393 504
rect 396 502 398 504
rect 401 502 403 504
rect 406 502 408 504
rect 411 502 413 504
rect 416 502 418 504
rect 421 502 423 504
rect 426 502 428 504
rect 431 502 433 504
rect 436 502 438 504
rect 441 502 443 504
rect 446 502 448 504
rect 451 502 453 504
rect 456 502 458 504
rect 461 502 463 504
rect 466 502 468 504
rect 471 502 473 504
rect 476 502 478 504
rect 481 502 483 504
rect 486 502 488 504
rect 491 502 493 504
rect 496 502 498 504
rect 501 502 503 504
rect 506 502 508 504
rect 511 502 513 504
rect 516 502 518 504
rect 521 502 523 504
rect 526 502 528 504
rect 531 502 533 504
rect 536 502 538 504
rect 541 502 543 504
rect 546 502 548 504
rect 551 502 553 504
rect 556 502 558 504
rect 561 502 563 504
rect 566 502 568 504
rect 571 502 573 504
rect 576 502 578 504
rect 581 502 583 504
rect 586 502 588 504
rect 591 502 593 504
rect 596 502 598 504
rect 601 502 603 504
rect 606 502 608 504
rect 611 502 613 504
rect 616 502 618 504
rect 621 502 623 504
rect 626 502 628 504
rect 631 502 633 504
rect 636 502 638 504
rect 641 502 643 504
rect 646 502 648 504
rect 651 502 653 504
rect 656 502 658 504
rect 661 502 663 504
rect 666 502 668 504
rect 671 502 673 504
rect 676 502 678 504
rect 681 502 683 504
rect 686 502 688 504
rect 691 502 693 504
rect 696 502 698 504
rect 701 502 703 504
rect 706 502 708 504
rect 711 502 713 504
rect 716 502 718 504
rect 721 502 723 504
rect 726 502 728 504
rect 731 502 733 504
rect 736 502 738 504
rect 741 502 743 504
rect 746 502 748 504
rect 751 502 753 504
rect 756 502 758 504
rect 761 502 763 504
rect 766 502 768 504
rect 771 502 773 504
rect 776 502 778 504
rect 781 502 783 504
rect 786 502 788 504
rect 791 502 793 504
rect 796 502 798 504
rect 801 502 803 504
rect 806 502 808 504
rect 811 502 813 504
rect 816 502 818 504
rect 821 502 823 504
rect 826 502 828 504
rect 831 502 833 504
rect 836 502 838 504
rect 841 502 843 504
rect 846 502 848 504
rect 851 502 853 504
rect 856 502 858 504
rect 861 502 863 504
rect 866 502 868 504
rect 871 502 873 504
rect 876 502 878 504
rect 881 502 883 504
rect 886 502 888 504
rect 891 502 893 504
rect 896 502 898 504
rect 901 502 903 504
rect 906 502 908 504
rect 911 502 913 504
rect 916 502 918 504
rect 921 502 923 504
rect 926 502 928 504
rect 931 502 933 504
rect 936 502 938 504
rect 941 502 943 504
rect 946 502 948 504
rect 951 502 953 504
rect 956 502 958 504
rect 961 502 963 504
rect 966 502 968 504
rect 971 502 973 504
rect 976 502 978 504
rect 981 502 983 504
rect 986 502 988 504
rect 991 502 993 504
rect 996 502 998 504
rect 331 497 333 499
rect 336 497 338 499
rect 341 497 343 499
rect 346 497 348 499
rect 351 497 353 499
rect 356 497 358 499
rect 361 497 363 499
rect 366 497 368 499
rect 371 497 373 499
rect 376 497 378 499
rect 381 497 383 499
rect 386 497 388 499
rect 391 497 393 499
rect 396 497 398 499
rect 401 497 403 499
rect 406 497 408 499
rect 411 497 413 499
rect 416 497 418 499
rect 421 497 423 499
rect 426 497 428 499
rect 431 497 433 499
rect 436 497 438 499
rect 441 497 443 499
rect 446 497 448 499
rect 451 497 453 499
rect 456 497 458 499
rect 461 497 463 499
rect 466 497 468 499
rect 471 497 473 499
rect 476 497 478 499
rect 481 497 483 499
rect 486 497 488 499
rect 491 497 493 499
rect 496 497 498 499
rect 501 497 503 499
rect 506 497 508 499
rect 511 497 513 499
rect 516 497 518 499
rect 521 497 523 499
rect 526 497 528 499
rect 531 497 533 499
rect 536 497 538 499
rect 541 497 543 499
rect 546 497 548 499
rect 551 497 553 499
rect 556 497 558 499
rect 561 497 563 499
rect 566 497 568 499
rect 571 497 573 499
rect 576 497 578 499
rect 581 497 583 499
rect 586 497 588 499
rect 591 497 593 499
rect 596 497 598 499
rect 601 497 603 499
rect 606 497 608 499
rect 611 497 613 499
rect 616 497 618 499
rect 621 497 623 499
rect 626 497 628 499
rect 631 497 633 499
rect 636 497 638 499
rect 641 497 643 499
rect 646 497 648 499
rect 651 497 653 499
rect 656 497 658 499
rect 661 497 663 499
rect 666 497 668 499
rect 671 497 673 499
rect 676 497 678 499
rect 681 497 683 499
rect 686 497 688 499
rect 691 497 693 499
rect 696 497 698 499
rect 701 497 703 499
rect 706 497 708 499
rect 711 497 713 499
rect 716 497 718 499
rect 721 497 723 499
rect 726 497 728 499
rect 731 497 733 499
rect 736 497 738 499
rect 741 497 743 499
rect 746 497 748 499
rect 751 497 753 499
rect 756 497 758 499
rect 761 497 763 499
rect 766 497 768 499
rect 771 497 773 499
rect 776 497 778 499
rect 781 497 783 499
rect 786 497 788 499
rect 791 497 793 499
rect 796 497 798 499
rect 801 497 803 499
rect 806 497 808 499
rect 811 497 813 499
rect 816 497 818 499
rect 821 497 823 499
rect 826 497 828 499
rect 831 497 833 499
rect 836 497 838 499
rect 841 497 843 499
rect 846 497 848 499
rect 851 497 853 499
rect 856 497 858 499
rect 861 497 863 499
rect 866 497 868 499
rect 871 497 873 499
rect 876 497 878 499
rect 881 497 883 499
rect 886 497 888 499
rect 891 497 893 499
rect 896 497 898 499
rect 901 497 903 499
rect 906 497 908 499
rect 911 497 913 499
rect 916 497 918 499
rect 921 497 923 499
rect 926 497 928 499
rect 931 497 933 499
rect 936 497 938 499
rect 941 497 943 499
rect 946 497 948 499
rect 951 497 953 499
rect 956 497 958 499
rect 961 497 963 499
rect 966 497 968 499
rect 971 497 973 499
rect 976 497 978 499
rect 981 497 983 499
rect 986 497 988 499
rect 991 497 993 499
rect 996 497 998 499
rect 331 492 333 494
rect 336 492 338 494
rect 341 492 343 494
rect 346 492 348 494
rect 351 492 353 494
rect 356 492 358 494
rect 361 492 363 494
rect 366 492 368 494
rect 371 492 373 494
rect 376 492 378 494
rect 381 492 383 494
rect 386 492 388 494
rect 391 492 393 494
rect 396 492 398 494
rect 401 492 403 494
rect 406 492 408 494
rect 411 492 413 494
rect 416 492 418 494
rect 421 492 423 494
rect 426 492 428 494
rect 431 492 433 494
rect 436 492 438 494
rect 441 492 443 494
rect 446 492 448 494
rect 451 492 453 494
rect 456 492 458 494
rect 461 492 463 494
rect 466 492 468 494
rect 471 492 473 494
rect 476 492 478 494
rect 481 492 483 494
rect 486 492 488 494
rect 491 492 493 494
rect 496 492 498 494
rect 501 492 503 494
rect 506 492 508 494
rect 511 492 513 494
rect 516 492 518 494
rect 521 492 523 494
rect 526 492 528 494
rect 531 492 533 494
rect 536 492 538 494
rect 541 492 543 494
rect 546 492 548 494
rect 551 492 553 494
rect 556 492 558 494
rect 561 492 563 494
rect 566 492 568 494
rect 571 492 573 494
rect 576 492 578 494
rect 581 492 583 494
rect 586 492 588 494
rect 591 492 593 494
rect 596 492 598 494
rect 601 492 603 494
rect 606 492 608 494
rect 611 492 613 494
rect 616 492 618 494
rect 621 492 623 494
rect 626 492 628 494
rect 631 492 633 494
rect 636 492 638 494
rect 641 492 643 494
rect 646 492 648 494
rect 651 492 653 494
rect 656 492 658 494
rect 661 492 663 494
rect 666 492 668 494
rect 671 492 673 494
rect 676 492 678 494
rect 681 492 683 494
rect 686 492 688 494
rect 691 492 693 494
rect 696 492 698 494
rect 701 492 703 494
rect 706 492 708 494
rect 711 492 713 494
rect 716 492 718 494
rect 721 492 723 494
rect 726 492 728 494
rect 731 492 733 494
rect 736 492 738 494
rect 741 492 743 494
rect 746 492 748 494
rect 751 492 753 494
rect 756 492 758 494
rect 761 492 763 494
rect 766 492 768 494
rect 771 492 773 494
rect 776 492 778 494
rect 781 492 783 494
rect 786 492 788 494
rect 791 492 793 494
rect 796 492 798 494
rect 801 492 803 494
rect 806 492 808 494
rect 811 492 813 494
rect 816 492 818 494
rect 821 492 823 494
rect 826 492 828 494
rect 831 492 833 494
rect 836 492 838 494
rect 841 492 843 494
rect 846 492 848 494
rect 851 492 853 494
rect 856 492 858 494
rect 861 492 863 494
rect 866 492 868 494
rect 871 492 873 494
rect 876 492 878 494
rect 881 492 883 494
rect 886 492 888 494
rect 891 492 893 494
rect 896 492 898 494
rect 901 492 903 494
rect 906 492 908 494
rect 911 492 913 494
rect 916 492 918 494
rect 921 492 923 494
rect 926 492 928 494
rect 931 492 933 494
rect 936 492 938 494
rect 941 492 943 494
rect 946 492 948 494
rect 951 492 953 494
rect 956 492 958 494
rect 961 492 963 494
rect 966 492 968 494
rect 971 492 973 494
rect 976 492 978 494
rect 981 492 983 494
rect 986 492 988 494
rect 991 492 993 494
rect 996 492 998 494
rect 331 487 333 489
rect 336 487 338 489
rect 341 487 343 489
rect 346 487 348 489
rect 351 487 353 489
rect 356 487 358 489
rect 361 487 363 489
rect 366 487 368 489
rect 371 487 373 489
rect 376 487 378 489
rect 381 487 383 489
rect 386 487 388 489
rect 391 487 393 489
rect 396 487 398 489
rect 401 487 403 489
rect 406 487 408 489
rect 411 487 413 489
rect 416 487 418 489
rect 421 487 423 489
rect 426 487 428 489
rect 431 487 433 489
rect 436 487 438 489
rect 441 487 443 489
rect 446 487 448 489
rect 451 487 453 489
rect 456 487 458 489
rect 461 487 463 489
rect 466 487 468 489
rect 471 487 473 489
rect 476 487 478 489
rect 481 487 483 489
rect 486 487 488 489
rect 491 487 493 489
rect 496 487 498 489
rect 501 487 503 489
rect 506 487 508 489
rect 511 487 513 489
rect 516 487 518 489
rect 521 487 523 489
rect 526 487 528 489
rect 531 487 533 489
rect 536 487 538 489
rect 541 487 543 489
rect 546 487 548 489
rect 551 487 553 489
rect 556 487 558 489
rect 561 487 563 489
rect 566 487 568 489
rect 571 487 573 489
rect 576 487 578 489
rect 581 487 583 489
rect 586 487 588 489
rect 591 487 593 489
rect 596 487 598 489
rect 601 487 603 489
rect 606 487 608 489
rect 611 487 613 489
rect 616 487 618 489
rect 621 487 623 489
rect 626 487 628 489
rect 631 487 633 489
rect 636 487 638 489
rect 641 487 643 489
rect 646 487 648 489
rect 651 487 653 489
rect 656 487 658 489
rect 661 487 663 489
rect 666 487 668 489
rect 671 487 673 489
rect 676 487 678 489
rect 681 487 683 489
rect 686 487 688 489
rect 691 487 693 489
rect 696 487 698 489
rect 701 487 703 489
rect 706 487 708 489
rect 711 487 713 489
rect 716 487 718 489
rect 721 487 723 489
rect 726 487 728 489
rect 731 487 733 489
rect 736 487 738 489
rect 741 487 743 489
rect 746 487 748 489
rect 751 487 753 489
rect 756 487 758 489
rect 761 487 763 489
rect 766 487 768 489
rect 771 487 773 489
rect 776 487 778 489
rect 781 487 783 489
rect 786 487 788 489
rect 791 487 793 489
rect 796 487 798 489
rect 801 487 803 489
rect 806 487 808 489
rect 811 487 813 489
rect 816 487 818 489
rect 821 487 823 489
rect 826 487 828 489
rect 831 487 833 489
rect 836 487 838 489
rect 841 487 843 489
rect 846 487 848 489
rect 851 487 853 489
rect 856 487 858 489
rect 861 487 863 489
rect 866 487 868 489
rect 871 487 873 489
rect 876 487 878 489
rect 881 487 883 489
rect 886 487 888 489
rect 891 487 893 489
rect 896 487 898 489
rect 901 487 903 489
rect 906 487 908 489
rect 911 487 913 489
rect 916 487 918 489
rect 921 487 923 489
rect 926 487 928 489
rect 931 487 933 489
rect 936 487 938 489
rect 941 487 943 489
rect 946 487 948 489
rect 951 487 953 489
rect 956 487 958 489
rect 961 487 963 489
rect 966 487 968 489
rect 971 487 973 489
rect 976 487 978 489
rect 981 487 983 489
rect 986 487 988 489
rect 991 487 993 489
rect 996 487 998 489
rect 331 482 333 484
rect 336 482 338 484
rect 341 482 343 484
rect 346 482 348 484
rect 351 482 353 484
rect 356 482 358 484
rect 361 482 363 484
rect 366 482 368 484
rect 371 482 373 484
rect 376 482 378 484
rect 381 482 383 484
rect 386 482 388 484
rect 391 482 393 484
rect 396 482 398 484
rect 401 482 403 484
rect 406 482 408 484
rect 411 482 413 484
rect 416 482 418 484
rect 421 482 423 484
rect 426 482 428 484
rect 431 482 433 484
rect 436 482 438 484
rect 441 482 443 484
rect 446 482 448 484
rect 451 482 453 484
rect 456 482 458 484
rect 461 482 463 484
rect 466 482 468 484
rect 471 482 473 484
rect 476 482 478 484
rect 481 482 483 484
rect 486 482 488 484
rect 491 482 493 484
rect 496 482 498 484
rect 501 482 503 484
rect 506 482 508 484
rect 511 482 513 484
rect 516 482 518 484
rect 521 482 523 484
rect 526 482 528 484
rect 531 482 533 484
rect 536 482 538 484
rect 541 482 543 484
rect 546 482 548 484
rect 551 482 553 484
rect 556 482 558 484
rect 561 482 563 484
rect 566 482 568 484
rect 571 482 573 484
rect 576 482 578 484
rect 581 482 583 484
rect 586 482 588 484
rect 591 482 593 484
rect 596 482 598 484
rect 601 482 603 484
rect 606 482 608 484
rect 611 482 613 484
rect 616 482 618 484
rect 621 482 623 484
rect 626 482 628 484
rect 631 482 633 484
rect 636 482 638 484
rect 641 482 643 484
rect 646 482 648 484
rect 651 482 653 484
rect 656 482 658 484
rect 661 482 663 484
rect 666 482 668 484
rect 671 482 673 484
rect 676 482 678 484
rect 681 482 683 484
rect 686 482 688 484
rect 691 482 693 484
rect 696 482 698 484
rect 701 482 703 484
rect 706 482 708 484
rect 711 482 713 484
rect 716 482 718 484
rect 721 482 723 484
rect 726 482 728 484
rect 731 482 733 484
rect 736 482 738 484
rect 741 482 743 484
rect 746 482 748 484
rect 751 482 753 484
rect 756 482 758 484
rect 761 482 763 484
rect 766 482 768 484
rect 771 482 773 484
rect 776 482 778 484
rect 781 482 783 484
rect 786 482 788 484
rect 791 482 793 484
rect 796 482 798 484
rect 801 482 803 484
rect 806 482 808 484
rect 811 482 813 484
rect 816 482 818 484
rect 821 482 823 484
rect 826 482 828 484
rect 831 482 833 484
rect 836 482 838 484
rect 841 482 843 484
rect 846 482 848 484
rect 851 482 853 484
rect 856 482 858 484
rect 861 482 863 484
rect 866 482 868 484
rect 871 482 873 484
rect 876 482 878 484
rect 881 482 883 484
rect 886 482 888 484
rect 891 482 893 484
rect 896 482 898 484
rect 901 482 903 484
rect 906 482 908 484
rect 911 482 913 484
rect 916 482 918 484
rect 921 482 923 484
rect 926 482 928 484
rect 931 482 933 484
rect 936 482 938 484
rect 941 482 943 484
rect 946 482 948 484
rect 951 482 953 484
rect 956 482 958 484
rect 961 482 963 484
rect 966 482 968 484
rect 971 482 973 484
rect 976 482 978 484
rect 981 482 983 484
rect 986 482 988 484
rect 991 482 993 484
rect 996 482 998 484
rect 331 477 333 479
rect 336 477 338 479
rect 341 477 343 479
rect 346 477 348 479
rect 351 477 353 479
rect 356 477 358 479
rect 361 477 363 479
rect 366 477 368 479
rect 371 477 373 479
rect 376 477 378 479
rect 381 477 383 479
rect 386 477 388 479
rect 391 477 393 479
rect 396 477 398 479
rect 401 477 403 479
rect 406 477 408 479
rect 411 477 413 479
rect 416 477 418 479
rect 421 477 423 479
rect 426 477 428 479
rect 431 477 433 479
rect 436 477 438 479
rect 441 477 443 479
rect 446 477 448 479
rect 451 477 453 479
rect 456 477 458 479
rect 461 477 463 479
rect 466 477 468 479
rect 471 477 473 479
rect 476 477 478 479
rect 481 477 483 479
rect 486 477 488 479
rect 491 477 493 479
rect 496 477 498 479
rect 501 477 503 479
rect 506 477 508 479
rect 511 477 513 479
rect 516 477 518 479
rect 521 477 523 479
rect 526 477 528 479
rect 531 477 533 479
rect 536 477 538 479
rect 541 477 543 479
rect 546 477 548 479
rect 551 477 553 479
rect 556 477 558 479
rect 561 477 563 479
rect 566 477 568 479
rect 571 477 573 479
rect 576 477 578 479
rect 581 477 583 479
rect 586 477 588 479
rect 591 477 593 479
rect 596 477 598 479
rect 601 477 603 479
rect 606 477 608 479
rect 611 477 613 479
rect 616 477 618 479
rect 621 477 623 479
rect 626 477 628 479
rect 631 477 633 479
rect 636 477 638 479
rect 641 477 643 479
rect 646 477 648 479
rect 651 477 653 479
rect 656 477 658 479
rect 661 477 663 479
rect 666 477 668 479
rect 671 477 673 479
rect 676 477 678 479
rect 681 477 683 479
rect 686 477 688 479
rect 691 477 693 479
rect 696 477 698 479
rect 701 477 703 479
rect 706 477 708 479
rect 711 477 713 479
rect 716 477 718 479
rect 721 477 723 479
rect 726 477 728 479
rect 731 477 733 479
rect 736 477 738 479
rect 741 477 743 479
rect 746 477 748 479
rect 751 477 753 479
rect 756 477 758 479
rect 761 477 763 479
rect 766 477 768 479
rect 771 477 773 479
rect 776 477 778 479
rect 781 477 783 479
rect 786 477 788 479
rect 791 477 793 479
rect 796 477 798 479
rect 801 477 803 479
rect 806 477 808 479
rect 811 477 813 479
rect 816 477 818 479
rect 821 477 823 479
rect 826 477 828 479
rect 831 477 833 479
rect 836 477 838 479
rect 841 477 843 479
rect 846 477 848 479
rect 851 477 853 479
rect 856 477 858 479
rect 861 477 863 479
rect 866 477 868 479
rect 871 477 873 479
rect 876 477 878 479
rect 881 477 883 479
rect 886 477 888 479
rect 891 477 893 479
rect 896 477 898 479
rect 901 477 903 479
rect 906 477 908 479
rect 911 477 913 479
rect 916 477 918 479
rect 921 477 923 479
rect 926 477 928 479
rect 931 477 933 479
rect 936 477 938 479
rect 941 477 943 479
rect 946 477 948 479
rect 951 477 953 479
rect 956 477 958 479
rect 961 477 963 479
rect 966 477 968 479
rect 971 477 973 479
rect 976 477 978 479
rect 981 477 983 479
rect 986 477 988 479
rect 991 477 993 479
rect 996 477 998 479
rect 331 472 333 474
rect 336 472 338 474
rect 341 472 343 474
rect 346 472 348 474
rect 351 472 353 474
rect 356 472 358 474
rect 361 472 363 474
rect 366 472 368 474
rect 371 472 373 474
rect 376 472 378 474
rect 381 472 383 474
rect 386 472 388 474
rect 391 472 393 474
rect 396 472 398 474
rect 401 472 403 474
rect 406 472 408 474
rect 411 472 413 474
rect 416 472 418 474
rect 421 472 423 474
rect 426 472 428 474
rect 431 472 433 474
rect 436 472 438 474
rect 441 472 443 474
rect 446 472 448 474
rect 451 472 453 474
rect 456 472 458 474
rect 461 472 463 474
rect 466 472 468 474
rect 471 472 473 474
rect 476 472 478 474
rect 481 472 483 474
rect 486 472 488 474
rect 491 472 493 474
rect 496 472 498 474
rect 501 472 503 474
rect 506 472 508 474
rect 511 472 513 474
rect 516 472 518 474
rect 521 472 523 474
rect 526 472 528 474
rect 531 472 533 474
rect 536 472 538 474
rect 541 472 543 474
rect 546 472 548 474
rect 551 472 553 474
rect 556 472 558 474
rect 561 472 563 474
rect 566 472 568 474
rect 571 472 573 474
rect 576 472 578 474
rect 581 472 583 474
rect 586 472 588 474
rect 591 472 593 474
rect 596 472 598 474
rect 601 472 603 474
rect 606 472 608 474
rect 611 472 613 474
rect 616 472 618 474
rect 621 472 623 474
rect 626 472 628 474
rect 631 472 633 474
rect 636 472 638 474
rect 641 472 643 474
rect 646 472 648 474
rect 651 472 653 474
rect 656 472 658 474
rect 661 472 663 474
rect 666 472 668 474
rect 671 472 673 474
rect 676 472 678 474
rect 681 472 683 474
rect 686 472 688 474
rect 691 472 693 474
rect 696 472 698 474
rect 701 472 703 474
rect 706 472 708 474
rect 711 472 713 474
rect 716 472 718 474
rect 721 472 723 474
rect 726 472 728 474
rect 731 472 733 474
rect 736 472 738 474
rect 741 472 743 474
rect 746 472 748 474
rect 751 472 753 474
rect 756 472 758 474
rect 761 472 763 474
rect 766 472 768 474
rect 771 472 773 474
rect 776 472 778 474
rect 781 472 783 474
rect 786 472 788 474
rect 791 472 793 474
rect 796 472 798 474
rect 801 472 803 474
rect 806 472 808 474
rect 811 472 813 474
rect 816 472 818 474
rect 821 472 823 474
rect 826 472 828 474
rect 831 472 833 474
rect 836 472 838 474
rect 841 472 843 474
rect 846 472 848 474
rect 851 472 853 474
rect 856 472 858 474
rect 861 472 863 474
rect 866 472 868 474
rect 871 472 873 474
rect 876 472 878 474
rect 881 472 883 474
rect 886 472 888 474
rect 891 472 893 474
rect 896 472 898 474
rect 901 472 903 474
rect 906 472 908 474
rect 911 472 913 474
rect 916 472 918 474
rect 921 472 923 474
rect 926 472 928 474
rect 931 472 933 474
rect 936 472 938 474
rect 941 472 943 474
rect 946 472 948 474
rect 951 472 953 474
rect 956 472 958 474
rect 961 472 963 474
rect 966 472 968 474
rect 971 472 973 474
rect 976 472 978 474
rect 981 472 983 474
rect 986 472 988 474
rect 991 472 993 474
rect 996 472 998 474
rect 331 467 333 469
rect 336 467 338 469
rect 341 467 343 469
rect 346 467 348 469
rect 351 467 353 469
rect 356 467 358 469
rect 361 467 363 469
rect 366 467 368 469
rect 371 467 373 469
rect 376 467 378 469
rect 381 467 383 469
rect 386 467 388 469
rect 391 467 393 469
rect 396 467 398 469
rect 401 467 403 469
rect 406 467 408 469
rect 411 467 413 469
rect 416 467 418 469
rect 421 467 423 469
rect 426 467 428 469
rect 431 467 433 469
rect 436 467 438 469
rect 441 467 443 469
rect 446 467 448 469
rect 451 467 453 469
rect 456 467 458 469
rect 461 467 463 469
rect 466 467 468 469
rect 471 467 473 469
rect 476 467 478 469
rect 481 467 483 469
rect 486 467 488 469
rect 491 467 493 469
rect 496 467 498 469
rect 501 467 503 469
rect 506 467 508 469
rect 511 467 513 469
rect 516 467 518 469
rect 521 467 523 469
rect 526 467 528 469
rect 531 467 533 469
rect 536 467 538 469
rect 541 467 543 469
rect 546 467 548 469
rect 551 467 553 469
rect 556 467 558 469
rect 561 467 563 469
rect 566 467 568 469
rect 571 467 573 469
rect 576 467 578 469
rect 581 467 583 469
rect 586 467 588 469
rect 591 467 593 469
rect 596 467 598 469
rect 601 467 603 469
rect 606 467 608 469
rect 611 467 613 469
rect 616 467 618 469
rect 621 467 623 469
rect 626 467 628 469
rect 631 467 633 469
rect 636 467 638 469
rect 641 467 643 469
rect 646 467 648 469
rect 651 467 653 469
rect 656 467 658 469
rect 661 467 663 469
rect 666 467 668 469
rect 671 467 673 469
rect 676 467 678 469
rect 681 467 683 469
rect 686 467 688 469
rect 691 467 693 469
rect 696 467 698 469
rect 701 467 703 469
rect 706 467 708 469
rect 711 467 713 469
rect 716 467 718 469
rect 721 467 723 469
rect 726 467 728 469
rect 731 467 733 469
rect 736 467 738 469
rect 741 467 743 469
rect 746 467 748 469
rect 751 467 753 469
rect 756 467 758 469
rect 761 467 763 469
rect 766 467 768 469
rect 771 467 773 469
rect 776 467 778 469
rect 781 467 783 469
rect 786 467 788 469
rect 791 467 793 469
rect 796 467 798 469
rect 801 467 803 469
rect 806 467 808 469
rect 811 467 813 469
rect 816 467 818 469
rect 821 467 823 469
rect 826 467 828 469
rect 831 467 833 469
rect 836 467 838 469
rect 841 467 843 469
rect 846 467 848 469
rect 851 467 853 469
rect 856 467 858 469
rect 861 467 863 469
rect 866 467 868 469
rect 871 467 873 469
rect 876 467 878 469
rect 881 467 883 469
rect 886 467 888 469
rect 891 467 893 469
rect 896 467 898 469
rect 901 467 903 469
rect 906 467 908 469
rect 911 467 913 469
rect 916 467 918 469
rect 921 467 923 469
rect 926 467 928 469
rect 931 467 933 469
rect 936 467 938 469
rect 941 467 943 469
rect 946 467 948 469
rect 951 467 953 469
rect 956 467 958 469
rect 961 467 963 469
rect 966 467 968 469
rect 971 467 973 469
rect 976 467 978 469
rect 981 467 983 469
rect 986 467 988 469
rect 991 467 993 469
rect 996 467 998 469
rect 331 462 333 464
rect 336 462 338 464
rect 341 462 343 464
rect 346 462 348 464
rect 351 462 353 464
rect 356 462 358 464
rect 361 462 363 464
rect 366 462 368 464
rect 371 462 373 464
rect 376 462 378 464
rect 381 462 383 464
rect 386 462 388 464
rect 391 462 393 464
rect 396 462 398 464
rect 401 462 403 464
rect 406 462 408 464
rect 411 462 413 464
rect 416 462 418 464
rect 421 462 423 464
rect 426 462 428 464
rect 431 462 433 464
rect 436 462 438 464
rect 441 462 443 464
rect 446 462 448 464
rect 451 462 453 464
rect 456 462 458 464
rect 461 462 463 464
rect 466 462 468 464
rect 471 462 473 464
rect 476 462 478 464
rect 481 462 483 464
rect 486 462 488 464
rect 491 462 493 464
rect 496 462 498 464
rect 501 462 503 464
rect 506 462 508 464
rect 511 462 513 464
rect 516 462 518 464
rect 521 462 523 464
rect 526 462 528 464
rect 531 462 533 464
rect 536 462 538 464
rect 541 462 543 464
rect 546 462 548 464
rect 551 462 553 464
rect 556 462 558 464
rect 561 462 563 464
rect 566 462 568 464
rect 571 462 573 464
rect 576 462 578 464
rect 581 462 583 464
rect 586 462 588 464
rect 591 462 593 464
rect 596 462 598 464
rect 601 462 603 464
rect 606 462 608 464
rect 611 462 613 464
rect 616 462 618 464
rect 621 462 623 464
rect 626 462 628 464
rect 631 462 633 464
rect 636 462 638 464
rect 641 462 643 464
rect 646 462 648 464
rect 651 462 653 464
rect 656 462 658 464
rect 661 462 663 464
rect 666 462 668 464
rect 671 462 673 464
rect 676 462 678 464
rect 681 462 683 464
rect 686 462 688 464
rect 691 462 693 464
rect 696 462 698 464
rect 701 462 703 464
rect 706 462 708 464
rect 711 462 713 464
rect 716 462 718 464
rect 721 462 723 464
rect 726 462 728 464
rect 731 462 733 464
rect 736 462 738 464
rect 741 462 743 464
rect 746 462 748 464
rect 751 462 753 464
rect 756 462 758 464
rect 761 462 763 464
rect 766 462 768 464
rect 771 462 773 464
rect 776 462 778 464
rect 781 462 783 464
rect 786 462 788 464
rect 791 462 793 464
rect 796 462 798 464
rect 801 462 803 464
rect 806 462 808 464
rect 811 462 813 464
rect 816 462 818 464
rect 821 462 823 464
rect 826 462 828 464
rect 831 462 833 464
rect 836 462 838 464
rect 841 462 843 464
rect 846 462 848 464
rect 851 462 853 464
rect 856 462 858 464
rect 861 462 863 464
rect 866 462 868 464
rect 871 462 873 464
rect 876 462 878 464
rect 881 462 883 464
rect 886 462 888 464
rect 891 462 893 464
rect 896 462 898 464
rect 901 462 903 464
rect 906 462 908 464
rect 911 462 913 464
rect 916 462 918 464
rect 921 462 923 464
rect 926 462 928 464
rect 931 462 933 464
rect 936 462 938 464
rect 941 462 943 464
rect 946 462 948 464
rect 951 462 953 464
rect 956 462 958 464
rect 961 462 963 464
rect 966 462 968 464
rect 971 462 973 464
rect 976 462 978 464
rect 981 462 983 464
rect 986 462 988 464
rect 991 462 993 464
rect 996 462 998 464
rect 331 457 333 459
rect 336 457 338 459
rect 341 457 343 459
rect 346 457 348 459
rect 351 457 353 459
rect 356 457 358 459
rect 361 457 363 459
rect 366 457 368 459
rect 371 457 373 459
rect 376 457 378 459
rect 381 457 383 459
rect 386 457 388 459
rect 391 457 393 459
rect 396 457 398 459
rect 401 457 403 459
rect 406 457 408 459
rect 411 457 413 459
rect 416 457 418 459
rect 421 457 423 459
rect 426 457 428 459
rect 431 457 433 459
rect 436 457 438 459
rect 441 457 443 459
rect 446 457 448 459
rect 451 457 453 459
rect 456 457 458 459
rect 461 457 463 459
rect 466 457 468 459
rect 471 457 473 459
rect 476 457 478 459
rect 481 457 483 459
rect 486 457 488 459
rect 491 457 493 459
rect 496 457 498 459
rect 501 457 503 459
rect 506 457 508 459
rect 511 457 513 459
rect 516 457 518 459
rect 521 457 523 459
rect 526 457 528 459
rect 531 457 533 459
rect 536 457 538 459
rect 541 457 543 459
rect 546 457 548 459
rect 551 457 553 459
rect 556 457 558 459
rect 561 457 563 459
rect 566 457 568 459
rect 571 457 573 459
rect 576 457 578 459
rect 581 457 583 459
rect 586 457 588 459
rect 591 457 593 459
rect 596 457 598 459
rect 601 457 603 459
rect 606 457 608 459
rect 611 457 613 459
rect 616 457 618 459
rect 621 457 623 459
rect 626 457 628 459
rect 631 457 633 459
rect 636 457 638 459
rect 641 457 643 459
rect 646 457 648 459
rect 651 457 653 459
rect 656 457 658 459
rect 661 457 663 459
rect 666 457 668 459
rect 671 457 673 459
rect 676 457 678 459
rect 681 457 683 459
rect 686 457 688 459
rect 691 457 693 459
rect 696 457 698 459
rect 701 457 703 459
rect 706 457 708 459
rect 711 457 713 459
rect 716 457 718 459
rect 721 457 723 459
rect 726 457 728 459
rect 731 457 733 459
rect 736 457 738 459
rect 741 457 743 459
rect 746 457 748 459
rect 751 457 753 459
rect 756 457 758 459
rect 761 457 763 459
rect 766 457 768 459
rect 771 457 773 459
rect 776 457 778 459
rect 781 457 783 459
rect 786 457 788 459
rect 791 457 793 459
rect 796 457 798 459
rect 801 457 803 459
rect 806 457 808 459
rect 811 457 813 459
rect 816 457 818 459
rect 821 457 823 459
rect 826 457 828 459
rect 831 457 833 459
rect 836 457 838 459
rect 841 457 843 459
rect 846 457 848 459
rect 851 457 853 459
rect 856 457 858 459
rect 861 457 863 459
rect 866 457 868 459
rect 871 457 873 459
rect 876 457 878 459
rect 881 457 883 459
rect 886 457 888 459
rect 891 457 893 459
rect 896 457 898 459
rect 901 457 903 459
rect 906 457 908 459
rect 911 457 913 459
rect 916 457 918 459
rect 921 457 923 459
rect 926 457 928 459
rect 931 457 933 459
rect 936 457 938 459
rect 941 457 943 459
rect 946 457 948 459
rect 951 457 953 459
rect 956 457 958 459
rect 961 457 963 459
rect 966 457 968 459
rect 971 457 973 459
rect 976 457 978 459
rect 981 457 983 459
rect 986 457 988 459
rect 991 457 993 459
rect 996 457 998 459
rect 331 452 333 454
rect 336 452 338 454
rect 341 452 343 454
rect 346 452 348 454
rect 351 452 353 454
rect 356 452 358 454
rect 361 452 363 454
rect 366 452 368 454
rect 371 452 373 454
rect 376 452 378 454
rect 381 452 383 454
rect 386 452 388 454
rect 391 452 393 454
rect 396 452 398 454
rect 401 452 403 454
rect 406 452 408 454
rect 411 452 413 454
rect 416 452 418 454
rect 421 452 423 454
rect 426 452 428 454
rect 431 452 433 454
rect 436 452 438 454
rect 441 452 443 454
rect 446 452 448 454
rect 451 452 453 454
rect 456 452 458 454
rect 461 452 463 454
rect 466 452 468 454
rect 471 452 473 454
rect 476 452 478 454
rect 481 452 483 454
rect 486 452 488 454
rect 491 452 493 454
rect 496 452 498 454
rect 501 452 503 454
rect 506 452 508 454
rect 511 452 513 454
rect 516 452 518 454
rect 521 452 523 454
rect 526 452 528 454
rect 531 452 533 454
rect 536 452 538 454
rect 541 452 543 454
rect 546 452 548 454
rect 551 452 553 454
rect 556 452 558 454
rect 561 452 563 454
rect 566 452 568 454
rect 571 452 573 454
rect 576 452 578 454
rect 581 452 583 454
rect 586 452 588 454
rect 591 452 593 454
rect 596 452 598 454
rect 601 452 603 454
rect 606 452 608 454
rect 611 452 613 454
rect 616 452 618 454
rect 621 452 623 454
rect 626 452 628 454
rect 631 452 633 454
rect 636 452 638 454
rect 641 452 643 454
rect 646 452 648 454
rect 651 452 653 454
rect 656 452 658 454
rect 661 452 663 454
rect 666 452 668 454
rect 671 452 673 454
rect 676 452 678 454
rect 681 452 683 454
rect 686 452 688 454
rect 691 452 693 454
rect 696 452 698 454
rect 701 452 703 454
rect 706 452 708 454
rect 711 452 713 454
rect 716 452 718 454
rect 721 452 723 454
rect 726 452 728 454
rect 731 452 733 454
rect 736 452 738 454
rect 741 452 743 454
rect 746 452 748 454
rect 751 452 753 454
rect 756 452 758 454
rect 761 452 763 454
rect 766 452 768 454
rect 771 452 773 454
rect 776 452 778 454
rect 781 452 783 454
rect 786 452 788 454
rect 791 452 793 454
rect 796 452 798 454
rect 801 452 803 454
rect 806 452 808 454
rect 811 452 813 454
rect 816 452 818 454
rect 821 452 823 454
rect 826 452 828 454
rect 831 452 833 454
rect 836 452 838 454
rect 841 452 843 454
rect 846 452 848 454
rect 851 452 853 454
rect 856 452 858 454
rect 861 452 863 454
rect 866 452 868 454
rect 871 452 873 454
rect 876 452 878 454
rect 881 452 883 454
rect 886 452 888 454
rect 891 452 893 454
rect 896 452 898 454
rect 901 452 903 454
rect 906 452 908 454
rect 911 452 913 454
rect 916 452 918 454
rect 921 452 923 454
rect 926 452 928 454
rect 931 452 933 454
rect 936 452 938 454
rect 941 452 943 454
rect 946 452 948 454
rect 951 452 953 454
rect 956 452 958 454
rect 961 452 963 454
rect 966 452 968 454
rect 971 452 973 454
rect 976 452 978 454
rect 981 452 983 454
rect 986 452 988 454
rect 991 452 993 454
rect 996 452 998 454
rect 331 447 333 449
rect 336 447 338 449
rect 341 447 343 449
rect 346 447 348 449
rect 351 447 353 449
rect 356 447 358 449
rect 361 447 363 449
rect 366 447 368 449
rect 371 447 373 449
rect 376 447 378 449
rect 381 447 383 449
rect 386 447 388 449
rect 391 447 393 449
rect 396 447 398 449
rect 401 447 403 449
rect 406 447 408 449
rect 411 447 413 449
rect 416 447 418 449
rect 421 447 423 449
rect 426 447 428 449
rect 431 447 433 449
rect 436 447 438 449
rect 441 447 443 449
rect 446 447 448 449
rect 451 447 453 449
rect 456 447 458 449
rect 461 447 463 449
rect 466 447 468 449
rect 471 447 473 449
rect 476 447 478 449
rect 481 447 483 449
rect 486 447 488 449
rect 491 447 493 449
rect 496 447 498 449
rect 501 447 503 449
rect 506 447 508 449
rect 511 447 513 449
rect 516 447 518 449
rect 521 447 523 449
rect 526 447 528 449
rect 531 447 533 449
rect 536 447 538 449
rect 541 447 543 449
rect 546 447 548 449
rect 551 447 553 449
rect 556 447 558 449
rect 561 447 563 449
rect 566 447 568 449
rect 571 447 573 449
rect 576 447 578 449
rect 581 447 583 449
rect 586 447 588 449
rect 591 447 593 449
rect 596 447 598 449
rect 601 447 603 449
rect 606 447 608 449
rect 611 447 613 449
rect 616 447 618 449
rect 621 447 623 449
rect 626 447 628 449
rect 631 447 633 449
rect 636 447 638 449
rect 641 447 643 449
rect 646 447 648 449
rect 651 447 653 449
rect 656 447 658 449
rect 661 447 663 449
rect 666 447 668 449
rect 671 447 673 449
rect 676 447 678 449
rect 681 447 683 449
rect 686 447 688 449
rect 691 447 693 449
rect 696 447 698 449
rect 701 447 703 449
rect 706 447 708 449
rect 711 447 713 449
rect 716 447 718 449
rect 721 447 723 449
rect 726 447 728 449
rect 731 447 733 449
rect 736 447 738 449
rect 741 447 743 449
rect 746 447 748 449
rect 751 447 753 449
rect 756 447 758 449
rect 761 447 763 449
rect 766 447 768 449
rect 771 447 773 449
rect 776 447 778 449
rect 781 447 783 449
rect 786 447 788 449
rect 791 447 793 449
rect 796 447 798 449
rect 801 447 803 449
rect 806 447 808 449
rect 811 447 813 449
rect 816 447 818 449
rect 821 447 823 449
rect 826 447 828 449
rect 831 447 833 449
rect 836 447 838 449
rect 841 447 843 449
rect 846 447 848 449
rect 851 447 853 449
rect 856 447 858 449
rect 861 447 863 449
rect 866 447 868 449
rect 871 447 873 449
rect 876 447 878 449
rect 881 447 883 449
rect 886 447 888 449
rect 891 447 893 449
rect 896 447 898 449
rect 901 447 903 449
rect 906 447 908 449
rect 911 447 913 449
rect 916 447 918 449
rect 921 447 923 449
rect 926 447 928 449
rect 931 447 933 449
rect 936 447 938 449
rect 941 447 943 449
rect 946 447 948 449
rect 951 447 953 449
rect 956 447 958 449
rect 961 447 963 449
rect 966 447 968 449
rect 971 447 973 449
rect 976 447 978 449
rect 981 447 983 449
rect 986 447 988 449
rect 991 447 993 449
rect 996 447 998 449
rect 331 442 333 444
rect 336 442 338 444
rect 341 442 343 444
rect 346 442 348 444
rect 351 442 353 444
rect 356 442 358 444
rect 361 442 363 444
rect 366 442 368 444
rect 371 442 373 444
rect 376 442 378 444
rect 381 442 383 444
rect 386 442 388 444
rect 391 442 393 444
rect 396 442 398 444
rect 401 442 403 444
rect 406 442 408 444
rect 411 442 413 444
rect 416 442 418 444
rect 421 442 423 444
rect 426 442 428 444
rect 431 442 433 444
rect 436 442 438 444
rect 441 442 443 444
rect 446 442 448 444
rect 451 442 453 444
rect 456 442 458 444
rect 461 442 463 444
rect 466 442 468 444
rect 471 442 473 444
rect 476 442 478 444
rect 481 442 483 444
rect 486 442 488 444
rect 491 442 493 444
rect 496 442 498 444
rect 501 442 503 444
rect 506 442 508 444
rect 511 442 513 444
rect 516 442 518 444
rect 521 442 523 444
rect 526 442 528 444
rect 531 442 533 444
rect 536 442 538 444
rect 541 442 543 444
rect 546 442 548 444
rect 551 442 553 444
rect 556 442 558 444
rect 561 442 563 444
rect 566 442 568 444
rect 571 442 573 444
rect 576 442 578 444
rect 581 442 583 444
rect 586 442 588 444
rect 591 442 593 444
rect 596 442 598 444
rect 601 442 603 444
rect 606 442 608 444
rect 611 442 613 444
rect 616 442 618 444
rect 621 442 623 444
rect 626 442 628 444
rect 631 442 633 444
rect 636 442 638 444
rect 641 442 643 444
rect 646 442 648 444
rect 651 442 653 444
rect 656 442 658 444
rect 661 442 663 444
rect 666 442 668 444
rect 671 442 673 444
rect 676 442 678 444
rect 681 442 683 444
rect 686 442 688 444
rect 691 442 693 444
rect 696 442 698 444
rect 701 442 703 444
rect 706 442 708 444
rect 711 442 713 444
rect 716 442 718 444
rect 721 442 723 444
rect 726 442 728 444
rect 731 442 733 444
rect 736 442 738 444
rect 741 442 743 444
rect 746 442 748 444
rect 751 442 753 444
rect 756 442 758 444
rect 761 442 763 444
rect 766 442 768 444
rect 771 442 773 444
rect 776 442 778 444
rect 781 442 783 444
rect 786 442 788 444
rect 791 442 793 444
rect 796 442 798 444
rect 801 442 803 444
rect 806 442 808 444
rect 811 442 813 444
rect 816 442 818 444
rect 821 442 823 444
rect 826 442 828 444
rect 831 442 833 444
rect 836 442 838 444
rect 841 442 843 444
rect 846 442 848 444
rect 851 442 853 444
rect 856 442 858 444
rect 861 442 863 444
rect 866 442 868 444
rect 871 442 873 444
rect 876 442 878 444
rect 881 442 883 444
rect 886 442 888 444
rect 891 442 893 444
rect 896 442 898 444
rect 901 442 903 444
rect 906 442 908 444
rect 911 442 913 444
rect 916 442 918 444
rect 921 442 923 444
rect 926 442 928 444
rect 931 442 933 444
rect 936 442 938 444
rect 941 442 943 444
rect 946 442 948 444
rect 951 442 953 444
rect 956 442 958 444
rect 961 442 963 444
rect 966 442 968 444
rect 971 442 973 444
rect 976 442 978 444
rect 981 442 983 444
rect 986 442 988 444
rect 991 442 993 444
rect 996 442 998 444
rect 331 421 333 423
rect 336 421 338 423
rect 341 421 343 423
rect 346 421 348 423
rect 351 421 353 423
rect 356 421 358 423
rect 361 421 363 423
rect 366 421 368 423
rect 371 421 373 423
rect 376 421 378 423
rect 381 421 383 423
rect 386 421 388 423
rect 391 421 393 423
rect 396 421 398 423
rect 401 421 403 423
rect 406 421 408 423
rect 411 421 413 423
rect 416 421 418 423
rect 421 421 423 423
rect 426 421 428 423
rect 431 421 433 423
rect 436 421 438 423
rect 441 421 443 423
rect 446 421 448 423
rect 451 421 453 423
rect 456 421 458 423
rect 461 421 463 423
rect 466 421 468 423
rect 471 421 473 423
rect 476 421 478 423
rect 481 421 483 423
rect 486 421 488 423
rect 491 421 493 423
rect 496 421 498 423
rect 501 421 503 423
rect 506 421 508 423
rect 511 421 513 423
rect 516 421 518 423
rect 521 421 523 423
rect 526 421 528 423
rect 531 421 533 423
rect 536 421 538 423
rect 541 421 543 423
rect 546 421 548 423
rect 551 421 553 423
rect 556 421 558 423
rect 331 416 333 418
rect 336 416 338 418
rect 341 416 343 418
rect 346 416 348 418
rect 351 416 353 418
rect 356 416 358 418
rect 361 416 363 418
rect 366 416 368 418
rect 371 416 373 418
rect 376 416 378 418
rect 381 416 383 418
rect 386 416 388 418
rect 391 416 393 418
rect 396 416 398 418
rect 401 416 403 418
rect 406 416 408 418
rect 411 416 413 418
rect 416 416 418 418
rect 421 416 423 418
rect 426 416 428 418
rect 431 416 433 418
rect 436 416 438 418
rect 441 416 443 418
rect 446 416 448 418
rect 451 416 453 418
rect 456 416 458 418
rect 461 416 463 418
rect 466 416 468 418
rect 471 416 473 418
rect 476 416 478 418
rect 481 416 483 418
rect 486 416 488 418
rect 491 416 493 418
rect 496 416 498 418
rect 501 416 503 418
rect 506 416 508 418
rect 511 416 513 418
rect 516 416 518 418
rect 521 416 523 418
rect 526 416 528 418
rect 531 416 533 418
rect 536 416 538 418
rect 541 416 543 418
rect 546 416 548 418
rect 551 416 553 418
rect 556 416 558 418
rect 331 411 333 413
rect 336 411 338 413
rect 341 411 343 413
rect 346 411 348 413
rect 351 411 353 413
rect 356 411 358 413
rect 361 411 363 413
rect 366 411 368 413
rect 371 411 373 413
rect 376 411 378 413
rect 381 411 383 413
rect 386 411 388 413
rect 391 411 393 413
rect 396 411 398 413
rect 401 411 403 413
rect 406 411 408 413
rect 411 411 413 413
rect 416 411 418 413
rect 421 411 423 413
rect 426 411 428 413
rect 431 411 433 413
rect 436 411 438 413
rect 441 411 443 413
rect 446 411 448 413
rect 451 411 453 413
rect 456 411 458 413
rect 461 411 463 413
rect 466 411 468 413
rect 471 411 473 413
rect 476 411 478 413
rect 481 411 483 413
rect 486 411 488 413
rect 491 411 493 413
rect 496 411 498 413
rect 501 411 503 413
rect 506 411 508 413
rect 511 411 513 413
rect 516 411 518 413
rect 521 411 523 413
rect 526 411 528 413
rect 531 411 533 413
rect 536 411 538 413
rect 541 411 543 413
rect 546 411 548 413
rect 551 411 553 413
rect 556 411 558 413
rect 331 406 333 408
rect 336 406 338 408
rect 341 406 343 408
rect 346 406 348 408
rect 351 406 353 408
rect 356 406 358 408
rect 361 406 363 408
rect 366 406 368 408
rect 371 406 373 408
rect 376 406 378 408
rect 381 406 383 408
rect 386 406 388 408
rect 391 406 393 408
rect 396 406 398 408
rect 401 406 403 408
rect 406 406 408 408
rect 411 406 413 408
rect 416 406 418 408
rect 421 406 423 408
rect 426 406 428 408
rect 431 406 433 408
rect 436 406 438 408
rect 441 406 443 408
rect 446 406 448 408
rect 451 406 453 408
rect 456 406 458 408
rect 461 406 463 408
rect 466 406 468 408
rect 471 406 473 408
rect 476 406 478 408
rect 481 406 483 408
rect 486 406 488 408
rect 491 406 493 408
rect 496 406 498 408
rect 501 406 503 408
rect 506 406 508 408
rect 511 406 513 408
rect 516 406 518 408
rect 521 406 523 408
rect 526 406 528 408
rect 531 406 533 408
rect 536 406 538 408
rect 541 406 543 408
rect 546 406 548 408
rect 551 406 553 408
rect 556 406 558 408
rect 331 401 333 403
rect 336 401 338 403
rect 341 401 343 403
rect 346 401 348 403
rect 351 401 353 403
rect 356 401 358 403
rect 361 401 363 403
rect 366 401 368 403
rect 371 401 373 403
rect 376 401 378 403
rect 381 401 383 403
rect 386 401 388 403
rect 391 401 393 403
rect 396 401 398 403
rect 401 401 403 403
rect 406 401 408 403
rect 411 401 413 403
rect 416 401 418 403
rect 421 401 423 403
rect 426 401 428 403
rect 431 401 433 403
rect 436 401 438 403
rect 441 401 443 403
rect 446 401 448 403
rect 451 401 453 403
rect 456 401 458 403
rect 461 401 463 403
rect 466 401 468 403
rect 471 401 473 403
rect 476 401 478 403
rect 481 401 483 403
rect 486 401 488 403
rect 491 401 493 403
rect 496 401 498 403
rect 501 401 503 403
rect 506 401 508 403
rect 511 401 513 403
rect 516 401 518 403
rect 521 401 523 403
rect 526 401 528 403
rect 531 401 533 403
rect 536 401 538 403
rect 541 401 543 403
rect 546 401 548 403
rect 551 401 553 403
rect 556 401 558 403
rect 331 396 333 398
rect 336 396 338 398
rect 341 396 343 398
rect 346 396 348 398
rect 351 396 353 398
rect 356 396 358 398
rect 361 396 363 398
rect 366 396 368 398
rect 371 396 373 398
rect 376 396 378 398
rect 381 396 383 398
rect 386 396 388 398
rect 391 396 393 398
rect 396 396 398 398
rect 401 396 403 398
rect 406 396 408 398
rect 411 396 413 398
rect 416 396 418 398
rect 421 396 423 398
rect 426 396 428 398
rect 431 396 433 398
rect 436 396 438 398
rect 441 396 443 398
rect 446 396 448 398
rect 451 396 453 398
rect 456 396 458 398
rect 461 396 463 398
rect 466 396 468 398
rect 471 396 473 398
rect 476 396 478 398
rect 481 396 483 398
rect 486 396 488 398
rect 491 396 493 398
rect 496 396 498 398
rect 501 396 503 398
rect 506 396 508 398
rect 511 396 513 398
rect 516 396 518 398
rect 521 396 523 398
rect 526 396 528 398
rect 531 396 533 398
rect 536 396 538 398
rect 541 396 543 398
rect 546 396 548 398
rect 551 396 553 398
rect 556 396 558 398
rect 331 391 333 393
rect 336 391 338 393
rect 341 391 343 393
rect 346 391 348 393
rect 351 391 353 393
rect 356 391 358 393
rect 361 391 363 393
rect 366 391 368 393
rect 371 391 373 393
rect 376 391 378 393
rect 381 391 383 393
rect 386 391 388 393
rect 391 391 393 393
rect 396 391 398 393
rect 401 391 403 393
rect 406 391 408 393
rect 411 391 413 393
rect 416 391 418 393
rect 421 391 423 393
rect 426 391 428 393
rect 431 391 433 393
rect 436 391 438 393
rect 441 391 443 393
rect 446 391 448 393
rect 451 391 453 393
rect 456 391 458 393
rect 461 391 463 393
rect 466 391 468 393
rect 471 391 473 393
rect 476 391 478 393
rect 481 391 483 393
rect 486 391 488 393
rect 491 391 493 393
rect 496 391 498 393
rect 501 391 503 393
rect 506 391 508 393
rect 511 391 513 393
rect 516 391 518 393
rect 521 391 523 393
rect 526 391 528 393
rect 531 391 533 393
rect 536 391 538 393
rect 541 391 543 393
rect 546 391 548 393
rect 551 391 553 393
rect 556 391 558 393
rect 331 386 333 388
rect 336 386 338 388
rect 341 386 343 388
rect 346 386 348 388
rect 351 386 353 388
rect 356 386 358 388
rect 361 386 363 388
rect 366 386 368 388
rect 371 386 373 388
rect 376 386 378 388
rect 381 386 383 388
rect 386 386 388 388
rect 391 386 393 388
rect 396 386 398 388
rect 401 386 403 388
rect 406 386 408 388
rect 411 386 413 388
rect 416 386 418 388
rect 421 386 423 388
rect 426 386 428 388
rect 431 386 433 388
rect 436 386 438 388
rect 441 386 443 388
rect 446 386 448 388
rect 451 386 453 388
rect 456 386 458 388
rect 461 386 463 388
rect 466 386 468 388
rect 471 386 473 388
rect 476 386 478 388
rect 481 386 483 388
rect 486 386 488 388
rect 491 386 493 388
rect 496 386 498 388
rect 501 386 503 388
rect 506 386 508 388
rect 511 386 513 388
rect 516 386 518 388
rect 521 386 523 388
rect 526 386 528 388
rect 531 386 533 388
rect 536 386 538 388
rect 541 386 543 388
rect 546 386 548 388
rect 551 386 553 388
rect 556 386 558 388
rect 331 381 333 383
rect 336 381 338 383
rect 341 381 343 383
rect 346 381 348 383
rect 351 381 353 383
rect 356 381 358 383
rect 361 381 363 383
rect 366 381 368 383
rect 371 381 373 383
rect 376 381 378 383
rect 381 381 383 383
rect 386 381 388 383
rect 391 381 393 383
rect 396 381 398 383
rect 401 381 403 383
rect 406 381 408 383
rect 411 381 413 383
rect 416 381 418 383
rect 421 381 423 383
rect 426 381 428 383
rect 431 381 433 383
rect 436 381 438 383
rect 441 381 443 383
rect 446 381 448 383
rect 451 381 453 383
rect 456 381 458 383
rect 461 381 463 383
rect 466 381 468 383
rect 471 381 473 383
rect 476 381 478 383
rect 481 381 483 383
rect 486 381 488 383
rect 491 381 493 383
rect 496 381 498 383
rect 501 381 503 383
rect 506 381 508 383
rect 511 381 513 383
rect 516 381 518 383
rect 521 381 523 383
rect 526 381 528 383
rect 531 381 533 383
rect 536 381 538 383
rect 541 381 543 383
rect 546 381 548 383
rect 551 381 553 383
rect 556 381 558 383
rect 331 376 333 378
rect 336 376 338 378
rect 341 376 343 378
rect 346 376 348 378
rect 351 376 353 378
rect 356 376 358 378
rect 361 376 363 378
rect 366 376 368 378
rect 371 376 373 378
rect 376 376 378 378
rect 381 376 383 378
rect 386 376 388 378
rect 391 376 393 378
rect 396 376 398 378
rect 401 376 403 378
rect 406 376 408 378
rect 411 376 413 378
rect 416 376 418 378
rect 421 376 423 378
rect 426 376 428 378
rect 431 376 433 378
rect 436 376 438 378
rect 441 376 443 378
rect 446 376 448 378
rect 451 376 453 378
rect 456 376 458 378
rect 461 376 463 378
rect 466 376 468 378
rect 471 376 473 378
rect 476 376 478 378
rect 481 376 483 378
rect 486 376 488 378
rect 491 376 493 378
rect 496 376 498 378
rect 501 376 503 378
rect 506 376 508 378
rect 511 376 513 378
rect 516 376 518 378
rect 521 376 523 378
rect 526 376 528 378
rect 531 376 533 378
rect 536 376 538 378
rect 541 376 543 378
rect 546 376 548 378
rect 551 376 553 378
rect 556 376 558 378
rect 331 371 333 373
rect 336 371 338 373
rect 341 371 343 373
rect 346 371 348 373
rect 351 371 353 373
rect 356 371 358 373
rect 361 371 363 373
rect 366 371 368 373
rect 371 371 373 373
rect 376 371 378 373
rect 381 371 383 373
rect 386 371 388 373
rect 391 371 393 373
rect 396 371 398 373
rect 401 371 403 373
rect 406 371 408 373
rect 411 371 413 373
rect 416 371 418 373
rect 421 371 423 373
rect 426 371 428 373
rect 431 371 433 373
rect 436 371 438 373
rect 441 371 443 373
rect 446 371 448 373
rect 451 371 453 373
rect 456 371 458 373
rect 461 371 463 373
rect 466 371 468 373
rect 471 371 473 373
rect 476 371 478 373
rect 481 371 483 373
rect 486 371 488 373
rect 491 371 493 373
rect 496 371 498 373
rect 501 371 503 373
rect 506 371 508 373
rect 511 371 513 373
rect 516 371 518 373
rect 521 371 523 373
rect 526 371 528 373
rect 531 371 533 373
rect 536 371 538 373
rect 541 371 543 373
rect 546 371 548 373
rect 551 371 553 373
rect 556 371 558 373
rect 331 366 333 368
rect 336 366 338 368
rect 341 366 343 368
rect 346 366 348 368
rect 351 366 353 368
rect 356 366 358 368
rect 361 366 363 368
rect 366 366 368 368
rect 371 366 373 368
rect 376 366 378 368
rect 381 366 383 368
rect 386 366 388 368
rect 391 366 393 368
rect 396 366 398 368
rect 401 366 403 368
rect 406 366 408 368
rect 411 366 413 368
rect 416 366 418 368
rect 421 366 423 368
rect 426 366 428 368
rect 431 366 433 368
rect 436 366 438 368
rect 441 366 443 368
rect 446 366 448 368
rect 451 366 453 368
rect 456 366 458 368
rect 461 366 463 368
rect 466 366 468 368
rect 471 366 473 368
rect 476 366 478 368
rect 481 366 483 368
rect 486 366 488 368
rect 491 366 493 368
rect 496 366 498 368
rect 501 366 503 368
rect 506 366 508 368
rect 511 366 513 368
rect 516 366 518 368
rect 521 366 523 368
rect 526 366 528 368
rect 531 366 533 368
rect 536 366 538 368
rect 541 366 543 368
rect 546 366 548 368
rect 551 366 553 368
rect 556 366 558 368
rect 331 361 333 363
rect 336 361 338 363
rect 341 361 343 363
rect 346 361 348 363
rect 351 361 353 363
rect 356 361 358 363
rect 361 361 363 363
rect 366 361 368 363
rect 371 361 373 363
rect 376 361 378 363
rect 381 361 383 363
rect 386 361 388 363
rect 391 361 393 363
rect 396 361 398 363
rect 401 361 403 363
rect 406 361 408 363
rect 411 361 413 363
rect 416 361 418 363
rect 421 361 423 363
rect 426 361 428 363
rect 431 361 433 363
rect 436 361 438 363
rect 441 361 443 363
rect 446 361 448 363
rect 451 361 453 363
rect 456 361 458 363
rect 461 361 463 363
rect 466 361 468 363
rect 471 361 473 363
rect 476 361 478 363
rect 481 361 483 363
rect 486 361 488 363
rect 491 361 493 363
rect 496 361 498 363
rect 501 361 503 363
rect 506 361 508 363
rect 511 361 513 363
rect 516 361 518 363
rect 521 361 523 363
rect 526 361 528 363
rect 531 361 533 363
rect 536 361 538 363
rect 541 361 543 363
rect 546 361 548 363
rect 551 361 553 363
rect 556 361 558 363
rect 331 356 333 358
rect 336 356 338 358
rect 341 356 343 358
rect 346 356 348 358
rect 351 356 353 358
rect 356 356 358 358
rect 361 356 363 358
rect 366 356 368 358
rect 371 356 373 358
rect 376 356 378 358
rect 381 356 383 358
rect 386 356 388 358
rect 391 356 393 358
rect 396 356 398 358
rect 401 356 403 358
rect 406 356 408 358
rect 411 356 413 358
rect 416 356 418 358
rect 421 356 423 358
rect 426 356 428 358
rect 431 356 433 358
rect 436 356 438 358
rect 441 356 443 358
rect 446 356 448 358
rect 451 356 453 358
rect 456 356 458 358
rect 461 356 463 358
rect 466 356 468 358
rect 471 356 473 358
rect 476 356 478 358
rect 481 356 483 358
rect 486 356 488 358
rect 491 356 493 358
rect 496 356 498 358
rect 501 356 503 358
rect 506 356 508 358
rect 511 356 513 358
rect 516 356 518 358
rect 521 356 523 358
rect 526 356 528 358
rect 531 356 533 358
rect 536 356 538 358
rect 541 356 543 358
rect 546 356 548 358
rect 551 356 553 358
rect 556 356 558 358
rect 331 351 333 353
rect 336 351 338 353
rect 341 351 343 353
rect 346 351 348 353
rect 351 351 353 353
rect 356 351 358 353
rect 361 351 363 353
rect 366 351 368 353
rect 371 351 373 353
rect 376 351 378 353
rect 381 351 383 353
rect 386 351 388 353
rect 391 351 393 353
rect 396 351 398 353
rect 401 351 403 353
rect 406 351 408 353
rect 411 351 413 353
rect 416 351 418 353
rect 421 351 423 353
rect 426 351 428 353
rect 431 351 433 353
rect 436 351 438 353
rect 441 351 443 353
rect 446 351 448 353
rect 451 351 453 353
rect 456 351 458 353
rect 461 351 463 353
rect 466 351 468 353
rect 471 351 473 353
rect 476 351 478 353
rect 481 351 483 353
rect 486 351 488 353
rect 491 351 493 353
rect 496 351 498 353
rect 501 351 503 353
rect 506 351 508 353
rect 511 351 513 353
rect 516 351 518 353
rect 521 351 523 353
rect 526 351 528 353
rect 531 351 533 353
rect 536 351 538 353
rect 541 351 543 353
rect 546 351 548 353
rect 551 351 553 353
rect 556 351 558 353
rect 331 346 333 348
rect 336 346 338 348
rect 341 346 343 348
rect 346 346 348 348
rect 351 346 353 348
rect 356 346 358 348
rect 361 346 363 348
rect 366 346 368 348
rect 371 346 373 348
rect 376 346 378 348
rect 381 346 383 348
rect 386 346 388 348
rect 391 346 393 348
rect 396 346 398 348
rect 401 346 403 348
rect 406 346 408 348
rect 411 346 413 348
rect 416 346 418 348
rect 421 346 423 348
rect 426 346 428 348
rect 431 346 433 348
rect 436 346 438 348
rect 441 346 443 348
rect 446 346 448 348
rect 451 346 453 348
rect 456 346 458 348
rect 461 346 463 348
rect 466 346 468 348
rect 471 346 473 348
rect 476 346 478 348
rect 481 346 483 348
rect 486 346 488 348
rect 491 346 493 348
rect 496 346 498 348
rect 501 346 503 348
rect 506 346 508 348
rect 511 346 513 348
rect 516 346 518 348
rect 521 346 523 348
rect 526 346 528 348
rect 531 346 533 348
rect 536 346 538 348
rect 541 346 543 348
rect 546 346 548 348
rect 551 346 553 348
rect 556 346 558 348
rect 331 341 333 343
rect 336 341 338 343
rect 341 341 343 343
rect 346 341 348 343
rect 351 341 353 343
rect 356 341 358 343
rect 361 341 363 343
rect 366 341 368 343
rect 371 341 373 343
rect 376 341 378 343
rect 381 341 383 343
rect 386 341 388 343
rect 391 341 393 343
rect 396 341 398 343
rect 401 341 403 343
rect 406 341 408 343
rect 411 341 413 343
rect 416 341 418 343
rect 421 341 423 343
rect 426 341 428 343
rect 431 341 433 343
rect 436 341 438 343
rect 441 341 443 343
rect 446 341 448 343
rect 451 341 453 343
rect 456 341 458 343
rect 461 341 463 343
rect 466 341 468 343
rect 471 341 473 343
rect 476 341 478 343
rect 481 341 483 343
rect 486 341 488 343
rect 491 341 493 343
rect 496 341 498 343
rect 501 341 503 343
rect 506 341 508 343
rect 511 341 513 343
rect 516 341 518 343
rect 521 341 523 343
rect 526 341 528 343
rect 531 341 533 343
rect 536 341 538 343
rect 541 341 543 343
rect 546 341 548 343
rect 551 341 553 343
rect 556 341 558 343
rect 331 336 333 338
rect 336 336 338 338
rect 341 336 343 338
rect 346 336 348 338
rect 351 336 353 338
rect 356 336 358 338
rect 361 336 363 338
rect 366 336 368 338
rect 371 336 373 338
rect 376 336 378 338
rect 381 336 383 338
rect 386 336 388 338
rect 391 336 393 338
rect 396 336 398 338
rect 401 336 403 338
rect 406 336 408 338
rect 411 336 413 338
rect 416 336 418 338
rect 421 336 423 338
rect 426 336 428 338
rect 431 336 433 338
rect 436 336 438 338
rect 441 336 443 338
rect 446 336 448 338
rect 451 336 453 338
rect 456 336 458 338
rect 461 336 463 338
rect 466 336 468 338
rect 471 336 473 338
rect 476 336 478 338
rect 481 336 483 338
rect 486 336 488 338
rect 491 336 493 338
rect 496 336 498 338
rect 501 336 503 338
rect 506 336 508 338
rect 511 336 513 338
rect 516 336 518 338
rect 521 336 523 338
rect 526 336 528 338
rect 531 336 533 338
rect 536 336 538 338
rect 541 336 543 338
rect 546 336 548 338
rect 551 336 553 338
rect 556 336 558 338
rect 331 331 333 333
rect 336 331 338 333
rect 341 331 343 333
rect 346 331 348 333
rect 351 331 353 333
rect 356 331 358 333
rect 361 331 363 333
rect 366 331 368 333
rect 371 331 373 333
rect 376 331 378 333
rect 381 331 383 333
rect 386 331 388 333
rect 391 331 393 333
rect 396 331 398 333
rect 401 331 403 333
rect 406 331 408 333
rect 411 331 413 333
rect 416 331 418 333
rect 421 331 423 333
rect 426 331 428 333
rect 431 331 433 333
rect 436 331 438 333
rect 441 331 443 333
rect 446 331 448 333
rect 451 331 453 333
rect 456 331 458 333
rect 461 331 463 333
rect 466 331 468 333
rect 471 331 473 333
rect 476 331 478 333
rect 481 331 483 333
rect 486 331 488 333
rect 491 331 493 333
rect 496 331 498 333
rect 501 331 503 333
rect 506 331 508 333
rect 511 331 513 333
rect 516 331 518 333
rect 521 331 523 333
rect 526 331 528 333
rect 531 331 533 333
rect 536 331 538 333
rect 541 331 543 333
rect 546 331 548 333
rect 551 331 553 333
rect 556 331 558 333
rect 331 326 333 328
rect 336 326 338 328
rect 341 326 343 328
rect 346 326 348 328
rect 351 326 353 328
rect 356 326 358 328
rect 361 326 363 328
rect 366 326 368 328
rect 371 326 373 328
rect 376 326 378 328
rect 381 326 383 328
rect 386 326 388 328
rect 391 326 393 328
rect 396 326 398 328
rect 401 326 403 328
rect 406 326 408 328
rect 411 326 413 328
rect 416 326 418 328
rect 421 326 423 328
rect 426 326 428 328
rect 431 326 433 328
rect 436 326 438 328
rect 441 326 443 328
rect 446 326 448 328
rect 451 326 453 328
rect 456 326 458 328
rect 461 326 463 328
rect 466 326 468 328
rect 471 326 473 328
rect 476 326 478 328
rect 481 326 483 328
rect 486 326 488 328
rect 491 326 493 328
rect 496 326 498 328
rect 501 326 503 328
rect 506 326 508 328
rect 511 326 513 328
rect 516 326 518 328
rect 521 326 523 328
rect 526 326 528 328
rect 531 326 533 328
rect 536 326 538 328
rect 541 326 543 328
rect 546 326 548 328
rect 551 326 553 328
rect 556 326 558 328
rect 331 321 333 323
rect 336 321 338 323
rect 341 321 343 323
rect 346 321 348 323
rect 351 321 353 323
rect 356 321 358 323
rect 361 321 363 323
rect 366 321 368 323
rect 371 321 373 323
rect 376 321 378 323
rect 381 321 383 323
rect 386 321 388 323
rect 391 321 393 323
rect 396 321 398 323
rect 401 321 403 323
rect 406 321 408 323
rect 411 321 413 323
rect 416 321 418 323
rect 421 321 423 323
rect 426 321 428 323
rect 431 321 433 323
rect 436 321 438 323
rect 441 321 443 323
rect 446 321 448 323
rect 451 321 453 323
rect 456 321 458 323
rect 461 321 463 323
rect 466 321 468 323
rect 471 321 473 323
rect 476 321 478 323
rect 481 321 483 323
rect 486 321 488 323
rect 491 321 493 323
rect 496 321 498 323
rect 501 321 503 323
rect 506 321 508 323
rect 511 321 513 323
rect 516 321 518 323
rect 521 321 523 323
rect 526 321 528 323
rect 531 321 533 323
rect 536 321 538 323
rect 541 321 543 323
rect 546 321 548 323
rect 551 321 553 323
rect 556 321 558 323
rect 331 316 333 318
rect 336 316 338 318
rect 341 316 343 318
rect 346 316 348 318
rect 351 316 353 318
rect 356 316 358 318
rect 361 316 363 318
rect 366 316 368 318
rect 371 316 373 318
rect 376 316 378 318
rect 381 316 383 318
rect 386 316 388 318
rect 391 316 393 318
rect 396 316 398 318
rect 401 316 403 318
rect 406 316 408 318
rect 411 316 413 318
rect 416 316 418 318
rect 421 316 423 318
rect 426 316 428 318
rect 431 316 433 318
rect 436 316 438 318
rect 441 316 443 318
rect 446 316 448 318
rect 451 316 453 318
rect 456 316 458 318
rect 461 316 463 318
rect 466 316 468 318
rect 471 316 473 318
rect 476 316 478 318
rect 481 316 483 318
rect 486 316 488 318
rect 491 316 493 318
rect 496 316 498 318
rect 501 316 503 318
rect 506 316 508 318
rect 511 316 513 318
rect 516 316 518 318
rect 521 316 523 318
rect 526 316 528 318
rect 531 316 533 318
rect 536 316 538 318
rect 541 316 543 318
rect 546 316 548 318
rect 551 316 553 318
rect 556 316 558 318
rect 331 311 333 313
rect 336 311 338 313
rect 341 311 343 313
rect 346 311 348 313
rect 351 311 353 313
rect 356 311 358 313
rect 361 311 363 313
rect 366 311 368 313
rect 371 311 373 313
rect 376 311 378 313
rect 381 311 383 313
rect 386 311 388 313
rect 391 311 393 313
rect 396 311 398 313
rect 401 311 403 313
rect 406 311 408 313
rect 411 311 413 313
rect 416 311 418 313
rect 421 311 423 313
rect 426 311 428 313
rect 431 311 433 313
rect 436 311 438 313
rect 441 311 443 313
rect 446 311 448 313
rect 451 311 453 313
rect 456 311 458 313
rect 461 311 463 313
rect 466 311 468 313
rect 471 311 473 313
rect 476 311 478 313
rect 481 311 483 313
rect 486 311 488 313
rect 491 311 493 313
rect 496 311 498 313
rect 501 311 503 313
rect 506 311 508 313
rect 511 311 513 313
rect 516 311 518 313
rect 521 311 523 313
rect 526 311 528 313
rect 531 311 533 313
rect 536 311 538 313
rect 541 311 543 313
rect 546 311 548 313
rect 551 311 553 313
rect 556 311 558 313
rect 331 306 333 308
rect 336 306 338 308
rect 341 306 343 308
rect 346 306 348 308
rect 351 306 353 308
rect 356 306 358 308
rect 361 306 363 308
rect 366 306 368 308
rect 371 306 373 308
rect 376 306 378 308
rect 381 306 383 308
rect 386 306 388 308
rect 391 306 393 308
rect 396 306 398 308
rect 401 306 403 308
rect 406 306 408 308
rect 411 306 413 308
rect 416 306 418 308
rect 421 306 423 308
rect 426 306 428 308
rect 431 306 433 308
rect 436 306 438 308
rect 441 306 443 308
rect 446 306 448 308
rect 451 306 453 308
rect 456 306 458 308
rect 461 306 463 308
rect 466 306 468 308
rect 471 306 473 308
rect 476 306 478 308
rect 481 306 483 308
rect 486 306 488 308
rect 491 306 493 308
rect 496 306 498 308
rect 501 306 503 308
rect 506 306 508 308
rect 511 306 513 308
rect 516 306 518 308
rect 521 306 523 308
rect 526 306 528 308
rect 531 306 533 308
rect 536 306 538 308
rect 541 306 543 308
rect 546 306 548 308
rect 551 306 553 308
rect 556 306 558 308
rect 331 301 333 303
rect 336 301 338 303
rect 341 301 343 303
rect 346 301 348 303
rect 351 301 353 303
rect 356 301 358 303
rect 361 301 363 303
rect 366 301 368 303
rect 371 301 373 303
rect 376 301 378 303
rect 381 301 383 303
rect 386 301 388 303
rect 391 301 393 303
rect 396 301 398 303
rect 401 301 403 303
rect 406 301 408 303
rect 411 301 413 303
rect 416 301 418 303
rect 421 301 423 303
rect 426 301 428 303
rect 431 301 433 303
rect 436 301 438 303
rect 441 301 443 303
rect 446 301 448 303
rect 451 301 453 303
rect 456 301 458 303
rect 461 301 463 303
rect 466 301 468 303
rect 471 301 473 303
rect 476 301 478 303
rect 481 301 483 303
rect 486 301 488 303
rect 491 301 493 303
rect 496 301 498 303
rect 501 301 503 303
rect 506 301 508 303
rect 511 301 513 303
rect 516 301 518 303
rect 521 301 523 303
rect 526 301 528 303
rect 531 301 533 303
rect 536 301 538 303
rect 541 301 543 303
rect 546 301 548 303
rect 551 301 553 303
rect 556 301 558 303
rect 331 296 333 298
rect 336 296 338 298
rect 341 296 343 298
rect 346 296 348 298
rect 351 296 353 298
rect 356 296 358 298
rect 361 296 363 298
rect 366 296 368 298
rect 371 296 373 298
rect 376 296 378 298
rect 381 296 383 298
rect 386 296 388 298
rect 391 296 393 298
rect 396 296 398 298
rect 401 296 403 298
rect 406 296 408 298
rect 411 296 413 298
rect 416 296 418 298
rect 421 296 423 298
rect 426 296 428 298
rect 431 296 433 298
rect 436 296 438 298
rect 441 296 443 298
rect 446 296 448 298
rect 451 296 453 298
rect 456 296 458 298
rect 461 296 463 298
rect 466 296 468 298
rect 471 296 473 298
rect 476 296 478 298
rect 481 296 483 298
rect 486 296 488 298
rect 491 296 493 298
rect 496 296 498 298
rect 501 296 503 298
rect 506 296 508 298
rect 511 296 513 298
rect 516 296 518 298
rect 521 296 523 298
rect 526 296 528 298
rect 531 296 533 298
rect 536 296 538 298
rect 541 296 543 298
rect 546 296 548 298
rect 551 296 553 298
rect 556 296 558 298
rect 331 291 333 293
rect 336 291 338 293
rect 341 291 343 293
rect 346 291 348 293
rect 351 291 353 293
rect 356 291 358 293
rect 361 291 363 293
rect 366 291 368 293
rect 371 291 373 293
rect 376 291 378 293
rect 381 291 383 293
rect 386 291 388 293
rect 391 291 393 293
rect 396 291 398 293
rect 401 291 403 293
rect 406 291 408 293
rect 411 291 413 293
rect 416 291 418 293
rect 421 291 423 293
rect 426 291 428 293
rect 431 291 433 293
rect 436 291 438 293
rect 441 291 443 293
rect 446 291 448 293
rect 451 291 453 293
rect 456 291 458 293
rect 461 291 463 293
rect 466 291 468 293
rect 471 291 473 293
rect 476 291 478 293
rect 481 291 483 293
rect 486 291 488 293
rect 491 291 493 293
rect 496 291 498 293
rect 501 291 503 293
rect 506 291 508 293
rect 511 291 513 293
rect 516 291 518 293
rect 521 291 523 293
rect 526 291 528 293
rect 531 291 533 293
rect 536 291 538 293
rect 541 291 543 293
rect 546 291 548 293
rect 551 291 553 293
rect 556 291 558 293
rect 331 286 333 288
rect 336 286 338 288
rect 341 286 343 288
rect 346 286 348 288
rect 351 286 353 288
rect 356 286 358 288
rect 361 286 363 288
rect 366 286 368 288
rect 371 286 373 288
rect 376 286 378 288
rect 381 286 383 288
rect 386 286 388 288
rect 391 286 393 288
rect 396 286 398 288
rect 401 286 403 288
rect 406 286 408 288
rect 411 286 413 288
rect 416 286 418 288
rect 421 286 423 288
rect 426 286 428 288
rect 431 286 433 288
rect 436 286 438 288
rect 441 286 443 288
rect 446 286 448 288
rect 451 286 453 288
rect 456 286 458 288
rect 461 286 463 288
rect 466 286 468 288
rect 471 286 473 288
rect 476 286 478 288
rect 481 286 483 288
rect 486 286 488 288
rect 491 286 493 288
rect 496 286 498 288
rect 501 286 503 288
rect 506 286 508 288
rect 511 286 513 288
rect 516 286 518 288
rect 521 286 523 288
rect 526 286 528 288
rect 531 286 533 288
rect 536 286 538 288
rect 541 286 543 288
rect 546 286 548 288
rect 551 286 553 288
rect 556 286 558 288
rect 331 281 333 283
rect 336 281 338 283
rect 341 281 343 283
rect 346 281 348 283
rect 351 281 353 283
rect 356 281 358 283
rect 361 281 363 283
rect 366 281 368 283
rect 371 281 373 283
rect 376 281 378 283
rect 381 281 383 283
rect 386 281 388 283
rect 391 281 393 283
rect 396 281 398 283
rect 401 281 403 283
rect 406 281 408 283
rect 411 281 413 283
rect 416 281 418 283
rect 421 281 423 283
rect 426 281 428 283
rect 431 281 433 283
rect 436 281 438 283
rect 441 281 443 283
rect 446 281 448 283
rect 451 281 453 283
rect 456 281 458 283
rect 461 281 463 283
rect 466 281 468 283
rect 471 281 473 283
rect 476 281 478 283
rect 481 281 483 283
rect 486 281 488 283
rect 491 281 493 283
rect 496 281 498 283
rect 501 281 503 283
rect 506 281 508 283
rect 511 281 513 283
rect 516 281 518 283
rect 521 281 523 283
rect 526 281 528 283
rect 531 281 533 283
rect 536 281 538 283
rect 541 281 543 283
rect 546 281 548 283
rect 551 281 553 283
rect 556 281 558 283
rect 331 276 333 278
rect 336 276 338 278
rect 341 276 343 278
rect 346 276 348 278
rect 351 276 353 278
rect 356 276 358 278
rect 361 276 363 278
rect 366 276 368 278
rect 371 276 373 278
rect 376 276 378 278
rect 381 276 383 278
rect 386 276 388 278
rect 391 276 393 278
rect 396 276 398 278
rect 401 276 403 278
rect 406 276 408 278
rect 411 276 413 278
rect 416 276 418 278
rect 421 276 423 278
rect 426 276 428 278
rect 431 276 433 278
rect 436 276 438 278
rect 441 276 443 278
rect 446 276 448 278
rect 451 276 453 278
rect 456 276 458 278
rect 461 276 463 278
rect 466 276 468 278
rect 471 276 473 278
rect 476 276 478 278
rect 481 276 483 278
rect 486 276 488 278
rect 491 276 493 278
rect 496 276 498 278
rect 501 276 503 278
rect 506 276 508 278
rect 511 276 513 278
rect 516 276 518 278
rect 521 276 523 278
rect 526 276 528 278
rect 531 276 533 278
rect 536 276 538 278
rect 541 276 543 278
rect 546 276 548 278
rect 551 276 553 278
rect 556 276 558 278
rect 331 271 333 273
rect 336 271 338 273
rect 341 271 343 273
rect 346 271 348 273
rect 351 271 353 273
rect 356 271 358 273
rect 361 271 363 273
rect 366 271 368 273
rect 371 271 373 273
rect 376 271 378 273
rect 381 271 383 273
rect 386 271 388 273
rect 391 271 393 273
rect 396 271 398 273
rect 401 271 403 273
rect 406 271 408 273
rect 411 271 413 273
rect 416 271 418 273
rect 421 271 423 273
rect 426 271 428 273
rect 431 271 433 273
rect 436 271 438 273
rect 441 271 443 273
rect 446 271 448 273
rect 451 271 453 273
rect 456 271 458 273
rect 461 271 463 273
rect 466 271 468 273
rect 471 271 473 273
rect 476 271 478 273
rect 481 271 483 273
rect 486 271 488 273
rect 491 271 493 273
rect 496 271 498 273
rect 501 271 503 273
rect 506 271 508 273
rect 511 271 513 273
rect 516 271 518 273
rect 521 271 523 273
rect 526 271 528 273
rect 531 271 533 273
rect 536 271 538 273
rect 541 271 543 273
rect 546 271 548 273
rect 551 271 553 273
rect 556 271 558 273
rect 331 266 333 268
rect 336 266 338 268
rect 341 266 343 268
rect 346 266 348 268
rect 351 266 353 268
rect 356 266 358 268
rect 361 266 363 268
rect 366 266 368 268
rect 371 266 373 268
rect 376 266 378 268
rect 381 266 383 268
rect 386 266 388 268
rect 391 266 393 268
rect 396 266 398 268
rect 401 266 403 268
rect 406 266 408 268
rect 411 266 413 268
rect 416 266 418 268
rect 421 266 423 268
rect 426 266 428 268
rect 431 266 433 268
rect 436 266 438 268
rect 441 266 443 268
rect 446 266 448 268
rect 451 266 453 268
rect 456 266 458 268
rect 461 266 463 268
rect 466 266 468 268
rect 471 266 473 268
rect 476 266 478 268
rect 481 266 483 268
rect 486 266 488 268
rect 491 266 493 268
rect 496 266 498 268
rect 501 266 503 268
rect 506 266 508 268
rect 511 266 513 268
rect 516 266 518 268
rect 521 266 523 268
rect 526 266 528 268
rect 531 266 533 268
rect 536 266 538 268
rect 541 266 543 268
rect 546 266 548 268
rect 551 266 553 268
rect 556 266 558 268
rect 331 261 333 263
rect 336 261 338 263
rect 341 261 343 263
rect 346 261 348 263
rect 351 261 353 263
rect 356 261 358 263
rect 361 261 363 263
rect 366 261 368 263
rect 371 261 373 263
rect 376 261 378 263
rect 381 261 383 263
rect 386 261 388 263
rect 391 261 393 263
rect 396 261 398 263
rect 401 261 403 263
rect 406 261 408 263
rect 411 261 413 263
rect 416 261 418 263
rect 421 261 423 263
rect 426 261 428 263
rect 431 261 433 263
rect 436 261 438 263
rect 441 261 443 263
rect 446 261 448 263
rect 451 261 453 263
rect 456 261 458 263
rect 461 261 463 263
rect 466 261 468 263
rect 471 261 473 263
rect 476 261 478 263
rect 481 261 483 263
rect 486 261 488 263
rect 491 261 493 263
rect 496 261 498 263
rect 501 261 503 263
rect 506 261 508 263
rect 511 261 513 263
rect 516 261 518 263
rect 521 261 523 263
rect 526 261 528 263
rect 531 261 533 263
rect 536 261 538 263
rect 541 261 543 263
rect 546 261 548 263
rect 551 261 553 263
rect 556 261 558 263
rect 331 256 333 258
rect 336 256 338 258
rect 341 256 343 258
rect 346 256 348 258
rect 351 256 353 258
rect 356 256 358 258
rect 361 256 363 258
rect 366 256 368 258
rect 371 256 373 258
rect 376 256 378 258
rect 381 256 383 258
rect 386 256 388 258
rect 391 256 393 258
rect 396 256 398 258
rect 401 256 403 258
rect 406 256 408 258
rect 411 256 413 258
rect 416 256 418 258
rect 421 256 423 258
rect 426 256 428 258
rect 431 256 433 258
rect 436 256 438 258
rect 441 256 443 258
rect 446 256 448 258
rect 451 256 453 258
rect 456 256 458 258
rect 461 256 463 258
rect 466 256 468 258
rect 471 256 473 258
rect 476 256 478 258
rect 481 256 483 258
rect 486 256 488 258
rect 491 256 493 258
rect 496 256 498 258
rect 501 256 503 258
rect 506 256 508 258
rect 511 256 513 258
rect 516 256 518 258
rect 521 256 523 258
rect 526 256 528 258
rect 531 256 533 258
rect 536 256 538 258
rect 541 256 543 258
rect 546 256 548 258
rect 551 256 553 258
rect 556 256 558 258
rect 331 251 333 253
rect 336 251 338 253
rect 341 251 343 253
rect 346 251 348 253
rect 351 251 353 253
rect 356 251 358 253
rect 361 251 363 253
rect 366 251 368 253
rect 371 251 373 253
rect 376 251 378 253
rect 381 251 383 253
rect 386 251 388 253
rect 391 251 393 253
rect 396 251 398 253
rect 401 251 403 253
rect 406 251 408 253
rect 411 251 413 253
rect 416 251 418 253
rect 421 251 423 253
rect 426 251 428 253
rect 431 251 433 253
rect 436 251 438 253
rect 441 251 443 253
rect 446 251 448 253
rect 451 251 453 253
rect 456 251 458 253
rect 461 251 463 253
rect 466 251 468 253
rect 471 251 473 253
rect 476 251 478 253
rect 481 251 483 253
rect 486 251 488 253
rect 491 251 493 253
rect 496 251 498 253
rect 501 251 503 253
rect 506 251 508 253
rect 511 251 513 253
rect 516 251 518 253
rect 521 251 523 253
rect 526 251 528 253
rect 531 251 533 253
rect 536 251 538 253
rect 541 251 543 253
rect 546 251 548 253
rect 551 251 553 253
rect 556 251 558 253
rect 331 246 333 248
rect 336 246 338 248
rect 341 246 343 248
rect 346 246 348 248
rect 351 246 353 248
rect 356 246 358 248
rect 361 246 363 248
rect 366 246 368 248
rect 371 246 373 248
rect 376 246 378 248
rect 381 246 383 248
rect 386 246 388 248
rect 391 246 393 248
rect 396 246 398 248
rect 401 246 403 248
rect 406 246 408 248
rect 411 246 413 248
rect 416 246 418 248
rect 421 246 423 248
rect 426 246 428 248
rect 431 246 433 248
rect 436 246 438 248
rect 441 246 443 248
rect 446 246 448 248
rect 451 246 453 248
rect 456 246 458 248
rect 461 246 463 248
rect 466 246 468 248
rect 471 246 473 248
rect 476 246 478 248
rect 481 246 483 248
rect 486 246 488 248
rect 491 246 493 248
rect 496 246 498 248
rect 501 246 503 248
rect 506 246 508 248
rect 511 246 513 248
rect 516 246 518 248
rect 521 246 523 248
rect 526 246 528 248
rect 531 246 533 248
rect 536 246 538 248
rect 541 246 543 248
rect 546 246 548 248
rect 551 246 553 248
rect 556 246 558 248
rect 331 241 333 243
rect 336 241 338 243
rect 341 241 343 243
rect 346 241 348 243
rect 351 241 353 243
rect 356 241 358 243
rect 361 241 363 243
rect 366 241 368 243
rect 371 241 373 243
rect 376 241 378 243
rect 381 241 383 243
rect 386 241 388 243
rect 391 241 393 243
rect 396 241 398 243
rect 401 241 403 243
rect 406 241 408 243
rect 411 241 413 243
rect 416 241 418 243
rect 421 241 423 243
rect 426 241 428 243
rect 431 241 433 243
rect 436 241 438 243
rect 441 241 443 243
rect 446 241 448 243
rect 451 241 453 243
rect 456 241 458 243
rect 461 241 463 243
rect 466 241 468 243
rect 471 241 473 243
rect 476 241 478 243
rect 481 241 483 243
rect 486 241 488 243
rect 491 241 493 243
rect 496 241 498 243
rect 501 241 503 243
rect 506 241 508 243
rect 511 241 513 243
rect 516 241 518 243
rect 521 241 523 243
rect 526 241 528 243
rect 531 241 533 243
rect 536 241 538 243
rect 541 241 543 243
rect 546 241 548 243
rect 551 241 553 243
rect 556 241 558 243
rect 331 236 333 238
rect 336 236 338 238
rect 341 236 343 238
rect 346 236 348 238
rect 351 236 353 238
rect 356 236 358 238
rect 361 236 363 238
rect 366 236 368 238
rect 371 236 373 238
rect 376 236 378 238
rect 381 236 383 238
rect 386 236 388 238
rect 391 236 393 238
rect 396 236 398 238
rect 401 236 403 238
rect 406 236 408 238
rect 411 236 413 238
rect 416 236 418 238
rect 421 236 423 238
rect 426 236 428 238
rect 431 236 433 238
rect 436 236 438 238
rect 441 236 443 238
rect 446 236 448 238
rect 451 236 453 238
rect 456 236 458 238
rect 461 236 463 238
rect 466 236 468 238
rect 471 236 473 238
rect 476 236 478 238
rect 481 236 483 238
rect 486 236 488 238
rect 491 236 493 238
rect 496 236 498 238
rect 501 236 503 238
rect 506 236 508 238
rect 511 236 513 238
rect 516 236 518 238
rect 521 236 523 238
rect 526 236 528 238
rect 531 236 533 238
rect 536 236 538 238
rect 541 236 543 238
rect 546 236 548 238
rect 551 236 553 238
rect 556 236 558 238
rect 331 231 333 233
rect 336 231 338 233
rect 341 231 343 233
rect 346 231 348 233
rect 351 231 353 233
rect 356 231 358 233
rect 361 231 363 233
rect 366 231 368 233
rect 371 231 373 233
rect 376 231 378 233
rect 381 231 383 233
rect 386 231 388 233
rect 391 231 393 233
rect 396 231 398 233
rect 401 231 403 233
rect 406 231 408 233
rect 411 231 413 233
rect 416 231 418 233
rect 421 231 423 233
rect 426 231 428 233
rect 431 231 433 233
rect 436 231 438 233
rect 441 231 443 233
rect 446 231 448 233
rect 451 231 453 233
rect 456 231 458 233
rect 461 231 463 233
rect 466 231 468 233
rect 471 231 473 233
rect 476 231 478 233
rect 481 231 483 233
rect 486 231 488 233
rect 491 231 493 233
rect 496 231 498 233
rect 501 231 503 233
rect 506 231 508 233
rect 511 231 513 233
rect 516 231 518 233
rect 521 231 523 233
rect 526 231 528 233
rect 531 231 533 233
rect 536 231 538 233
rect 541 231 543 233
rect 546 231 548 233
rect 551 231 553 233
rect 556 231 558 233
rect 331 226 333 228
rect 336 226 338 228
rect 341 226 343 228
rect 346 226 348 228
rect 351 226 353 228
rect 356 226 358 228
rect 361 226 363 228
rect 366 226 368 228
rect 371 226 373 228
rect 376 226 378 228
rect 381 226 383 228
rect 386 226 388 228
rect 391 226 393 228
rect 396 226 398 228
rect 401 226 403 228
rect 406 226 408 228
rect 411 226 413 228
rect 416 226 418 228
rect 421 226 423 228
rect 426 226 428 228
rect 431 226 433 228
rect 436 226 438 228
rect 441 226 443 228
rect 446 226 448 228
rect 451 226 453 228
rect 456 226 458 228
rect 461 226 463 228
rect 466 226 468 228
rect 471 226 473 228
rect 476 226 478 228
rect 481 226 483 228
rect 486 226 488 228
rect 491 226 493 228
rect 496 226 498 228
rect 501 226 503 228
rect 506 226 508 228
rect 511 226 513 228
rect 516 226 518 228
rect 521 226 523 228
rect 526 226 528 228
rect 531 226 533 228
rect 536 226 538 228
rect 541 226 543 228
rect 546 226 548 228
rect 551 226 553 228
rect 556 226 558 228
rect 771 227 773 229
rect 776 227 778 229
rect 781 227 783 229
rect 786 227 788 229
rect 791 227 793 229
rect 796 227 798 229
rect 801 227 803 229
rect 806 227 808 229
rect 811 227 813 229
rect 816 227 818 229
rect 821 227 823 229
rect 826 227 828 229
rect 831 227 833 229
rect 836 227 838 229
rect 841 227 843 229
rect 846 227 848 229
rect 851 227 853 229
rect 856 227 858 229
rect 861 227 863 229
rect 866 227 868 229
rect 871 227 873 229
rect 876 227 878 229
rect 881 227 883 229
rect 886 227 888 229
rect 891 227 893 229
rect 896 227 898 229
rect 901 227 903 229
rect 906 227 908 229
rect 911 227 913 229
rect 916 227 918 229
rect 921 227 923 229
rect 926 227 928 229
rect 931 227 933 229
rect 936 227 938 229
rect 941 227 943 229
rect 946 227 948 229
rect 951 227 953 229
rect 956 227 958 229
rect 961 227 963 229
rect 966 227 968 229
rect 971 227 973 229
rect 976 227 978 229
rect 981 227 983 229
rect 986 227 988 229
rect 991 227 993 229
rect 996 227 998 229
rect 331 221 333 223
rect 336 221 338 223
rect 341 221 343 223
rect 346 221 348 223
rect 351 221 353 223
rect 356 221 358 223
rect 361 221 363 223
rect 366 221 368 223
rect 371 221 373 223
rect 376 221 378 223
rect 381 221 383 223
rect 386 221 388 223
rect 391 221 393 223
rect 396 221 398 223
rect 401 221 403 223
rect 406 221 408 223
rect 411 221 413 223
rect 416 221 418 223
rect 421 221 423 223
rect 426 221 428 223
rect 431 221 433 223
rect 436 221 438 223
rect 441 221 443 223
rect 446 221 448 223
rect 451 221 453 223
rect 456 221 458 223
rect 461 221 463 223
rect 466 221 468 223
rect 471 221 473 223
rect 476 221 478 223
rect 481 221 483 223
rect 486 221 488 223
rect 491 221 493 223
rect 496 221 498 223
rect 501 221 503 223
rect 506 221 508 223
rect 511 221 513 223
rect 516 221 518 223
rect 521 221 523 223
rect 526 221 528 223
rect 531 221 533 223
rect 536 221 538 223
rect 541 221 543 223
rect 546 221 548 223
rect 551 221 553 223
rect 556 221 558 223
rect 771 222 773 224
rect 776 222 778 224
rect 781 222 783 224
rect 786 222 788 224
rect 791 222 793 224
rect 796 222 798 224
rect 801 222 803 224
rect 806 222 808 224
rect 811 222 813 224
rect 816 222 818 224
rect 821 222 823 224
rect 826 222 828 224
rect 831 222 833 224
rect 836 222 838 224
rect 841 222 843 224
rect 846 222 848 224
rect 851 222 853 224
rect 856 222 858 224
rect 861 222 863 224
rect 866 222 868 224
rect 871 222 873 224
rect 876 222 878 224
rect 881 222 883 224
rect 886 222 888 224
rect 891 222 893 224
rect 896 222 898 224
rect 901 222 903 224
rect 906 222 908 224
rect 911 222 913 224
rect 916 222 918 224
rect 921 222 923 224
rect 926 222 928 224
rect 931 222 933 224
rect 936 222 938 224
rect 941 222 943 224
rect 946 222 948 224
rect 951 222 953 224
rect 956 222 958 224
rect 961 222 963 224
rect 966 222 968 224
rect 971 222 973 224
rect 976 222 978 224
rect 981 222 983 224
rect 986 222 988 224
rect 991 222 993 224
rect 996 222 998 224
rect 331 216 333 218
rect 336 216 338 218
rect 341 216 343 218
rect 346 216 348 218
rect 351 216 353 218
rect 356 216 358 218
rect 361 216 363 218
rect 366 216 368 218
rect 371 216 373 218
rect 376 216 378 218
rect 381 216 383 218
rect 386 216 388 218
rect 391 216 393 218
rect 396 216 398 218
rect 401 216 403 218
rect 406 216 408 218
rect 411 216 413 218
rect 416 216 418 218
rect 421 216 423 218
rect 426 216 428 218
rect 431 216 433 218
rect 436 216 438 218
rect 441 216 443 218
rect 446 216 448 218
rect 451 216 453 218
rect 456 216 458 218
rect 461 216 463 218
rect 466 216 468 218
rect 471 216 473 218
rect 476 216 478 218
rect 481 216 483 218
rect 486 216 488 218
rect 491 216 493 218
rect 496 216 498 218
rect 501 216 503 218
rect 506 216 508 218
rect 511 216 513 218
rect 516 216 518 218
rect 521 216 523 218
rect 526 216 528 218
rect 531 216 533 218
rect 536 216 538 218
rect 541 216 543 218
rect 546 216 548 218
rect 551 216 553 218
rect 556 216 558 218
rect 771 217 773 219
rect 776 217 778 219
rect 781 217 783 219
rect 786 217 788 219
rect 791 217 793 219
rect 796 217 798 219
rect 801 217 803 219
rect 806 217 808 219
rect 811 217 813 219
rect 816 217 818 219
rect 821 217 823 219
rect 826 217 828 219
rect 831 217 833 219
rect 836 217 838 219
rect 841 217 843 219
rect 846 217 848 219
rect 851 217 853 219
rect 856 217 858 219
rect 861 217 863 219
rect 866 217 868 219
rect 871 217 873 219
rect 876 217 878 219
rect 881 217 883 219
rect 886 217 888 219
rect 891 217 893 219
rect 896 217 898 219
rect 901 217 903 219
rect 906 217 908 219
rect 911 217 913 219
rect 916 217 918 219
rect 921 217 923 219
rect 926 217 928 219
rect 931 217 933 219
rect 936 217 938 219
rect 941 217 943 219
rect 946 217 948 219
rect 951 217 953 219
rect 956 217 958 219
rect 961 217 963 219
rect 966 217 968 219
rect 971 217 973 219
rect 976 217 978 219
rect 981 217 983 219
rect 986 217 988 219
rect 991 217 993 219
rect 996 217 998 219
rect 331 211 333 213
rect 336 211 338 213
rect 341 211 343 213
rect 346 211 348 213
rect 351 211 353 213
rect 356 211 358 213
rect 361 211 363 213
rect 366 211 368 213
rect 371 211 373 213
rect 376 211 378 213
rect 381 211 383 213
rect 386 211 388 213
rect 391 211 393 213
rect 396 211 398 213
rect 401 211 403 213
rect 406 211 408 213
rect 411 211 413 213
rect 416 211 418 213
rect 421 211 423 213
rect 426 211 428 213
rect 431 211 433 213
rect 436 211 438 213
rect 441 211 443 213
rect 446 211 448 213
rect 451 211 453 213
rect 456 211 458 213
rect 461 211 463 213
rect 466 211 468 213
rect 471 211 473 213
rect 476 211 478 213
rect 481 211 483 213
rect 486 211 488 213
rect 491 211 493 213
rect 496 211 498 213
rect 501 211 503 213
rect 506 211 508 213
rect 511 211 513 213
rect 516 211 518 213
rect 521 211 523 213
rect 526 211 528 213
rect 531 211 533 213
rect 536 211 538 213
rect 541 211 543 213
rect 546 211 548 213
rect 551 211 553 213
rect 556 211 558 213
rect 771 212 773 214
rect 776 212 778 214
rect 781 212 783 214
rect 786 212 788 214
rect 791 212 793 214
rect 796 212 798 214
rect 801 212 803 214
rect 806 212 808 214
rect 811 212 813 214
rect 816 212 818 214
rect 821 212 823 214
rect 826 212 828 214
rect 831 212 833 214
rect 836 212 838 214
rect 841 212 843 214
rect 846 212 848 214
rect 851 212 853 214
rect 856 212 858 214
rect 861 212 863 214
rect 866 212 868 214
rect 871 212 873 214
rect 876 212 878 214
rect 881 212 883 214
rect 886 212 888 214
rect 891 212 893 214
rect 896 212 898 214
rect 901 212 903 214
rect 906 212 908 214
rect 911 212 913 214
rect 916 212 918 214
rect 921 212 923 214
rect 926 212 928 214
rect 931 212 933 214
rect 936 212 938 214
rect 941 212 943 214
rect 946 212 948 214
rect 951 212 953 214
rect 956 212 958 214
rect 961 212 963 214
rect 966 212 968 214
rect 971 212 973 214
rect 976 212 978 214
rect 981 212 983 214
rect 986 212 988 214
rect 991 212 993 214
rect 996 212 998 214
rect 331 206 333 208
rect 336 206 338 208
rect 341 206 343 208
rect 346 206 348 208
rect 351 206 353 208
rect 356 206 358 208
rect 361 206 363 208
rect 366 206 368 208
rect 371 206 373 208
rect 376 206 378 208
rect 381 206 383 208
rect 386 206 388 208
rect 391 206 393 208
rect 396 206 398 208
rect 401 206 403 208
rect 406 206 408 208
rect 411 206 413 208
rect 416 206 418 208
rect 421 206 423 208
rect 426 206 428 208
rect 431 206 433 208
rect 436 206 438 208
rect 441 206 443 208
rect 446 206 448 208
rect 451 206 453 208
rect 456 206 458 208
rect 461 206 463 208
rect 466 206 468 208
rect 471 206 473 208
rect 476 206 478 208
rect 481 206 483 208
rect 486 206 488 208
rect 491 206 493 208
rect 496 206 498 208
rect 501 206 503 208
rect 506 206 508 208
rect 511 206 513 208
rect 516 206 518 208
rect 521 206 523 208
rect 526 206 528 208
rect 531 206 533 208
rect 536 206 538 208
rect 541 206 543 208
rect 546 206 548 208
rect 551 206 553 208
rect 556 206 558 208
rect 771 207 773 209
rect 776 207 778 209
rect 781 207 783 209
rect 786 207 788 209
rect 791 207 793 209
rect 796 207 798 209
rect 801 207 803 209
rect 806 207 808 209
rect 811 207 813 209
rect 816 207 818 209
rect 821 207 823 209
rect 826 207 828 209
rect 831 207 833 209
rect 836 207 838 209
rect 841 207 843 209
rect 846 207 848 209
rect 851 207 853 209
rect 856 207 858 209
rect 861 207 863 209
rect 866 207 868 209
rect 871 207 873 209
rect 876 207 878 209
rect 881 207 883 209
rect 886 207 888 209
rect 891 207 893 209
rect 896 207 898 209
rect 901 207 903 209
rect 906 207 908 209
rect 911 207 913 209
rect 916 207 918 209
rect 921 207 923 209
rect 926 207 928 209
rect 931 207 933 209
rect 936 207 938 209
rect 941 207 943 209
rect 946 207 948 209
rect 951 207 953 209
rect 956 207 958 209
rect 961 207 963 209
rect 966 207 968 209
rect 971 207 973 209
rect 976 207 978 209
rect 981 207 983 209
rect 986 207 988 209
rect 991 207 993 209
rect 996 207 998 209
rect 331 201 333 203
rect 336 201 338 203
rect 341 201 343 203
rect 346 201 348 203
rect 351 201 353 203
rect 356 201 358 203
rect 361 201 363 203
rect 366 201 368 203
rect 371 201 373 203
rect 376 201 378 203
rect 381 201 383 203
rect 386 201 388 203
rect 391 201 393 203
rect 396 201 398 203
rect 401 201 403 203
rect 406 201 408 203
rect 411 201 413 203
rect 416 201 418 203
rect 421 201 423 203
rect 426 201 428 203
rect 431 201 433 203
rect 436 201 438 203
rect 441 201 443 203
rect 446 201 448 203
rect 451 201 453 203
rect 456 201 458 203
rect 461 201 463 203
rect 466 201 468 203
rect 471 201 473 203
rect 476 201 478 203
rect 481 201 483 203
rect 486 201 488 203
rect 491 201 493 203
rect 496 201 498 203
rect 501 201 503 203
rect 506 201 508 203
rect 511 201 513 203
rect 516 201 518 203
rect 521 201 523 203
rect 526 201 528 203
rect 531 201 533 203
rect 536 201 538 203
rect 541 201 543 203
rect 546 201 548 203
rect 551 201 553 203
rect 556 201 558 203
rect 771 202 773 204
rect 776 202 778 204
rect 781 202 783 204
rect 786 202 788 204
rect 791 202 793 204
rect 796 202 798 204
rect 801 202 803 204
rect 806 202 808 204
rect 811 202 813 204
rect 816 202 818 204
rect 821 202 823 204
rect 826 202 828 204
rect 831 202 833 204
rect 836 202 838 204
rect 841 202 843 204
rect 846 202 848 204
rect 851 202 853 204
rect 856 202 858 204
rect 861 202 863 204
rect 866 202 868 204
rect 871 202 873 204
rect 876 202 878 204
rect 881 202 883 204
rect 886 202 888 204
rect 891 202 893 204
rect 896 202 898 204
rect 901 202 903 204
rect 906 202 908 204
rect 911 202 913 204
rect 916 202 918 204
rect 921 202 923 204
rect 926 202 928 204
rect 931 202 933 204
rect 936 202 938 204
rect 941 202 943 204
rect 946 202 948 204
rect 951 202 953 204
rect 956 202 958 204
rect 961 202 963 204
rect 966 202 968 204
rect 971 202 973 204
rect 976 202 978 204
rect 981 202 983 204
rect 986 202 988 204
rect 991 202 993 204
rect 996 202 998 204
rect 331 196 333 198
rect 336 196 338 198
rect 341 196 343 198
rect 346 196 348 198
rect 351 196 353 198
rect 356 196 358 198
rect 361 196 363 198
rect 366 196 368 198
rect 371 196 373 198
rect 376 196 378 198
rect 381 196 383 198
rect 386 196 388 198
rect 391 196 393 198
rect 396 196 398 198
rect 401 196 403 198
rect 406 196 408 198
rect 411 196 413 198
rect 416 196 418 198
rect 421 196 423 198
rect 426 196 428 198
rect 431 196 433 198
rect 436 196 438 198
rect 441 196 443 198
rect 446 196 448 198
rect 451 196 453 198
rect 456 196 458 198
rect 461 196 463 198
rect 466 196 468 198
rect 471 196 473 198
rect 476 196 478 198
rect 481 196 483 198
rect 486 196 488 198
rect 491 196 493 198
rect 496 196 498 198
rect 501 196 503 198
rect 506 196 508 198
rect 511 196 513 198
rect 516 196 518 198
rect 521 196 523 198
rect 526 196 528 198
rect 531 196 533 198
rect 536 196 538 198
rect 541 196 543 198
rect 546 196 548 198
rect 551 196 553 198
rect 556 196 558 198
rect 771 197 773 199
rect 776 197 778 199
rect 781 197 783 199
rect 786 197 788 199
rect 791 197 793 199
rect 796 197 798 199
rect 801 197 803 199
rect 806 197 808 199
rect 811 197 813 199
rect 816 197 818 199
rect 821 197 823 199
rect 826 197 828 199
rect 831 197 833 199
rect 836 197 838 199
rect 841 197 843 199
rect 846 197 848 199
rect 851 197 853 199
rect 856 197 858 199
rect 861 197 863 199
rect 866 197 868 199
rect 871 197 873 199
rect 876 197 878 199
rect 881 197 883 199
rect 886 197 888 199
rect 891 197 893 199
rect 896 197 898 199
rect 901 197 903 199
rect 906 197 908 199
rect 911 197 913 199
rect 916 197 918 199
rect 921 197 923 199
rect 926 197 928 199
rect 931 197 933 199
rect 936 197 938 199
rect 941 197 943 199
rect 946 197 948 199
rect 951 197 953 199
rect 956 197 958 199
rect 961 197 963 199
rect 966 197 968 199
rect 971 197 973 199
rect 976 197 978 199
rect 981 197 983 199
rect 986 197 988 199
rect 991 197 993 199
rect 996 197 998 199
rect 331 191 333 193
rect 336 191 338 193
rect 341 191 343 193
rect 346 191 348 193
rect 351 191 353 193
rect 356 191 358 193
rect 361 191 363 193
rect 366 191 368 193
rect 371 191 373 193
rect 376 191 378 193
rect 381 191 383 193
rect 386 191 388 193
rect 391 191 393 193
rect 396 191 398 193
rect 401 191 403 193
rect 406 191 408 193
rect 411 191 413 193
rect 416 191 418 193
rect 421 191 423 193
rect 426 191 428 193
rect 431 191 433 193
rect 436 191 438 193
rect 441 191 443 193
rect 446 191 448 193
rect 451 191 453 193
rect 456 191 458 193
rect 461 191 463 193
rect 466 191 468 193
rect 471 191 473 193
rect 476 191 478 193
rect 481 191 483 193
rect 486 191 488 193
rect 491 191 493 193
rect 496 191 498 193
rect 501 191 503 193
rect 506 191 508 193
rect 511 191 513 193
rect 516 191 518 193
rect 521 191 523 193
rect 526 191 528 193
rect 531 191 533 193
rect 536 191 538 193
rect 541 191 543 193
rect 546 191 548 193
rect 551 191 553 193
rect 556 191 558 193
rect 771 192 773 194
rect 776 192 778 194
rect 781 192 783 194
rect 786 192 788 194
rect 791 192 793 194
rect 796 192 798 194
rect 801 192 803 194
rect 806 192 808 194
rect 811 192 813 194
rect 816 192 818 194
rect 821 192 823 194
rect 826 192 828 194
rect 831 192 833 194
rect 836 192 838 194
rect 841 192 843 194
rect 846 192 848 194
rect 851 192 853 194
rect 856 192 858 194
rect 861 192 863 194
rect 866 192 868 194
rect 871 192 873 194
rect 876 192 878 194
rect 881 192 883 194
rect 886 192 888 194
rect 891 192 893 194
rect 896 192 898 194
rect 901 192 903 194
rect 906 192 908 194
rect 911 192 913 194
rect 916 192 918 194
rect 921 192 923 194
rect 926 192 928 194
rect 931 192 933 194
rect 936 192 938 194
rect 941 192 943 194
rect 946 192 948 194
rect 951 192 953 194
rect 956 192 958 194
rect 961 192 963 194
rect 966 192 968 194
rect 971 192 973 194
rect 976 192 978 194
rect 981 192 983 194
rect 986 192 988 194
rect 991 192 993 194
rect 996 192 998 194
rect 331 186 333 188
rect 336 186 338 188
rect 341 186 343 188
rect 346 186 348 188
rect 351 186 353 188
rect 356 186 358 188
rect 361 186 363 188
rect 366 186 368 188
rect 371 186 373 188
rect 376 186 378 188
rect 381 186 383 188
rect 386 186 388 188
rect 391 186 393 188
rect 396 186 398 188
rect 401 186 403 188
rect 406 186 408 188
rect 411 186 413 188
rect 416 186 418 188
rect 421 186 423 188
rect 426 186 428 188
rect 431 186 433 188
rect 436 186 438 188
rect 441 186 443 188
rect 446 186 448 188
rect 451 186 453 188
rect 456 186 458 188
rect 461 186 463 188
rect 466 186 468 188
rect 471 186 473 188
rect 476 186 478 188
rect 481 186 483 188
rect 486 186 488 188
rect 491 186 493 188
rect 496 186 498 188
rect 501 186 503 188
rect 506 186 508 188
rect 511 186 513 188
rect 516 186 518 188
rect 521 186 523 188
rect 526 186 528 188
rect 531 186 533 188
rect 536 186 538 188
rect 541 186 543 188
rect 546 186 548 188
rect 551 186 553 188
rect 556 186 558 188
rect 771 187 773 189
rect 776 187 778 189
rect 781 187 783 189
rect 786 187 788 189
rect 791 187 793 189
rect 796 187 798 189
rect 801 187 803 189
rect 806 187 808 189
rect 811 187 813 189
rect 816 187 818 189
rect 821 187 823 189
rect 826 187 828 189
rect 831 187 833 189
rect 836 187 838 189
rect 841 187 843 189
rect 846 187 848 189
rect 851 187 853 189
rect 856 187 858 189
rect 861 187 863 189
rect 866 187 868 189
rect 871 187 873 189
rect 876 187 878 189
rect 881 187 883 189
rect 886 187 888 189
rect 891 187 893 189
rect 896 187 898 189
rect 901 187 903 189
rect 906 187 908 189
rect 911 187 913 189
rect 916 187 918 189
rect 921 187 923 189
rect 926 187 928 189
rect 931 187 933 189
rect 936 187 938 189
rect 941 187 943 189
rect 946 187 948 189
rect 951 187 953 189
rect 956 187 958 189
rect 961 187 963 189
rect 966 187 968 189
rect 971 187 973 189
rect 976 187 978 189
rect 981 187 983 189
rect 986 187 988 189
rect 991 187 993 189
rect 996 187 998 189
rect 331 181 333 183
rect 336 181 338 183
rect 341 181 343 183
rect 346 181 348 183
rect 351 181 353 183
rect 356 181 358 183
rect 361 181 363 183
rect 366 181 368 183
rect 371 181 373 183
rect 376 181 378 183
rect 381 181 383 183
rect 386 181 388 183
rect 391 181 393 183
rect 396 181 398 183
rect 401 181 403 183
rect 406 181 408 183
rect 411 181 413 183
rect 416 181 418 183
rect 421 181 423 183
rect 426 181 428 183
rect 431 181 433 183
rect 436 181 438 183
rect 441 181 443 183
rect 446 181 448 183
rect 451 181 453 183
rect 456 181 458 183
rect 461 181 463 183
rect 466 181 468 183
rect 471 181 473 183
rect 476 181 478 183
rect 481 181 483 183
rect 486 181 488 183
rect 491 181 493 183
rect 496 181 498 183
rect 501 181 503 183
rect 506 181 508 183
rect 511 181 513 183
rect 516 181 518 183
rect 521 181 523 183
rect 526 181 528 183
rect 531 181 533 183
rect 536 181 538 183
rect 541 181 543 183
rect 546 181 548 183
rect 551 181 553 183
rect 556 181 558 183
rect 771 182 773 184
rect 776 182 778 184
rect 781 182 783 184
rect 786 182 788 184
rect 791 182 793 184
rect 796 182 798 184
rect 801 182 803 184
rect 806 182 808 184
rect 811 182 813 184
rect 816 182 818 184
rect 821 182 823 184
rect 826 182 828 184
rect 831 182 833 184
rect 836 182 838 184
rect 841 182 843 184
rect 846 182 848 184
rect 851 182 853 184
rect 856 182 858 184
rect 861 182 863 184
rect 866 182 868 184
rect 871 182 873 184
rect 876 182 878 184
rect 881 182 883 184
rect 886 182 888 184
rect 891 182 893 184
rect 896 182 898 184
rect 901 182 903 184
rect 906 182 908 184
rect 911 182 913 184
rect 916 182 918 184
rect 921 182 923 184
rect 926 182 928 184
rect 931 182 933 184
rect 936 182 938 184
rect 941 182 943 184
rect 946 182 948 184
rect 951 182 953 184
rect 956 182 958 184
rect 961 182 963 184
rect 966 182 968 184
rect 971 182 973 184
rect 976 182 978 184
rect 981 182 983 184
rect 986 182 988 184
rect 991 182 993 184
rect 996 182 998 184
rect 331 176 333 178
rect 336 176 338 178
rect 341 176 343 178
rect 346 176 348 178
rect 351 176 353 178
rect 356 176 358 178
rect 361 176 363 178
rect 366 176 368 178
rect 371 176 373 178
rect 376 176 378 178
rect 381 176 383 178
rect 386 176 388 178
rect 391 176 393 178
rect 396 176 398 178
rect 401 176 403 178
rect 406 176 408 178
rect 411 176 413 178
rect 416 176 418 178
rect 421 176 423 178
rect 426 176 428 178
rect 431 176 433 178
rect 436 176 438 178
rect 441 176 443 178
rect 446 176 448 178
rect 451 176 453 178
rect 456 176 458 178
rect 461 176 463 178
rect 466 176 468 178
rect 471 176 473 178
rect 476 176 478 178
rect 481 176 483 178
rect 486 176 488 178
rect 491 176 493 178
rect 496 176 498 178
rect 501 176 503 178
rect 506 176 508 178
rect 511 176 513 178
rect 516 176 518 178
rect 521 176 523 178
rect 526 176 528 178
rect 531 176 533 178
rect 536 176 538 178
rect 541 176 543 178
rect 546 176 548 178
rect 551 176 553 178
rect 556 176 558 178
rect 771 177 773 179
rect 776 177 778 179
rect 781 177 783 179
rect 786 177 788 179
rect 791 177 793 179
rect 796 177 798 179
rect 801 177 803 179
rect 806 177 808 179
rect 811 177 813 179
rect 816 177 818 179
rect 821 177 823 179
rect 826 177 828 179
rect 831 177 833 179
rect 836 177 838 179
rect 841 177 843 179
rect 846 177 848 179
rect 851 177 853 179
rect 856 177 858 179
rect 861 177 863 179
rect 866 177 868 179
rect 871 177 873 179
rect 876 177 878 179
rect 881 177 883 179
rect 886 177 888 179
rect 891 177 893 179
rect 896 177 898 179
rect 901 177 903 179
rect 906 177 908 179
rect 911 177 913 179
rect 916 177 918 179
rect 921 177 923 179
rect 926 177 928 179
rect 931 177 933 179
rect 936 177 938 179
rect 941 177 943 179
rect 946 177 948 179
rect 951 177 953 179
rect 956 177 958 179
rect 961 177 963 179
rect 966 177 968 179
rect 971 177 973 179
rect 976 177 978 179
rect 981 177 983 179
rect 986 177 988 179
rect 991 177 993 179
rect 996 177 998 179
rect 331 171 333 173
rect 336 171 338 173
rect 341 171 343 173
rect 346 171 348 173
rect 351 171 353 173
rect 356 171 358 173
rect 361 171 363 173
rect 366 171 368 173
rect 371 171 373 173
rect 376 171 378 173
rect 381 171 383 173
rect 386 171 388 173
rect 391 171 393 173
rect 396 171 398 173
rect 401 171 403 173
rect 406 171 408 173
rect 411 171 413 173
rect 416 171 418 173
rect 421 171 423 173
rect 426 171 428 173
rect 431 171 433 173
rect 436 171 438 173
rect 441 171 443 173
rect 446 171 448 173
rect 451 171 453 173
rect 456 171 458 173
rect 461 171 463 173
rect 466 171 468 173
rect 471 171 473 173
rect 476 171 478 173
rect 481 171 483 173
rect 486 171 488 173
rect 491 171 493 173
rect 496 171 498 173
rect 501 171 503 173
rect 506 171 508 173
rect 511 171 513 173
rect 516 171 518 173
rect 521 171 523 173
rect 526 171 528 173
rect 531 171 533 173
rect 536 171 538 173
rect 541 171 543 173
rect 546 171 548 173
rect 551 171 553 173
rect 556 171 558 173
rect 771 172 773 174
rect 776 172 778 174
rect 781 172 783 174
rect 786 172 788 174
rect 791 172 793 174
rect 796 172 798 174
rect 801 172 803 174
rect 806 172 808 174
rect 811 172 813 174
rect 816 172 818 174
rect 821 172 823 174
rect 826 172 828 174
rect 831 172 833 174
rect 836 172 838 174
rect 841 172 843 174
rect 846 172 848 174
rect 851 172 853 174
rect 856 172 858 174
rect 861 172 863 174
rect 866 172 868 174
rect 871 172 873 174
rect 876 172 878 174
rect 881 172 883 174
rect 886 172 888 174
rect 891 172 893 174
rect 896 172 898 174
rect 901 172 903 174
rect 906 172 908 174
rect 911 172 913 174
rect 916 172 918 174
rect 921 172 923 174
rect 926 172 928 174
rect 931 172 933 174
rect 936 172 938 174
rect 941 172 943 174
rect 946 172 948 174
rect 951 172 953 174
rect 956 172 958 174
rect 961 172 963 174
rect 966 172 968 174
rect 971 172 973 174
rect 976 172 978 174
rect 981 172 983 174
rect 986 172 988 174
rect 991 172 993 174
rect 996 172 998 174
rect 331 166 333 168
rect 336 166 338 168
rect 341 166 343 168
rect 346 166 348 168
rect 351 166 353 168
rect 356 166 358 168
rect 361 166 363 168
rect 366 166 368 168
rect 371 166 373 168
rect 376 166 378 168
rect 381 166 383 168
rect 386 166 388 168
rect 391 166 393 168
rect 396 166 398 168
rect 401 166 403 168
rect 406 166 408 168
rect 411 166 413 168
rect 416 166 418 168
rect 421 166 423 168
rect 426 166 428 168
rect 431 166 433 168
rect 436 166 438 168
rect 441 166 443 168
rect 446 166 448 168
rect 451 166 453 168
rect 456 166 458 168
rect 461 166 463 168
rect 466 166 468 168
rect 471 166 473 168
rect 476 166 478 168
rect 481 166 483 168
rect 486 166 488 168
rect 491 166 493 168
rect 496 166 498 168
rect 501 166 503 168
rect 506 166 508 168
rect 511 166 513 168
rect 516 166 518 168
rect 521 166 523 168
rect 526 166 528 168
rect 531 166 533 168
rect 536 166 538 168
rect 541 166 543 168
rect 546 166 548 168
rect 551 166 553 168
rect 556 166 558 168
rect 771 167 773 169
rect 776 167 778 169
rect 781 167 783 169
rect 786 167 788 169
rect 791 167 793 169
rect 796 167 798 169
rect 801 167 803 169
rect 806 167 808 169
rect 811 167 813 169
rect 816 167 818 169
rect 821 167 823 169
rect 826 167 828 169
rect 831 167 833 169
rect 836 167 838 169
rect 841 167 843 169
rect 846 167 848 169
rect 851 167 853 169
rect 856 167 858 169
rect 861 167 863 169
rect 866 167 868 169
rect 871 167 873 169
rect 876 167 878 169
rect 881 167 883 169
rect 886 167 888 169
rect 891 167 893 169
rect 896 167 898 169
rect 901 167 903 169
rect 906 167 908 169
rect 911 167 913 169
rect 916 167 918 169
rect 921 167 923 169
rect 926 167 928 169
rect 931 167 933 169
rect 936 167 938 169
rect 941 167 943 169
rect 946 167 948 169
rect 951 167 953 169
rect 956 167 958 169
rect 961 167 963 169
rect 966 167 968 169
rect 971 167 973 169
rect 976 167 978 169
rect 981 167 983 169
rect 986 167 988 169
rect 991 167 993 169
rect 996 167 998 169
rect 331 161 333 163
rect 336 161 338 163
rect 341 161 343 163
rect 346 161 348 163
rect 351 161 353 163
rect 356 161 358 163
rect 361 161 363 163
rect 366 161 368 163
rect 371 161 373 163
rect 376 161 378 163
rect 381 161 383 163
rect 386 161 388 163
rect 391 161 393 163
rect 396 161 398 163
rect 401 161 403 163
rect 406 161 408 163
rect 411 161 413 163
rect 416 161 418 163
rect 421 161 423 163
rect 426 161 428 163
rect 431 161 433 163
rect 436 161 438 163
rect 441 161 443 163
rect 446 161 448 163
rect 451 161 453 163
rect 456 161 458 163
rect 461 161 463 163
rect 466 161 468 163
rect 471 161 473 163
rect 476 161 478 163
rect 481 161 483 163
rect 486 161 488 163
rect 491 161 493 163
rect 496 161 498 163
rect 501 161 503 163
rect 506 161 508 163
rect 511 161 513 163
rect 516 161 518 163
rect 521 161 523 163
rect 526 161 528 163
rect 531 161 533 163
rect 536 161 538 163
rect 541 161 543 163
rect 546 161 548 163
rect 551 161 553 163
rect 556 161 558 163
rect 771 162 773 164
rect 776 162 778 164
rect 781 162 783 164
rect 786 162 788 164
rect 791 162 793 164
rect 796 162 798 164
rect 801 162 803 164
rect 806 162 808 164
rect 811 162 813 164
rect 816 162 818 164
rect 821 162 823 164
rect 826 162 828 164
rect 831 162 833 164
rect 836 162 838 164
rect 841 162 843 164
rect 846 162 848 164
rect 851 162 853 164
rect 856 162 858 164
rect 861 162 863 164
rect 866 162 868 164
rect 871 162 873 164
rect 876 162 878 164
rect 881 162 883 164
rect 886 162 888 164
rect 891 162 893 164
rect 896 162 898 164
rect 901 162 903 164
rect 906 162 908 164
rect 911 162 913 164
rect 916 162 918 164
rect 921 162 923 164
rect 926 162 928 164
rect 931 162 933 164
rect 936 162 938 164
rect 941 162 943 164
rect 946 162 948 164
rect 951 162 953 164
rect 956 162 958 164
rect 961 162 963 164
rect 966 162 968 164
rect 971 162 973 164
rect 976 162 978 164
rect 981 162 983 164
rect 986 162 988 164
rect 991 162 993 164
rect 996 162 998 164
rect 331 156 333 158
rect 336 156 338 158
rect 341 156 343 158
rect 346 156 348 158
rect 351 156 353 158
rect 356 156 358 158
rect 361 156 363 158
rect 366 156 368 158
rect 371 156 373 158
rect 376 156 378 158
rect 381 156 383 158
rect 386 156 388 158
rect 391 156 393 158
rect 396 156 398 158
rect 401 156 403 158
rect 406 156 408 158
rect 411 156 413 158
rect 416 156 418 158
rect 421 156 423 158
rect 426 156 428 158
rect 431 156 433 158
rect 436 156 438 158
rect 441 156 443 158
rect 446 156 448 158
rect 451 156 453 158
rect 456 156 458 158
rect 461 156 463 158
rect 466 156 468 158
rect 471 156 473 158
rect 476 156 478 158
rect 481 156 483 158
rect 486 156 488 158
rect 491 156 493 158
rect 496 156 498 158
rect 501 156 503 158
rect 506 156 508 158
rect 511 156 513 158
rect 516 156 518 158
rect 521 156 523 158
rect 526 156 528 158
rect 531 156 533 158
rect 536 156 538 158
rect 541 156 543 158
rect 546 156 548 158
rect 551 156 553 158
rect 556 156 558 158
rect 771 157 773 159
rect 776 157 778 159
rect 781 157 783 159
rect 786 157 788 159
rect 791 157 793 159
rect 796 157 798 159
rect 801 157 803 159
rect 806 157 808 159
rect 811 157 813 159
rect 816 157 818 159
rect 821 157 823 159
rect 826 157 828 159
rect 831 157 833 159
rect 836 157 838 159
rect 841 157 843 159
rect 846 157 848 159
rect 851 157 853 159
rect 856 157 858 159
rect 861 157 863 159
rect 866 157 868 159
rect 871 157 873 159
rect 876 157 878 159
rect 881 157 883 159
rect 886 157 888 159
rect 891 157 893 159
rect 896 157 898 159
rect 901 157 903 159
rect 906 157 908 159
rect 911 157 913 159
rect 916 157 918 159
rect 921 157 923 159
rect 926 157 928 159
rect 931 157 933 159
rect 936 157 938 159
rect 941 157 943 159
rect 946 157 948 159
rect 951 157 953 159
rect 956 157 958 159
rect 961 157 963 159
rect 966 157 968 159
rect 971 157 973 159
rect 976 157 978 159
rect 981 157 983 159
rect 986 157 988 159
rect 991 157 993 159
rect 996 157 998 159
rect 331 151 333 153
rect 336 151 338 153
rect 341 151 343 153
rect 346 151 348 153
rect 351 151 353 153
rect 356 151 358 153
rect 361 151 363 153
rect 366 151 368 153
rect 371 151 373 153
rect 376 151 378 153
rect 381 151 383 153
rect 386 151 388 153
rect 391 151 393 153
rect 396 151 398 153
rect 401 151 403 153
rect 406 151 408 153
rect 411 151 413 153
rect 416 151 418 153
rect 421 151 423 153
rect 426 151 428 153
rect 431 151 433 153
rect 436 151 438 153
rect 441 151 443 153
rect 446 151 448 153
rect 451 151 453 153
rect 456 151 458 153
rect 461 151 463 153
rect 466 151 468 153
rect 471 151 473 153
rect 476 151 478 153
rect 481 151 483 153
rect 486 151 488 153
rect 491 151 493 153
rect 496 151 498 153
rect 501 151 503 153
rect 506 151 508 153
rect 511 151 513 153
rect 516 151 518 153
rect 521 151 523 153
rect 526 151 528 153
rect 531 151 533 153
rect 536 151 538 153
rect 541 151 543 153
rect 546 151 548 153
rect 551 151 553 153
rect 556 151 558 153
rect 771 152 773 154
rect 776 152 778 154
rect 781 152 783 154
rect 786 152 788 154
rect 791 152 793 154
rect 796 152 798 154
rect 801 152 803 154
rect 806 152 808 154
rect 811 152 813 154
rect 816 152 818 154
rect 821 152 823 154
rect 826 152 828 154
rect 831 152 833 154
rect 836 152 838 154
rect 841 152 843 154
rect 846 152 848 154
rect 851 152 853 154
rect 856 152 858 154
rect 861 152 863 154
rect 866 152 868 154
rect 871 152 873 154
rect 876 152 878 154
rect 881 152 883 154
rect 886 152 888 154
rect 891 152 893 154
rect 896 152 898 154
rect 901 152 903 154
rect 906 152 908 154
rect 911 152 913 154
rect 916 152 918 154
rect 921 152 923 154
rect 926 152 928 154
rect 931 152 933 154
rect 936 152 938 154
rect 941 152 943 154
rect 946 152 948 154
rect 951 152 953 154
rect 956 152 958 154
rect 961 152 963 154
rect 966 152 968 154
rect 971 152 973 154
rect 976 152 978 154
rect 981 152 983 154
rect 986 152 988 154
rect 991 152 993 154
rect 996 152 998 154
rect 331 146 333 148
rect 336 146 338 148
rect 341 146 343 148
rect 346 146 348 148
rect 351 146 353 148
rect 356 146 358 148
rect 361 146 363 148
rect 366 146 368 148
rect 371 146 373 148
rect 376 146 378 148
rect 381 146 383 148
rect 386 146 388 148
rect 391 146 393 148
rect 396 146 398 148
rect 401 146 403 148
rect 406 146 408 148
rect 411 146 413 148
rect 416 146 418 148
rect 421 146 423 148
rect 426 146 428 148
rect 431 146 433 148
rect 436 146 438 148
rect 441 146 443 148
rect 446 146 448 148
rect 451 146 453 148
rect 456 146 458 148
rect 461 146 463 148
rect 466 146 468 148
rect 471 146 473 148
rect 476 146 478 148
rect 481 146 483 148
rect 486 146 488 148
rect 491 146 493 148
rect 496 146 498 148
rect 501 146 503 148
rect 506 146 508 148
rect 511 146 513 148
rect 516 146 518 148
rect 521 146 523 148
rect 526 146 528 148
rect 531 146 533 148
rect 536 146 538 148
rect 541 146 543 148
rect 546 146 548 148
rect 551 146 553 148
rect 556 146 558 148
rect 771 147 773 149
rect 776 147 778 149
rect 781 147 783 149
rect 786 147 788 149
rect 791 147 793 149
rect 796 147 798 149
rect 801 147 803 149
rect 806 147 808 149
rect 811 147 813 149
rect 816 147 818 149
rect 821 147 823 149
rect 826 147 828 149
rect 831 147 833 149
rect 836 147 838 149
rect 841 147 843 149
rect 846 147 848 149
rect 851 147 853 149
rect 856 147 858 149
rect 861 147 863 149
rect 866 147 868 149
rect 871 147 873 149
rect 876 147 878 149
rect 881 147 883 149
rect 886 147 888 149
rect 891 147 893 149
rect 896 147 898 149
rect 901 147 903 149
rect 906 147 908 149
rect 911 147 913 149
rect 916 147 918 149
rect 921 147 923 149
rect 926 147 928 149
rect 931 147 933 149
rect 936 147 938 149
rect 941 147 943 149
rect 946 147 948 149
rect 951 147 953 149
rect 956 147 958 149
rect 961 147 963 149
rect 966 147 968 149
rect 971 147 973 149
rect 976 147 978 149
rect 981 147 983 149
rect 986 147 988 149
rect 991 147 993 149
rect 996 147 998 149
rect 331 141 333 143
rect 336 141 338 143
rect 341 141 343 143
rect 346 141 348 143
rect 351 141 353 143
rect 356 141 358 143
rect 361 141 363 143
rect 366 141 368 143
rect 371 141 373 143
rect 376 141 378 143
rect 381 141 383 143
rect 386 141 388 143
rect 391 141 393 143
rect 396 141 398 143
rect 401 141 403 143
rect 406 141 408 143
rect 411 141 413 143
rect 416 141 418 143
rect 421 141 423 143
rect 426 141 428 143
rect 431 141 433 143
rect 436 141 438 143
rect 441 141 443 143
rect 446 141 448 143
rect 451 141 453 143
rect 456 141 458 143
rect 461 141 463 143
rect 466 141 468 143
rect 471 141 473 143
rect 476 141 478 143
rect 481 141 483 143
rect 486 141 488 143
rect 491 141 493 143
rect 496 141 498 143
rect 501 141 503 143
rect 506 141 508 143
rect 511 141 513 143
rect 516 141 518 143
rect 521 141 523 143
rect 526 141 528 143
rect 531 141 533 143
rect 536 141 538 143
rect 541 141 543 143
rect 546 141 548 143
rect 551 141 553 143
rect 556 141 558 143
rect 771 142 773 144
rect 776 142 778 144
rect 781 142 783 144
rect 786 142 788 144
rect 791 142 793 144
rect 796 142 798 144
rect 801 142 803 144
rect 806 142 808 144
rect 811 142 813 144
rect 816 142 818 144
rect 821 142 823 144
rect 826 142 828 144
rect 831 142 833 144
rect 836 142 838 144
rect 841 142 843 144
rect 846 142 848 144
rect 851 142 853 144
rect 856 142 858 144
rect 861 142 863 144
rect 866 142 868 144
rect 871 142 873 144
rect 876 142 878 144
rect 881 142 883 144
rect 886 142 888 144
rect 891 142 893 144
rect 896 142 898 144
rect 901 142 903 144
rect 906 142 908 144
rect 911 142 913 144
rect 916 142 918 144
rect 921 142 923 144
rect 926 142 928 144
rect 931 142 933 144
rect 936 142 938 144
rect 941 142 943 144
rect 946 142 948 144
rect 951 142 953 144
rect 956 142 958 144
rect 961 142 963 144
rect 966 142 968 144
rect 971 142 973 144
rect 976 142 978 144
rect 981 142 983 144
rect 986 142 988 144
rect 991 142 993 144
rect 996 142 998 144
rect 331 136 333 138
rect 336 136 338 138
rect 341 136 343 138
rect 346 136 348 138
rect 351 136 353 138
rect 356 136 358 138
rect 361 136 363 138
rect 366 136 368 138
rect 371 136 373 138
rect 376 136 378 138
rect 381 136 383 138
rect 386 136 388 138
rect 391 136 393 138
rect 396 136 398 138
rect 401 136 403 138
rect 406 136 408 138
rect 411 136 413 138
rect 416 136 418 138
rect 421 136 423 138
rect 426 136 428 138
rect 431 136 433 138
rect 436 136 438 138
rect 441 136 443 138
rect 446 136 448 138
rect 451 136 453 138
rect 456 136 458 138
rect 461 136 463 138
rect 466 136 468 138
rect 471 136 473 138
rect 476 136 478 138
rect 481 136 483 138
rect 486 136 488 138
rect 491 136 493 138
rect 496 136 498 138
rect 501 136 503 138
rect 506 136 508 138
rect 511 136 513 138
rect 516 136 518 138
rect 521 136 523 138
rect 526 136 528 138
rect 531 136 533 138
rect 536 136 538 138
rect 541 136 543 138
rect 546 136 548 138
rect 551 136 553 138
rect 556 136 558 138
rect 771 137 773 139
rect 776 137 778 139
rect 781 137 783 139
rect 786 137 788 139
rect 791 137 793 139
rect 796 137 798 139
rect 801 137 803 139
rect 806 137 808 139
rect 811 137 813 139
rect 816 137 818 139
rect 821 137 823 139
rect 826 137 828 139
rect 831 137 833 139
rect 836 137 838 139
rect 841 137 843 139
rect 846 137 848 139
rect 851 137 853 139
rect 856 137 858 139
rect 861 137 863 139
rect 866 137 868 139
rect 871 137 873 139
rect 876 137 878 139
rect 881 137 883 139
rect 886 137 888 139
rect 891 137 893 139
rect 896 137 898 139
rect 901 137 903 139
rect 906 137 908 139
rect 911 137 913 139
rect 916 137 918 139
rect 921 137 923 139
rect 926 137 928 139
rect 931 137 933 139
rect 936 137 938 139
rect 941 137 943 139
rect 946 137 948 139
rect 951 137 953 139
rect 956 137 958 139
rect 961 137 963 139
rect 966 137 968 139
rect 971 137 973 139
rect 976 137 978 139
rect 981 137 983 139
rect 986 137 988 139
rect 991 137 993 139
rect 996 137 998 139
rect 331 131 333 133
rect 336 131 338 133
rect 341 131 343 133
rect 346 131 348 133
rect 351 131 353 133
rect 356 131 358 133
rect 361 131 363 133
rect 366 131 368 133
rect 371 131 373 133
rect 376 131 378 133
rect 381 131 383 133
rect 386 131 388 133
rect 391 131 393 133
rect 396 131 398 133
rect 401 131 403 133
rect 406 131 408 133
rect 411 131 413 133
rect 416 131 418 133
rect 421 131 423 133
rect 426 131 428 133
rect 431 131 433 133
rect 436 131 438 133
rect 441 131 443 133
rect 446 131 448 133
rect 451 131 453 133
rect 456 131 458 133
rect 461 131 463 133
rect 466 131 468 133
rect 471 131 473 133
rect 476 131 478 133
rect 481 131 483 133
rect 486 131 488 133
rect 491 131 493 133
rect 496 131 498 133
rect 501 131 503 133
rect 506 131 508 133
rect 511 131 513 133
rect 516 131 518 133
rect 521 131 523 133
rect 526 131 528 133
rect 531 131 533 133
rect 536 131 538 133
rect 541 131 543 133
rect 546 131 548 133
rect 551 131 553 133
rect 556 131 558 133
rect 771 132 773 134
rect 776 132 778 134
rect 781 132 783 134
rect 786 132 788 134
rect 791 132 793 134
rect 796 132 798 134
rect 801 132 803 134
rect 806 132 808 134
rect 811 132 813 134
rect 816 132 818 134
rect 821 132 823 134
rect 826 132 828 134
rect 831 132 833 134
rect 836 132 838 134
rect 841 132 843 134
rect 846 132 848 134
rect 851 132 853 134
rect 856 132 858 134
rect 861 132 863 134
rect 866 132 868 134
rect 871 132 873 134
rect 876 132 878 134
rect 881 132 883 134
rect 886 132 888 134
rect 891 132 893 134
rect 896 132 898 134
rect 901 132 903 134
rect 906 132 908 134
rect 911 132 913 134
rect 916 132 918 134
rect 921 132 923 134
rect 926 132 928 134
rect 931 132 933 134
rect 936 132 938 134
rect 941 132 943 134
rect 946 132 948 134
rect 951 132 953 134
rect 956 132 958 134
rect 961 132 963 134
rect 966 132 968 134
rect 971 132 973 134
rect 976 132 978 134
rect 981 132 983 134
rect 986 132 988 134
rect 991 132 993 134
rect 996 132 998 134
rect 331 126 333 128
rect 336 126 338 128
rect 341 126 343 128
rect 346 126 348 128
rect 351 126 353 128
rect 356 126 358 128
rect 361 126 363 128
rect 366 126 368 128
rect 371 126 373 128
rect 376 126 378 128
rect 381 126 383 128
rect 386 126 388 128
rect 391 126 393 128
rect 396 126 398 128
rect 401 126 403 128
rect 406 126 408 128
rect 411 126 413 128
rect 416 126 418 128
rect 421 126 423 128
rect 426 126 428 128
rect 431 126 433 128
rect 436 126 438 128
rect 441 126 443 128
rect 446 126 448 128
rect 451 126 453 128
rect 456 126 458 128
rect 461 126 463 128
rect 466 126 468 128
rect 471 126 473 128
rect 476 126 478 128
rect 481 126 483 128
rect 486 126 488 128
rect 491 126 493 128
rect 496 126 498 128
rect 501 126 503 128
rect 506 126 508 128
rect 511 126 513 128
rect 516 126 518 128
rect 521 126 523 128
rect 526 126 528 128
rect 531 126 533 128
rect 536 126 538 128
rect 541 126 543 128
rect 546 126 548 128
rect 551 126 553 128
rect 556 126 558 128
rect 771 127 773 129
rect 776 127 778 129
rect 781 127 783 129
rect 786 127 788 129
rect 791 127 793 129
rect 796 127 798 129
rect 801 127 803 129
rect 806 127 808 129
rect 811 127 813 129
rect 816 127 818 129
rect 821 127 823 129
rect 826 127 828 129
rect 831 127 833 129
rect 836 127 838 129
rect 841 127 843 129
rect 846 127 848 129
rect 851 127 853 129
rect 856 127 858 129
rect 861 127 863 129
rect 866 127 868 129
rect 871 127 873 129
rect 876 127 878 129
rect 881 127 883 129
rect 886 127 888 129
rect 891 127 893 129
rect 896 127 898 129
rect 901 127 903 129
rect 906 127 908 129
rect 911 127 913 129
rect 916 127 918 129
rect 921 127 923 129
rect 926 127 928 129
rect 931 127 933 129
rect 936 127 938 129
rect 941 127 943 129
rect 946 127 948 129
rect 951 127 953 129
rect 956 127 958 129
rect 961 127 963 129
rect 966 127 968 129
rect 971 127 973 129
rect 976 127 978 129
rect 981 127 983 129
rect 986 127 988 129
rect 991 127 993 129
rect 996 127 998 129
rect 331 121 333 123
rect 336 121 338 123
rect 341 121 343 123
rect 346 121 348 123
rect 351 121 353 123
rect 356 121 358 123
rect 361 121 363 123
rect 366 121 368 123
rect 371 121 373 123
rect 376 121 378 123
rect 381 121 383 123
rect 386 121 388 123
rect 391 121 393 123
rect 396 121 398 123
rect 401 121 403 123
rect 406 121 408 123
rect 411 121 413 123
rect 416 121 418 123
rect 421 121 423 123
rect 426 121 428 123
rect 431 121 433 123
rect 436 121 438 123
rect 441 121 443 123
rect 446 121 448 123
rect 451 121 453 123
rect 456 121 458 123
rect 461 121 463 123
rect 466 121 468 123
rect 471 121 473 123
rect 476 121 478 123
rect 481 121 483 123
rect 486 121 488 123
rect 491 121 493 123
rect 496 121 498 123
rect 501 121 503 123
rect 506 121 508 123
rect 511 121 513 123
rect 516 121 518 123
rect 521 121 523 123
rect 526 121 528 123
rect 531 121 533 123
rect 536 121 538 123
rect 541 121 543 123
rect 546 121 548 123
rect 551 121 553 123
rect 556 121 558 123
rect 771 122 773 124
rect 776 122 778 124
rect 781 122 783 124
rect 786 122 788 124
rect 791 122 793 124
rect 796 122 798 124
rect 801 122 803 124
rect 806 122 808 124
rect 811 122 813 124
rect 816 122 818 124
rect 821 122 823 124
rect 826 122 828 124
rect 831 122 833 124
rect 836 122 838 124
rect 841 122 843 124
rect 846 122 848 124
rect 851 122 853 124
rect 856 122 858 124
rect 861 122 863 124
rect 866 122 868 124
rect 871 122 873 124
rect 876 122 878 124
rect 881 122 883 124
rect 886 122 888 124
rect 891 122 893 124
rect 896 122 898 124
rect 901 122 903 124
rect 906 122 908 124
rect 911 122 913 124
rect 916 122 918 124
rect 921 122 923 124
rect 926 122 928 124
rect 931 122 933 124
rect 936 122 938 124
rect 941 122 943 124
rect 946 122 948 124
rect 951 122 953 124
rect 956 122 958 124
rect 961 122 963 124
rect 966 122 968 124
rect 971 122 973 124
rect 976 122 978 124
rect 981 122 983 124
rect 986 122 988 124
rect 991 122 993 124
rect 996 122 998 124
rect 331 116 333 118
rect 336 116 338 118
rect 341 116 343 118
rect 346 116 348 118
rect 351 116 353 118
rect 356 116 358 118
rect 361 116 363 118
rect 366 116 368 118
rect 371 116 373 118
rect 376 116 378 118
rect 381 116 383 118
rect 386 116 388 118
rect 391 116 393 118
rect 396 116 398 118
rect 401 116 403 118
rect 406 116 408 118
rect 411 116 413 118
rect 416 116 418 118
rect 421 116 423 118
rect 426 116 428 118
rect 431 116 433 118
rect 436 116 438 118
rect 441 116 443 118
rect 446 116 448 118
rect 451 116 453 118
rect 456 116 458 118
rect 461 116 463 118
rect 466 116 468 118
rect 471 116 473 118
rect 476 116 478 118
rect 481 116 483 118
rect 486 116 488 118
rect 491 116 493 118
rect 496 116 498 118
rect 501 116 503 118
rect 506 116 508 118
rect 511 116 513 118
rect 516 116 518 118
rect 521 116 523 118
rect 526 116 528 118
rect 531 116 533 118
rect 536 116 538 118
rect 541 116 543 118
rect 546 116 548 118
rect 551 116 553 118
rect 556 116 558 118
rect 771 117 773 119
rect 776 117 778 119
rect 781 117 783 119
rect 786 117 788 119
rect 791 117 793 119
rect 796 117 798 119
rect 801 117 803 119
rect 806 117 808 119
rect 811 117 813 119
rect 816 117 818 119
rect 821 117 823 119
rect 826 117 828 119
rect 831 117 833 119
rect 836 117 838 119
rect 841 117 843 119
rect 846 117 848 119
rect 851 117 853 119
rect 856 117 858 119
rect 861 117 863 119
rect 866 117 868 119
rect 871 117 873 119
rect 876 117 878 119
rect 881 117 883 119
rect 886 117 888 119
rect 891 117 893 119
rect 896 117 898 119
rect 901 117 903 119
rect 906 117 908 119
rect 911 117 913 119
rect 916 117 918 119
rect 921 117 923 119
rect 926 117 928 119
rect 931 117 933 119
rect 936 117 938 119
rect 941 117 943 119
rect 946 117 948 119
rect 951 117 953 119
rect 956 117 958 119
rect 961 117 963 119
rect 966 117 968 119
rect 971 117 973 119
rect 976 117 978 119
rect 981 117 983 119
rect 986 117 988 119
rect 991 117 993 119
rect 996 117 998 119
rect 331 111 333 113
rect 336 111 338 113
rect 341 111 343 113
rect 346 111 348 113
rect 351 111 353 113
rect 356 111 358 113
rect 361 111 363 113
rect 366 111 368 113
rect 371 111 373 113
rect 376 111 378 113
rect 381 111 383 113
rect 386 111 388 113
rect 391 111 393 113
rect 396 111 398 113
rect 401 111 403 113
rect 406 111 408 113
rect 411 111 413 113
rect 416 111 418 113
rect 421 111 423 113
rect 426 111 428 113
rect 431 111 433 113
rect 436 111 438 113
rect 441 111 443 113
rect 446 111 448 113
rect 451 111 453 113
rect 456 111 458 113
rect 461 111 463 113
rect 466 111 468 113
rect 471 111 473 113
rect 476 111 478 113
rect 481 111 483 113
rect 486 111 488 113
rect 491 111 493 113
rect 496 111 498 113
rect 501 111 503 113
rect 506 111 508 113
rect 511 111 513 113
rect 516 111 518 113
rect 521 111 523 113
rect 526 111 528 113
rect 531 111 533 113
rect 536 111 538 113
rect 541 111 543 113
rect 546 111 548 113
rect 551 111 553 113
rect 556 111 558 113
rect 771 112 773 114
rect 776 112 778 114
rect 781 112 783 114
rect 786 112 788 114
rect 791 112 793 114
rect 796 112 798 114
rect 801 112 803 114
rect 806 112 808 114
rect 811 112 813 114
rect 816 112 818 114
rect 821 112 823 114
rect 826 112 828 114
rect 831 112 833 114
rect 836 112 838 114
rect 841 112 843 114
rect 846 112 848 114
rect 851 112 853 114
rect 856 112 858 114
rect 861 112 863 114
rect 866 112 868 114
rect 871 112 873 114
rect 876 112 878 114
rect 881 112 883 114
rect 886 112 888 114
rect 891 112 893 114
rect 896 112 898 114
rect 901 112 903 114
rect 906 112 908 114
rect 911 112 913 114
rect 916 112 918 114
rect 921 112 923 114
rect 926 112 928 114
rect 931 112 933 114
rect 936 112 938 114
rect 941 112 943 114
rect 946 112 948 114
rect 951 112 953 114
rect 956 112 958 114
rect 961 112 963 114
rect 966 112 968 114
rect 971 112 973 114
rect 976 112 978 114
rect 981 112 983 114
rect 986 112 988 114
rect 991 112 993 114
rect 996 112 998 114
rect 331 106 333 108
rect 336 106 338 108
rect 341 106 343 108
rect 346 106 348 108
rect 351 106 353 108
rect 356 106 358 108
rect 361 106 363 108
rect 366 106 368 108
rect 371 106 373 108
rect 376 106 378 108
rect 381 106 383 108
rect 386 106 388 108
rect 391 106 393 108
rect 396 106 398 108
rect 401 106 403 108
rect 406 106 408 108
rect 411 106 413 108
rect 416 106 418 108
rect 421 106 423 108
rect 426 106 428 108
rect 431 106 433 108
rect 436 106 438 108
rect 441 106 443 108
rect 446 106 448 108
rect 451 106 453 108
rect 456 106 458 108
rect 461 106 463 108
rect 466 106 468 108
rect 471 106 473 108
rect 476 106 478 108
rect 481 106 483 108
rect 486 106 488 108
rect 491 106 493 108
rect 496 106 498 108
rect 501 106 503 108
rect 506 106 508 108
rect 511 106 513 108
rect 516 106 518 108
rect 521 106 523 108
rect 526 106 528 108
rect 531 106 533 108
rect 536 106 538 108
rect 541 106 543 108
rect 546 106 548 108
rect 551 106 553 108
rect 556 106 558 108
rect 771 107 773 109
rect 776 107 778 109
rect 781 107 783 109
rect 786 107 788 109
rect 791 107 793 109
rect 796 107 798 109
rect 801 107 803 109
rect 806 107 808 109
rect 811 107 813 109
rect 816 107 818 109
rect 821 107 823 109
rect 826 107 828 109
rect 831 107 833 109
rect 836 107 838 109
rect 841 107 843 109
rect 846 107 848 109
rect 851 107 853 109
rect 856 107 858 109
rect 861 107 863 109
rect 866 107 868 109
rect 871 107 873 109
rect 876 107 878 109
rect 881 107 883 109
rect 886 107 888 109
rect 891 107 893 109
rect 896 107 898 109
rect 901 107 903 109
rect 906 107 908 109
rect 911 107 913 109
rect 916 107 918 109
rect 921 107 923 109
rect 926 107 928 109
rect 931 107 933 109
rect 936 107 938 109
rect 941 107 943 109
rect 946 107 948 109
rect 951 107 953 109
rect 956 107 958 109
rect 961 107 963 109
rect 966 107 968 109
rect 971 107 973 109
rect 976 107 978 109
rect 981 107 983 109
rect 986 107 988 109
rect 991 107 993 109
rect 996 107 998 109
rect 331 101 333 103
rect 336 101 338 103
rect 341 101 343 103
rect 346 101 348 103
rect 351 101 353 103
rect 356 101 358 103
rect 361 101 363 103
rect 366 101 368 103
rect 371 101 373 103
rect 376 101 378 103
rect 381 101 383 103
rect 386 101 388 103
rect 391 101 393 103
rect 396 101 398 103
rect 401 101 403 103
rect 406 101 408 103
rect 411 101 413 103
rect 416 101 418 103
rect 421 101 423 103
rect 426 101 428 103
rect 431 101 433 103
rect 436 101 438 103
rect 441 101 443 103
rect 446 101 448 103
rect 451 101 453 103
rect 456 101 458 103
rect 461 101 463 103
rect 466 101 468 103
rect 471 101 473 103
rect 476 101 478 103
rect 481 101 483 103
rect 486 101 488 103
rect 491 101 493 103
rect 496 101 498 103
rect 501 101 503 103
rect 506 101 508 103
rect 511 101 513 103
rect 516 101 518 103
rect 521 101 523 103
rect 526 101 528 103
rect 531 101 533 103
rect 536 101 538 103
rect 541 101 543 103
rect 546 101 548 103
rect 551 101 553 103
rect 556 101 558 103
rect 771 102 773 104
rect 776 102 778 104
rect 781 102 783 104
rect 786 102 788 104
rect 791 102 793 104
rect 796 102 798 104
rect 801 102 803 104
rect 806 102 808 104
rect 811 102 813 104
rect 816 102 818 104
rect 821 102 823 104
rect 826 102 828 104
rect 831 102 833 104
rect 836 102 838 104
rect 841 102 843 104
rect 846 102 848 104
rect 851 102 853 104
rect 856 102 858 104
rect 861 102 863 104
rect 866 102 868 104
rect 871 102 873 104
rect 876 102 878 104
rect 881 102 883 104
rect 886 102 888 104
rect 891 102 893 104
rect 896 102 898 104
rect 901 102 903 104
rect 906 102 908 104
rect 911 102 913 104
rect 916 102 918 104
rect 921 102 923 104
rect 926 102 928 104
rect 931 102 933 104
rect 936 102 938 104
rect 941 102 943 104
rect 946 102 948 104
rect 951 102 953 104
rect 956 102 958 104
rect 961 102 963 104
rect 966 102 968 104
rect 971 102 973 104
rect 976 102 978 104
rect 981 102 983 104
rect 986 102 988 104
rect 991 102 993 104
rect 996 102 998 104
rect 331 96 333 98
rect 336 96 338 98
rect 341 96 343 98
rect 346 96 348 98
rect 351 96 353 98
rect 356 96 358 98
rect 361 96 363 98
rect 366 96 368 98
rect 371 96 373 98
rect 376 96 378 98
rect 381 96 383 98
rect 386 96 388 98
rect 391 96 393 98
rect 396 96 398 98
rect 401 96 403 98
rect 406 96 408 98
rect 411 96 413 98
rect 416 96 418 98
rect 421 96 423 98
rect 426 96 428 98
rect 431 96 433 98
rect 436 96 438 98
rect 441 96 443 98
rect 446 96 448 98
rect 451 96 453 98
rect 456 96 458 98
rect 461 96 463 98
rect 466 96 468 98
rect 471 96 473 98
rect 476 96 478 98
rect 481 96 483 98
rect 486 96 488 98
rect 491 96 493 98
rect 496 96 498 98
rect 501 96 503 98
rect 506 96 508 98
rect 511 96 513 98
rect 516 96 518 98
rect 521 96 523 98
rect 526 96 528 98
rect 531 96 533 98
rect 536 96 538 98
rect 541 96 543 98
rect 546 96 548 98
rect 551 96 553 98
rect 556 96 558 98
rect 771 97 773 99
rect 776 97 778 99
rect 781 97 783 99
rect 786 97 788 99
rect 791 97 793 99
rect 796 97 798 99
rect 801 97 803 99
rect 806 97 808 99
rect 811 97 813 99
rect 816 97 818 99
rect 821 97 823 99
rect 826 97 828 99
rect 831 97 833 99
rect 836 97 838 99
rect 841 97 843 99
rect 846 97 848 99
rect 851 97 853 99
rect 856 97 858 99
rect 861 97 863 99
rect 866 97 868 99
rect 871 97 873 99
rect 876 97 878 99
rect 881 97 883 99
rect 886 97 888 99
rect 891 97 893 99
rect 896 97 898 99
rect 901 97 903 99
rect 906 97 908 99
rect 911 97 913 99
rect 916 97 918 99
rect 921 97 923 99
rect 926 97 928 99
rect 931 97 933 99
rect 936 97 938 99
rect 941 97 943 99
rect 946 97 948 99
rect 951 97 953 99
rect 956 97 958 99
rect 961 97 963 99
rect 966 97 968 99
rect 971 97 973 99
rect 976 97 978 99
rect 981 97 983 99
rect 986 97 988 99
rect 991 97 993 99
rect 996 97 998 99
rect 331 91 333 93
rect 336 91 338 93
rect 341 91 343 93
rect 346 91 348 93
rect 351 91 353 93
rect 356 91 358 93
rect 361 91 363 93
rect 366 91 368 93
rect 371 91 373 93
rect 376 91 378 93
rect 381 91 383 93
rect 386 91 388 93
rect 391 91 393 93
rect 396 91 398 93
rect 401 91 403 93
rect 406 91 408 93
rect 411 91 413 93
rect 416 91 418 93
rect 421 91 423 93
rect 426 91 428 93
rect 431 91 433 93
rect 436 91 438 93
rect 441 91 443 93
rect 446 91 448 93
rect 451 91 453 93
rect 456 91 458 93
rect 461 91 463 93
rect 466 91 468 93
rect 471 91 473 93
rect 476 91 478 93
rect 481 91 483 93
rect 486 91 488 93
rect 491 91 493 93
rect 496 91 498 93
rect 501 91 503 93
rect 506 91 508 93
rect 511 91 513 93
rect 516 91 518 93
rect 521 91 523 93
rect 526 91 528 93
rect 531 91 533 93
rect 536 91 538 93
rect 541 91 543 93
rect 546 91 548 93
rect 551 91 553 93
rect 556 91 558 93
rect 771 92 773 94
rect 776 92 778 94
rect 781 92 783 94
rect 786 92 788 94
rect 791 92 793 94
rect 796 92 798 94
rect 801 92 803 94
rect 806 92 808 94
rect 811 92 813 94
rect 816 92 818 94
rect 821 92 823 94
rect 826 92 828 94
rect 831 92 833 94
rect 836 92 838 94
rect 841 92 843 94
rect 846 92 848 94
rect 851 92 853 94
rect 856 92 858 94
rect 861 92 863 94
rect 866 92 868 94
rect 871 92 873 94
rect 876 92 878 94
rect 881 92 883 94
rect 886 92 888 94
rect 891 92 893 94
rect 896 92 898 94
rect 901 92 903 94
rect 906 92 908 94
rect 911 92 913 94
rect 916 92 918 94
rect 921 92 923 94
rect 926 92 928 94
rect 931 92 933 94
rect 936 92 938 94
rect 941 92 943 94
rect 946 92 948 94
rect 951 92 953 94
rect 956 92 958 94
rect 961 92 963 94
rect 966 92 968 94
rect 971 92 973 94
rect 976 92 978 94
rect 981 92 983 94
rect 986 92 988 94
rect 991 92 993 94
rect 996 92 998 94
rect 331 86 333 88
rect 336 86 338 88
rect 341 86 343 88
rect 346 86 348 88
rect 351 86 353 88
rect 356 86 358 88
rect 361 86 363 88
rect 366 86 368 88
rect 371 86 373 88
rect 376 86 378 88
rect 381 86 383 88
rect 386 86 388 88
rect 391 86 393 88
rect 396 86 398 88
rect 401 86 403 88
rect 406 86 408 88
rect 411 86 413 88
rect 416 86 418 88
rect 421 86 423 88
rect 426 86 428 88
rect 431 86 433 88
rect 436 86 438 88
rect 441 86 443 88
rect 446 86 448 88
rect 451 86 453 88
rect 456 86 458 88
rect 461 86 463 88
rect 466 86 468 88
rect 471 86 473 88
rect 476 86 478 88
rect 481 86 483 88
rect 486 86 488 88
rect 491 86 493 88
rect 496 86 498 88
rect 501 86 503 88
rect 506 86 508 88
rect 511 86 513 88
rect 516 86 518 88
rect 521 86 523 88
rect 526 86 528 88
rect 531 86 533 88
rect 536 86 538 88
rect 541 86 543 88
rect 546 86 548 88
rect 551 86 553 88
rect 556 86 558 88
rect 771 87 773 89
rect 776 87 778 89
rect 781 87 783 89
rect 786 87 788 89
rect 791 87 793 89
rect 796 87 798 89
rect 801 87 803 89
rect 806 87 808 89
rect 811 87 813 89
rect 816 87 818 89
rect 821 87 823 89
rect 826 87 828 89
rect 831 87 833 89
rect 836 87 838 89
rect 841 87 843 89
rect 846 87 848 89
rect 851 87 853 89
rect 856 87 858 89
rect 861 87 863 89
rect 866 87 868 89
rect 871 87 873 89
rect 876 87 878 89
rect 881 87 883 89
rect 886 87 888 89
rect 891 87 893 89
rect 896 87 898 89
rect 901 87 903 89
rect 906 87 908 89
rect 911 87 913 89
rect 916 87 918 89
rect 921 87 923 89
rect 926 87 928 89
rect 931 87 933 89
rect 936 87 938 89
rect 941 87 943 89
rect 946 87 948 89
rect 951 87 953 89
rect 956 87 958 89
rect 961 87 963 89
rect 966 87 968 89
rect 971 87 973 89
rect 976 87 978 89
rect 981 87 983 89
rect 986 87 988 89
rect 991 87 993 89
rect 996 87 998 89
rect 331 81 333 83
rect 336 81 338 83
rect 341 81 343 83
rect 346 81 348 83
rect 351 81 353 83
rect 356 81 358 83
rect 361 81 363 83
rect 366 81 368 83
rect 371 81 373 83
rect 376 81 378 83
rect 381 81 383 83
rect 386 81 388 83
rect 391 81 393 83
rect 396 81 398 83
rect 401 81 403 83
rect 406 81 408 83
rect 411 81 413 83
rect 416 81 418 83
rect 421 81 423 83
rect 426 81 428 83
rect 431 81 433 83
rect 436 81 438 83
rect 441 81 443 83
rect 446 81 448 83
rect 451 81 453 83
rect 456 81 458 83
rect 461 81 463 83
rect 466 81 468 83
rect 471 81 473 83
rect 476 81 478 83
rect 481 81 483 83
rect 486 81 488 83
rect 491 81 493 83
rect 496 81 498 83
rect 501 81 503 83
rect 506 81 508 83
rect 511 81 513 83
rect 516 81 518 83
rect 521 81 523 83
rect 526 81 528 83
rect 531 81 533 83
rect 536 81 538 83
rect 541 81 543 83
rect 546 81 548 83
rect 551 81 553 83
rect 556 81 558 83
rect 771 82 773 84
rect 776 82 778 84
rect 781 82 783 84
rect 786 82 788 84
rect 791 82 793 84
rect 796 82 798 84
rect 801 82 803 84
rect 806 82 808 84
rect 811 82 813 84
rect 816 82 818 84
rect 821 82 823 84
rect 826 82 828 84
rect 831 82 833 84
rect 836 82 838 84
rect 841 82 843 84
rect 846 82 848 84
rect 851 82 853 84
rect 856 82 858 84
rect 861 82 863 84
rect 866 82 868 84
rect 871 82 873 84
rect 876 82 878 84
rect 881 82 883 84
rect 886 82 888 84
rect 891 82 893 84
rect 896 82 898 84
rect 901 82 903 84
rect 906 82 908 84
rect 911 82 913 84
rect 916 82 918 84
rect 921 82 923 84
rect 926 82 928 84
rect 931 82 933 84
rect 936 82 938 84
rect 941 82 943 84
rect 946 82 948 84
rect 951 82 953 84
rect 956 82 958 84
rect 961 82 963 84
rect 966 82 968 84
rect 971 82 973 84
rect 976 82 978 84
rect 981 82 983 84
rect 986 82 988 84
rect 991 82 993 84
rect 996 82 998 84
rect 331 76 333 78
rect 336 76 338 78
rect 341 76 343 78
rect 346 76 348 78
rect 351 76 353 78
rect 356 76 358 78
rect 361 76 363 78
rect 366 76 368 78
rect 371 76 373 78
rect 376 76 378 78
rect 381 76 383 78
rect 386 76 388 78
rect 391 76 393 78
rect 396 76 398 78
rect 401 76 403 78
rect 406 76 408 78
rect 411 76 413 78
rect 416 76 418 78
rect 421 76 423 78
rect 426 76 428 78
rect 431 76 433 78
rect 436 76 438 78
rect 441 76 443 78
rect 446 76 448 78
rect 451 76 453 78
rect 456 76 458 78
rect 461 76 463 78
rect 466 76 468 78
rect 471 76 473 78
rect 476 76 478 78
rect 481 76 483 78
rect 486 76 488 78
rect 491 76 493 78
rect 496 76 498 78
rect 501 76 503 78
rect 506 76 508 78
rect 511 76 513 78
rect 516 76 518 78
rect 521 76 523 78
rect 526 76 528 78
rect 531 76 533 78
rect 536 76 538 78
rect 541 76 543 78
rect 546 76 548 78
rect 551 76 553 78
rect 556 76 558 78
rect 771 77 773 79
rect 776 77 778 79
rect 781 77 783 79
rect 786 77 788 79
rect 791 77 793 79
rect 796 77 798 79
rect 801 77 803 79
rect 806 77 808 79
rect 811 77 813 79
rect 816 77 818 79
rect 821 77 823 79
rect 826 77 828 79
rect 831 77 833 79
rect 836 77 838 79
rect 841 77 843 79
rect 846 77 848 79
rect 851 77 853 79
rect 856 77 858 79
rect 861 77 863 79
rect 866 77 868 79
rect 871 77 873 79
rect 876 77 878 79
rect 881 77 883 79
rect 886 77 888 79
rect 891 77 893 79
rect 896 77 898 79
rect 901 77 903 79
rect 906 77 908 79
rect 911 77 913 79
rect 916 77 918 79
rect 921 77 923 79
rect 926 77 928 79
rect 931 77 933 79
rect 936 77 938 79
rect 941 77 943 79
rect 946 77 948 79
rect 951 77 953 79
rect 956 77 958 79
rect 961 77 963 79
rect 966 77 968 79
rect 971 77 973 79
rect 976 77 978 79
rect 981 77 983 79
rect 986 77 988 79
rect 991 77 993 79
rect 996 77 998 79
rect 331 71 333 73
rect 336 71 338 73
rect 341 71 343 73
rect 346 71 348 73
rect 351 71 353 73
rect 356 71 358 73
rect 361 71 363 73
rect 366 71 368 73
rect 371 71 373 73
rect 376 71 378 73
rect 381 71 383 73
rect 386 71 388 73
rect 391 71 393 73
rect 396 71 398 73
rect 401 71 403 73
rect 406 71 408 73
rect 411 71 413 73
rect 416 71 418 73
rect 421 71 423 73
rect 426 71 428 73
rect 431 71 433 73
rect 436 71 438 73
rect 441 71 443 73
rect 446 71 448 73
rect 451 71 453 73
rect 456 71 458 73
rect 461 71 463 73
rect 466 71 468 73
rect 471 71 473 73
rect 476 71 478 73
rect 481 71 483 73
rect 486 71 488 73
rect 491 71 493 73
rect 496 71 498 73
rect 501 71 503 73
rect 506 71 508 73
rect 511 71 513 73
rect 516 71 518 73
rect 521 71 523 73
rect 526 71 528 73
rect 531 71 533 73
rect 536 71 538 73
rect 541 71 543 73
rect 546 71 548 73
rect 551 71 553 73
rect 556 71 558 73
rect 771 72 773 74
rect 776 72 778 74
rect 781 72 783 74
rect 786 72 788 74
rect 791 72 793 74
rect 796 72 798 74
rect 801 72 803 74
rect 806 72 808 74
rect 811 72 813 74
rect 816 72 818 74
rect 821 72 823 74
rect 826 72 828 74
rect 831 72 833 74
rect 836 72 838 74
rect 841 72 843 74
rect 846 72 848 74
rect 851 72 853 74
rect 856 72 858 74
rect 861 72 863 74
rect 866 72 868 74
rect 871 72 873 74
rect 876 72 878 74
rect 881 72 883 74
rect 886 72 888 74
rect 891 72 893 74
rect 896 72 898 74
rect 901 72 903 74
rect 906 72 908 74
rect 911 72 913 74
rect 916 72 918 74
rect 921 72 923 74
rect 926 72 928 74
rect 931 72 933 74
rect 936 72 938 74
rect 941 72 943 74
rect 946 72 948 74
rect 951 72 953 74
rect 956 72 958 74
rect 961 72 963 74
rect 966 72 968 74
rect 971 72 973 74
rect 976 72 978 74
rect 981 72 983 74
rect 986 72 988 74
rect 991 72 993 74
rect 996 72 998 74
rect 331 66 333 68
rect 336 66 338 68
rect 341 66 343 68
rect 346 66 348 68
rect 351 66 353 68
rect 356 66 358 68
rect 361 66 363 68
rect 366 66 368 68
rect 371 66 373 68
rect 376 66 378 68
rect 381 66 383 68
rect 386 66 388 68
rect 391 66 393 68
rect 396 66 398 68
rect 401 66 403 68
rect 406 66 408 68
rect 411 66 413 68
rect 416 66 418 68
rect 421 66 423 68
rect 426 66 428 68
rect 431 66 433 68
rect 436 66 438 68
rect 441 66 443 68
rect 446 66 448 68
rect 451 66 453 68
rect 456 66 458 68
rect 461 66 463 68
rect 466 66 468 68
rect 471 66 473 68
rect 476 66 478 68
rect 481 66 483 68
rect 486 66 488 68
rect 491 66 493 68
rect 496 66 498 68
rect 501 66 503 68
rect 506 66 508 68
rect 511 66 513 68
rect 516 66 518 68
rect 521 66 523 68
rect 526 66 528 68
rect 531 66 533 68
rect 536 66 538 68
rect 541 66 543 68
rect 546 66 548 68
rect 551 66 553 68
rect 556 66 558 68
rect 771 67 773 69
rect 776 67 778 69
rect 781 67 783 69
rect 786 67 788 69
rect 791 67 793 69
rect 796 67 798 69
rect 801 67 803 69
rect 806 67 808 69
rect 811 67 813 69
rect 816 67 818 69
rect 821 67 823 69
rect 826 67 828 69
rect 831 67 833 69
rect 836 67 838 69
rect 841 67 843 69
rect 846 67 848 69
rect 851 67 853 69
rect 856 67 858 69
rect 861 67 863 69
rect 866 67 868 69
rect 871 67 873 69
rect 876 67 878 69
rect 881 67 883 69
rect 886 67 888 69
rect 891 67 893 69
rect 896 67 898 69
rect 901 67 903 69
rect 906 67 908 69
rect 911 67 913 69
rect 916 67 918 69
rect 921 67 923 69
rect 926 67 928 69
rect 931 67 933 69
rect 936 67 938 69
rect 941 67 943 69
rect 946 67 948 69
rect 951 67 953 69
rect 956 67 958 69
rect 961 67 963 69
rect 966 67 968 69
rect 971 67 973 69
rect 976 67 978 69
rect 981 67 983 69
rect 986 67 988 69
rect 991 67 993 69
rect 996 67 998 69
rect 331 61 333 63
rect 336 61 338 63
rect 341 61 343 63
rect 346 61 348 63
rect 351 61 353 63
rect 356 61 358 63
rect 361 61 363 63
rect 366 61 368 63
rect 371 61 373 63
rect 376 61 378 63
rect 381 61 383 63
rect 386 61 388 63
rect 391 61 393 63
rect 396 61 398 63
rect 401 61 403 63
rect 406 61 408 63
rect 411 61 413 63
rect 416 61 418 63
rect 421 61 423 63
rect 426 61 428 63
rect 431 61 433 63
rect 436 61 438 63
rect 441 61 443 63
rect 446 61 448 63
rect 451 61 453 63
rect 456 61 458 63
rect 461 61 463 63
rect 466 61 468 63
rect 471 61 473 63
rect 476 61 478 63
rect 481 61 483 63
rect 486 61 488 63
rect 491 61 493 63
rect 496 61 498 63
rect 501 61 503 63
rect 506 61 508 63
rect 511 61 513 63
rect 516 61 518 63
rect 521 61 523 63
rect 526 61 528 63
rect 531 61 533 63
rect 536 61 538 63
rect 541 61 543 63
rect 546 61 548 63
rect 551 61 553 63
rect 556 61 558 63
rect 771 62 773 64
rect 776 62 778 64
rect 781 62 783 64
rect 786 62 788 64
rect 791 62 793 64
rect 796 62 798 64
rect 801 62 803 64
rect 806 62 808 64
rect 811 62 813 64
rect 816 62 818 64
rect 821 62 823 64
rect 826 62 828 64
rect 831 62 833 64
rect 836 62 838 64
rect 841 62 843 64
rect 846 62 848 64
rect 851 62 853 64
rect 856 62 858 64
rect 861 62 863 64
rect 866 62 868 64
rect 871 62 873 64
rect 876 62 878 64
rect 881 62 883 64
rect 886 62 888 64
rect 891 62 893 64
rect 896 62 898 64
rect 901 62 903 64
rect 906 62 908 64
rect 911 62 913 64
rect 916 62 918 64
rect 921 62 923 64
rect 926 62 928 64
rect 931 62 933 64
rect 936 62 938 64
rect 941 62 943 64
rect 946 62 948 64
rect 951 62 953 64
rect 956 62 958 64
rect 961 62 963 64
rect 966 62 968 64
rect 971 62 973 64
rect 976 62 978 64
rect 981 62 983 64
rect 986 62 988 64
rect 991 62 993 64
rect 996 62 998 64
rect 331 56 333 58
rect 336 56 338 58
rect 341 56 343 58
rect 346 56 348 58
rect 351 56 353 58
rect 356 56 358 58
rect 361 56 363 58
rect 366 56 368 58
rect 371 56 373 58
rect 376 56 378 58
rect 381 56 383 58
rect 386 56 388 58
rect 391 56 393 58
rect 396 56 398 58
rect 401 56 403 58
rect 406 56 408 58
rect 411 56 413 58
rect 416 56 418 58
rect 421 56 423 58
rect 426 56 428 58
rect 431 56 433 58
rect 436 56 438 58
rect 441 56 443 58
rect 446 56 448 58
rect 451 56 453 58
rect 456 56 458 58
rect 461 56 463 58
rect 466 56 468 58
rect 471 56 473 58
rect 476 56 478 58
rect 481 56 483 58
rect 486 56 488 58
rect 491 56 493 58
rect 496 56 498 58
rect 501 56 503 58
rect 506 56 508 58
rect 511 56 513 58
rect 516 56 518 58
rect 521 56 523 58
rect 526 56 528 58
rect 531 56 533 58
rect 536 56 538 58
rect 541 56 543 58
rect 546 56 548 58
rect 551 56 553 58
rect 556 56 558 58
rect 771 57 773 59
rect 776 57 778 59
rect 781 57 783 59
rect 786 57 788 59
rect 791 57 793 59
rect 796 57 798 59
rect 801 57 803 59
rect 806 57 808 59
rect 811 57 813 59
rect 816 57 818 59
rect 821 57 823 59
rect 826 57 828 59
rect 831 57 833 59
rect 836 57 838 59
rect 841 57 843 59
rect 846 57 848 59
rect 851 57 853 59
rect 856 57 858 59
rect 861 57 863 59
rect 866 57 868 59
rect 871 57 873 59
rect 876 57 878 59
rect 881 57 883 59
rect 886 57 888 59
rect 891 57 893 59
rect 896 57 898 59
rect 901 57 903 59
rect 906 57 908 59
rect 911 57 913 59
rect 916 57 918 59
rect 921 57 923 59
rect 926 57 928 59
rect 931 57 933 59
rect 936 57 938 59
rect 941 57 943 59
rect 946 57 948 59
rect 951 57 953 59
rect 956 57 958 59
rect 961 57 963 59
rect 966 57 968 59
rect 971 57 973 59
rect 976 57 978 59
rect 981 57 983 59
rect 986 57 988 59
rect 991 57 993 59
rect 996 57 998 59
rect 331 51 333 53
rect 336 51 338 53
rect 341 51 343 53
rect 346 51 348 53
rect 351 51 353 53
rect 356 51 358 53
rect 361 51 363 53
rect 366 51 368 53
rect 371 51 373 53
rect 376 51 378 53
rect 381 51 383 53
rect 386 51 388 53
rect 391 51 393 53
rect 396 51 398 53
rect 401 51 403 53
rect 406 51 408 53
rect 411 51 413 53
rect 416 51 418 53
rect 421 51 423 53
rect 426 51 428 53
rect 431 51 433 53
rect 436 51 438 53
rect 441 51 443 53
rect 446 51 448 53
rect 451 51 453 53
rect 456 51 458 53
rect 461 51 463 53
rect 466 51 468 53
rect 471 51 473 53
rect 476 51 478 53
rect 481 51 483 53
rect 486 51 488 53
rect 491 51 493 53
rect 496 51 498 53
rect 501 51 503 53
rect 506 51 508 53
rect 511 51 513 53
rect 516 51 518 53
rect 521 51 523 53
rect 526 51 528 53
rect 531 51 533 53
rect 536 51 538 53
rect 541 51 543 53
rect 546 51 548 53
rect 551 51 553 53
rect 556 51 558 53
rect 771 52 773 54
rect 776 52 778 54
rect 781 52 783 54
rect 786 52 788 54
rect 791 52 793 54
rect 796 52 798 54
rect 801 52 803 54
rect 806 52 808 54
rect 811 52 813 54
rect 816 52 818 54
rect 821 52 823 54
rect 826 52 828 54
rect 831 52 833 54
rect 836 52 838 54
rect 841 52 843 54
rect 846 52 848 54
rect 851 52 853 54
rect 856 52 858 54
rect 861 52 863 54
rect 866 52 868 54
rect 871 52 873 54
rect 876 52 878 54
rect 881 52 883 54
rect 886 52 888 54
rect 891 52 893 54
rect 896 52 898 54
rect 901 52 903 54
rect 906 52 908 54
rect 911 52 913 54
rect 916 52 918 54
rect 921 52 923 54
rect 926 52 928 54
rect 931 52 933 54
rect 936 52 938 54
rect 941 52 943 54
rect 946 52 948 54
rect 951 52 953 54
rect 956 52 958 54
rect 961 52 963 54
rect 966 52 968 54
rect 971 52 973 54
rect 976 52 978 54
rect 981 52 983 54
rect 986 52 988 54
rect 991 52 993 54
rect 996 52 998 54
rect 331 46 333 48
rect 336 46 338 48
rect 341 46 343 48
rect 346 46 348 48
rect 351 46 353 48
rect 356 46 358 48
rect 361 46 363 48
rect 366 46 368 48
rect 371 46 373 48
rect 376 46 378 48
rect 381 46 383 48
rect 386 46 388 48
rect 391 46 393 48
rect 396 46 398 48
rect 401 46 403 48
rect 406 46 408 48
rect 411 46 413 48
rect 416 46 418 48
rect 421 46 423 48
rect 426 46 428 48
rect 431 46 433 48
rect 436 46 438 48
rect 441 46 443 48
rect 446 46 448 48
rect 451 46 453 48
rect 456 46 458 48
rect 461 46 463 48
rect 466 46 468 48
rect 471 46 473 48
rect 476 46 478 48
rect 481 46 483 48
rect 486 46 488 48
rect 491 46 493 48
rect 496 46 498 48
rect 501 46 503 48
rect 506 46 508 48
rect 511 46 513 48
rect 516 46 518 48
rect 521 46 523 48
rect 526 46 528 48
rect 531 46 533 48
rect 536 46 538 48
rect 541 46 543 48
rect 546 46 548 48
rect 551 46 553 48
rect 556 46 558 48
rect 771 47 773 49
rect 776 47 778 49
rect 781 47 783 49
rect 786 47 788 49
rect 791 47 793 49
rect 796 47 798 49
rect 801 47 803 49
rect 806 47 808 49
rect 811 47 813 49
rect 816 47 818 49
rect 821 47 823 49
rect 826 47 828 49
rect 831 47 833 49
rect 836 47 838 49
rect 841 47 843 49
rect 846 47 848 49
rect 851 47 853 49
rect 856 47 858 49
rect 861 47 863 49
rect 866 47 868 49
rect 871 47 873 49
rect 876 47 878 49
rect 881 47 883 49
rect 886 47 888 49
rect 891 47 893 49
rect 896 47 898 49
rect 901 47 903 49
rect 906 47 908 49
rect 911 47 913 49
rect 916 47 918 49
rect 921 47 923 49
rect 926 47 928 49
rect 931 47 933 49
rect 936 47 938 49
rect 941 47 943 49
rect 946 47 948 49
rect 951 47 953 49
rect 956 47 958 49
rect 961 47 963 49
rect 966 47 968 49
rect 971 47 973 49
rect 976 47 978 49
rect 981 47 983 49
rect 986 47 988 49
rect 991 47 993 49
rect 996 47 998 49
rect 331 41 333 43
rect 336 41 338 43
rect 341 41 343 43
rect 346 41 348 43
rect 351 41 353 43
rect 356 41 358 43
rect 361 41 363 43
rect 366 41 368 43
rect 371 41 373 43
rect 376 41 378 43
rect 381 41 383 43
rect 386 41 388 43
rect 391 41 393 43
rect 396 41 398 43
rect 401 41 403 43
rect 406 41 408 43
rect 411 41 413 43
rect 416 41 418 43
rect 421 41 423 43
rect 426 41 428 43
rect 431 41 433 43
rect 436 41 438 43
rect 441 41 443 43
rect 446 41 448 43
rect 451 41 453 43
rect 456 41 458 43
rect 461 41 463 43
rect 466 41 468 43
rect 471 41 473 43
rect 476 41 478 43
rect 481 41 483 43
rect 486 41 488 43
rect 491 41 493 43
rect 496 41 498 43
rect 501 41 503 43
rect 506 41 508 43
rect 511 41 513 43
rect 516 41 518 43
rect 521 41 523 43
rect 526 41 528 43
rect 531 41 533 43
rect 536 41 538 43
rect 541 41 543 43
rect 546 41 548 43
rect 551 41 553 43
rect 556 41 558 43
rect 771 42 773 44
rect 776 42 778 44
rect 781 42 783 44
rect 786 42 788 44
rect 791 42 793 44
rect 796 42 798 44
rect 801 42 803 44
rect 806 42 808 44
rect 811 42 813 44
rect 816 42 818 44
rect 821 42 823 44
rect 826 42 828 44
rect 831 42 833 44
rect 836 42 838 44
rect 841 42 843 44
rect 846 42 848 44
rect 851 42 853 44
rect 856 42 858 44
rect 861 42 863 44
rect 866 42 868 44
rect 871 42 873 44
rect 876 42 878 44
rect 881 42 883 44
rect 886 42 888 44
rect 891 42 893 44
rect 896 42 898 44
rect 901 42 903 44
rect 906 42 908 44
rect 911 42 913 44
rect 916 42 918 44
rect 921 42 923 44
rect 926 42 928 44
rect 931 42 933 44
rect 936 42 938 44
rect 941 42 943 44
rect 946 42 948 44
rect 951 42 953 44
rect 956 42 958 44
rect 961 42 963 44
rect 966 42 968 44
rect 971 42 973 44
rect 976 42 978 44
rect 981 42 983 44
rect 986 42 988 44
rect 991 42 993 44
rect 996 42 998 44
rect 331 36 333 38
rect 336 36 338 38
rect 341 36 343 38
rect 346 36 348 38
rect 351 36 353 38
rect 356 36 358 38
rect 361 36 363 38
rect 366 36 368 38
rect 371 36 373 38
rect 376 36 378 38
rect 381 36 383 38
rect 386 36 388 38
rect 391 36 393 38
rect 396 36 398 38
rect 401 36 403 38
rect 406 36 408 38
rect 411 36 413 38
rect 416 36 418 38
rect 421 36 423 38
rect 426 36 428 38
rect 431 36 433 38
rect 436 36 438 38
rect 441 36 443 38
rect 446 36 448 38
rect 451 36 453 38
rect 456 36 458 38
rect 461 36 463 38
rect 466 36 468 38
rect 471 36 473 38
rect 476 36 478 38
rect 481 36 483 38
rect 486 36 488 38
rect 491 36 493 38
rect 496 36 498 38
rect 501 36 503 38
rect 506 36 508 38
rect 511 36 513 38
rect 516 36 518 38
rect 521 36 523 38
rect 526 36 528 38
rect 531 36 533 38
rect 536 36 538 38
rect 541 36 543 38
rect 546 36 548 38
rect 551 36 553 38
rect 556 36 558 38
rect 771 37 773 39
rect 776 37 778 39
rect 781 37 783 39
rect 786 37 788 39
rect 791 37 793 39
rect 796 37 798 39
rect 801 37 803 39
rect 806 37 808 39
rect 811 37 813 39
rect 816 37 818 39
rect 821 37 823 39
rect 826 37 828 39
rect 831 37 833 39
rect 836 37 838 39
rect 841 37 843 39
rect 846 37 848 39
rect 851 37 853 39
rect 856 37 858 39
rect 861 37 863 39
rect 866 37 868 39
rect 871 37 873 39
rect 876 37 878 39
rect 881 37 883 39
rect 886 37 888 39
rect 891 37 893 39
rect 896 37 898 39
rect 901 37 903 39
rect 906 37 908 39
rect 911 37 913 39
rect 916 37 918 39
rect 921 37 923 39
rect 926 37 928 39
rect 931 37 933 39
rect 936 37 938 39
rect 941 37 943 39
rect 946 37 948 39
rect 951 37 953 39
rect 956 37 958 39
rect 961 37 963 39
rect 966 37 968 39
rect 971 37 973 39
rect 976 37 978 39
rect 981 37 983 39
rect 986 37 988 39
rect 991 37 993 39
rect 996 37 998 39
rect 331 31 333 33
rect 336 31 338 33
rect 341 31 343 33
rect 346 31 348 33
rect 351 31 353 33
rect 356 31 358 33
rect 361 31 363 33
rect 366 31 368 33
rect 371 31 373 33
rect 376 31 378 33
rect 381 31 383 33
rect 386 31 388 33
rect 391 31 393 33
rect 396 31 398 33
rect 401 31 403 33
rect 406 31 408 33
rect 411 31 413 33
rect 416 31 418 33
rect 421 31 423 33
rect 426 31 428 33
rect 431 31 433 33
rect 436 31 438 33
rect 441 31 443 33
rect 446 31 448 33
rect 451 31 453 33
rect 456 31 458 33
rect 461 31 463 33
rect 466 31 468 33
rect 471 31 473 33
rect 476 31 478 33
rect 481 31 483 33
rect 486 31 488 33
rect 491 31 493 33
rect 496 31 498 33
rect 501 31 503 33
rect 506 31 508 33
rect 511 31 513 33
rect 516 31 518 33
rect 521 31 523 33
rect 526 31 528 33
rect 531 31 533 33
rect 536 31 538 33
rect 541 31 543 33
rect 546 31 548 33
rect 551 31 553 33
rect 556 31 558 33
rect 771 32 773 34
rect 776 32 778 34
rect 781 32 783 34
rect 786 32 788 34
rect 791 32 793 34
rect 796 32 798 34
rect 801 32 803 34
rect 806 32 808 34
rect 811 32 813 34
rect 816 32 818 34
rect 821 32 823 34
rect 826 32 828 34
rect 831 32 833 34
rect 836 32 838 34
rect 841 32 843 34
rect 846 32 848 34
rect 851 32 853 34
rect 856 32 858 34
rect 861 32 863 34
rect 866 32 868 34
rect 871 32 873 34
rect 876 32 878 34
rect 881 32 883 34
rect 886 32 888 34
rect 891 32 893 34
rect 896 32 898 34
rect 901 32 903 34
rect 906 32 908 34
rect 911 32 913 34
rect 916 32 918 34
rect 921 32 923 34
rect 926 32 928 34
rect 931 32 933 34
rect 936 32 938 34
rect 941 32 943 34
rect 946 32 948 34
rect 951 32 953 34
rect 956 32 958 34
rect 961 32 963 34
rect 966 32 968 34
rect 971 32 973 34
rect 976 32 978 34
rect 981 32 983 34
rect 986 32 988 34
rect 991 32 993 34
rect 996 32 998 34
rect 331 26 333 28
rect 336 26 338 28
rect 341 26 343 28
rect 346 26 348 28
rect 351 26 353 28
rect 356 26 358 28
rect 361 26 363 28
rect 366 26 368 28
rect 371 26 373 28
rect 376 26 378 28
rect 381 26 383 28
rect 386 26 388 28
rect 391 26 393 28
rect 396 26 398 28
rect 401 26 403 28
rect 406 26 408 28
rect 411 26 413 28
rect 416 26 418 28
rect 421 26 423 28
rect 426 26 428 28
rect 431 26 433 28
rect 436 26 438 28
rect 441 26 443 28
rect 446 26 448 28
rect 451 26 453 28
rect 456 26 458 28
rect 461 26 463 28
rect 466 26 468 28
rect 471 26 473 28
rect 476 26 478 28
rect 481 26 483 28
rect 486 26 488 28
rect 491 26 493 28
rect 496 26 498 28
rect 501 26 503 28
rect 506 26 508 28
rect 511 26 513 28
rect 516 26 518 28
rect 521 26 523 28
rect 526 26 528 28
rect 531 26 533 28
rect 536 26 538 28
rect 541 26 543 28
rect 546 26 548 28
rect 551 26 553 28
rect 556 26 558 28
rect 771 27 773 29
rect 776 27 778 29
rect 781 27 783 29
rect 786 27 788 29
rect 791 27 793 29
rect 796 27 798 29
rect 801 27 803 29
rect 806 27 808 29
rect 811 27 813 29
rect 816 27 818 29
rect 821 27 823 29
rect 826 27 828 29
rect 831 27 833 29
rect 836 27 838 29
rect 841 27 843 29
rect 846 27 848 29
rect 851 27 853 29
rect 856 27 858 29
rect 861 27 863 29
rect 866 27 868 29
rect 871 27 873 29
rect 876 27 878 29
rect 881 27 883 29
rect 886 27 888 29
rect 891 27 893 29
rect 896 27 898 29
rect 901 27 903 29
rect 906 27 908 29
rect 911 27 913 29
rect 916 27 918 29
rect 921 27 923 29
rect 926 27 928 29
rect 931 27 933 29
rect 936 27 938 29
rect 941 27 943 29
rect 946 27 948 29
rect 951 27 953 29
rect 956 27 958 29
rect 961 27 963 29
rect 966 27 968 29
rect 971 27 973 29
rect 976 27 978 29
rect 981 27 983 29
rect 986 27 988 29
rect 991 27 993 29
rect 996 27 998 29
rect 331 21 333 23
rect 336 21 338 23
rect 341 21 343 23
rect 346 21 348 23
rect 351 21 353 23
rect 356 21 358 23
rect 361 21 363 23
rect 366 21 368 23
rect 371 21 373 23
rect 376 21 378 23
rect 381 21 383 23
rect 386 21 388 23
rect 391 21 393 23
rect 396 21 398 23
rect 401 21 403 23
rect 406 21 408 23
rect 411 21 413 23
rect 416 21 418 23
rect 421 21 423 23
rect 426 21 428 23
rect 431 21 433 23
rect 436 21 438 23
rect 441 21 443 23
rect 446 21 448 23
rect 451 21 453 23
rect 456 21 458 23
rect 461 21 463 23
rect 466 21 468 23
rect 471 21 473 23
rect 476 21 478 23
rect 481 21 483 23
rect 486 21 488 23
rect 491 21 493 23
rect 496 21 498 23
rect 501 21 503 23
rect 506 21 508 23
rect 511 21 513 23
rect 516 21 518 23
rect 521 21 523 23
rect 526 21 528 23
rect 531 21 533 23
rect 536 21 538 23
rect 541 21 543 23
rect 546 21 548 23
rect 551 21 553 23
rect 556 21 558 23
rect 771 22 773 24
rect 776 22 778 24
rect 781 22 783 24
rect 786 22 788 24
rect 791 22 793 24
rect 796 22 798 24
rect 801 22 803 24
rect 806 22 808 24
rect 811 22 813 24
rect 816 22 818 24
rect 821 22 823 24
rect 826 22 828 24
rect 831 22 833 24
rect 836 22 838 24
rect 841 22 843 24
rect 846 22 848 24
rect 851 22 853 24
rect 856 22 858 24
rect 861 22 863 24
rect 866 22 868 24
rect 871 22 873 24
rect 876 22 878 24
rect 881 22 883 24
rect 886 22 888 24
rect 891 22 893 24
rect 896 22 898 24
rect 901 22 903 24
rect 906 22 908 24
rect 911 22 913 24
rect 916 22 918 24
rect 921 22 923 24
rect 926 22 928 24
rect 931 22 933 24
rect 936 22 938 24
rect 941 22 943 24
rect 946 22 948 24
rect 951 22 953 24
rect 956 22 958 24
rect 961 22 963 24
rect 966 22 968 24
rect 971 22 973 24
rect 976 22 978 24
rect 981 22 983 24
rect 986 22 988 24
rect 991 22 993 24
rect 996 22 998 24
rect 331 16 333 18
rect 336 16 338 18
rect 341 16 343 18
rect 346 16 348 18
rect 351 16 353 18
rect 356 16 358 18
rect 361 16 363 18
rect 366 16 368 18
rect 371 16 373 18
rect 376 16 378 18
rect 381 16 383 18
rect 386 16 388 18
rect 391 16 393 18
rect 396 16 398 18
rect 401 16 403 18
rect 406 16 408 18
rect 411 16 413 18
rect 416 16 418 18
rect 421 16 423 18
rect 426 16 428 18
rect 431 16 433 18
rect 436 16 438 18
rect 441 16 443 18
rect 446 16 448 18
rect 451 16 453 18
rect 456 16 458 18
rect 461 16 463 18
rect 466 16 468 18
rect 471 16 473 18
rect 476 16 478 18
rect 481 16 483 18
rect 486 16 488 18
rect 491 16 493 18
rect 496 16 498 18
rect 501 16 503 18
rect 506 16 508 18
rect 511 16 513 18
rect 516 16 518 18
rect 521 16 523 18
rect 526 16 528 18
rect 531 16 533 18
rect 536 16 538 18
rect 541 16 543 18
rect 546 16 548 18
rect 551 16 553 18
rect 556 16 558 18
rect 771 17 773 19
rect 776 17 778 19
rect 781 17 783 19
rect 786 17 788 19
rect 791 17 793 19
rect 796 17 798 19
rect 801 17 803 19
rect 806 17 808 19
rect 811 17 813 19
rect 816 17 818 19
rect 821 17 823 19
rect 826 17 828 19
rect 831 17 833 19
rect 836 17 838 19
rect 841 17 843 19
rect 846 17 848 19
rect 851 17 853 19
rect 856 17 858 19
rect 861 17 863 19
rect 866 17 868 19
rect 871 17 873 19
rect 876 17 878 19
rect 881 17 883 19
rect 886 17 888 19
rect 891 17 893 19
rect 896 17 898 19
rect 901 17 903 19
rect 906 17 908 19
rect 911 17 913 19
rect 916 17 918 19
rect 921 17 923 19
rect 926 17 928 19
rect 931 17 933 19
rect 936 17 938 19
rect 941 17 943 19
rect 946 17 948 19
rect 951 17 953 19
rect 956 17 958 19
rect 961 17 963 19
rect 966 17 968 19
rect 971 17 973 19
rect 976 17 978 19
rect 981 17 983 19
rect 986 17 988 19
rect 991 17 993 19
rect 996 17 998 19
rect 331 11 333 13
rect 336 11 338 13
rect 341 11 343 13
rect 346 11 348 13
rect 351 11 353 13
rect 356 11 358 13
rect 361 11 363 13
rect 366 11 368 13
rect 371 11 373 13
rect 376 11 378 13
rect 381 11 383 13
rect 386 11 388 13
rect 391 11 393 13
rect 396 11 398 13
rect 401 11 403 13
rect 406 11 408 13
rect 411 11 413 13
rect 416 11 418 13
rect 421 11 423 13
rect 426 11 428 13
rect 431 11 433 13
rect 436 11 438 13
rect 441 11 443 13
rect 446 11 448 13
rect 451 11 453 13
rect 456 11 458 13
rect 461 11 463 13
rect 466 11 468 13
rect 471 11 473 13
rect 476 11 478 13
rect 481 11 483 13
rect 486 11 488 13
rect 491 11 493 13
rect 496 11 498 13
rect 501 11 503 13
rect 506 11 508 13
rect 511 11 513 13
rect 516 11 518 13
rect 521 11 523 13
rect 526 11 528 13
rect 531 11 533 13
rect 536 11 538 13
rect 541 11 543 13
rect 546 11 548 13
rect 551 11 553 13
rect 556 11 558 13
rect 771 12 773 14
rect 776 12 778 14
rect 781 12 783 14
rect 786 12 788 14
rect 791 12 793 14
rect 796 12 798 14
rect 801 12 803 14
rect 806 12 808 14
rect 811 12 813 14
rect 816 12 818 14
rect 821 12 823 14
rect 826 12 828 14
rect 831 12 833 14
rect 836 12 838 14
rect 841 12 843 14
rect 846 12 848 14
rect 851 12 853 14
rect 856 12 858 14
rect 861 12 863 14
rect 866 12 868 14
rect 871 12 873 14
rect 876 12 878 14
rect 881 12 883 14
rect 886 12 888 14
rect 891 12 893 14
rect 896 12 898 14
rect 901 12 903 14
rect 906 12 908 14
rect 911 12 913 14
rect 916 12 918 14
rect 921 12 923 14
rect 926 12 928 14
rect 931 12 933 14
rect 936 12 938 14
rect 941 12 943 14
rect 946 12 948 14
rect 951 12 953 14
rect 956 12 958 14
rect 961 12 963 14
rect 966 12 968 14
rect 971 12 973 14
rect 976 12 978 14
rect 981 12 983 14
rect 986 12 988 14
rect 991 12 993 14
rect 996 12 998 14
rect 331 6 333 8
rect 336 6 338 8
rect 341 6 343 8
rect 346 6 348 8
rect 351 6 353 8
rect 356 6 358 8
rect 361 6 363 8
rect 366 6 368 8
rect 371 6 373 8
rect 376 6 378 8
rect 381 6 383 8
rect 386 6 388 8
rect 391 6 393 8
rect 396 6 398 8
rect 401 6 403 8
rect 406 6 408 8
rect 411 6 413 8
rect 416 6 418 8
rect 421 6 423 8
rect 426 6 428 8
rect 431 6 433 8
rect 436 6 438 8
rect 441 6 443 8
rect 446 6 448 8
rect 451 6 453 8
rect 456 6 458 8
rect 461 6 463 8
rect 466 6 468 8
rect 471 6 473 8
rect 476 6 478 8
rect 481 6 483 8
rect 486 6 488 8
rect 491 6 493 8
rect 496 6 498 8
rect 501 6 503 8
rect 506 6 508 8
rect 511 6 513 8
rect 516 6 518 8
rect 521 6 523 8
rect 526 6 528 8
rect 531 6 533 8
rect 536 6 538 8
rect 541 6 543 8
rect 546 6 548 8
rect 551 6 553 8
rect 556 6 558 8
rect 771 7 773 9
rect 776 7 778 9
rect 781 7 783 9
rect 786 7 788 9
rect 791 7 793 9
rect 796 7 798 9
rect 801 7 803 9
rect 806 7 808 9
rect 811 7 813 9
rect 816 7 818 9
rect 821 7 823 9
rect 826 7 828 9
rect 831 7 833 9
rect 836 7 838 9
rect 841 7 843 9
rect 846 7 848 9
rect 851 7 853 9
rect 856 7 858 9
rect 861 7 863 9
rect 866 7 868 9
rect 871 7 873 9
rect 876 7 878 9
rect 881 7 883 9
rect 886 7 888 9
rect 891 7 893 9
rect 896 7 898 9
rect 901 7 903 9
rect 906 7 908 9
rect 911 7 913 9
rect 916 7 918 9
rect 921 7 923 9
rect 926 7 928 9
rect 931 7 933 9
rect 936 7 938 9
rect 941 7 943 9
rect 946 7 948 9
rect 951 7 953 9
rect 956 7 958 9
rect 961 7 963 9
rect 966 7 968 9
rect 971 7 973 9
rect 976 7 978 9
rect 981 7 983 9
rect 986 7 988 9
rect 991 7 993 9
rect 996 7 998 9
rect 331 1 333 3
rect 336 1 338 3
rect 341 1 343 3
rect 346 1 348 3
rect 351 1 353 3
rect 356 1 358 3
rect 361 1 363 3
rect 366 1 368 3
rect 371 1 373 3
rect 376 1 378 3
rect 381 1 383 3
rect 386 1 388 3
rect 391 1 393 3
rect 396 1 398 3
rect 401 1 403 3
rect 406 1 408 3
rect 411 1 413 3
rect 416 1 418 3
rect 421 1 423 3
rect 426 1 428 3
rect 431 1 433 3
rect 436 1 438 3
rect 441 1 443 3
rect 446 1 448 3
rect 451 1 453 3
rect 456 1 458 3
rect 461 1 463 3
rect 466 1 468 3
rect 471 1 473 3
rect 476 1 478 3
rect 481 1 483 3
rect 486 1 488 3
rect 491 1 493 3
rect 496 1 498 3
rect 501 1 503 3
rect 506 1 508 3
rect 511 1 513 3
rect 516 1 518 3
rect 521 1 523 3
rect 526 1 528 3
rect 531 1 533 3
rect 536 1 538 3
rect 541 1 543 3
rect 546 1 548 3
rect 551 1 553 3
rect 556 1 558 3
rect 771 2 773 4
rect 776 2 778 4
rect 781 2 783 4
rect 786 2 788 4
rect 791 2 793 4
rect 796 2 798 4
rect 801 2 803 4
rect 806 2 808 4
rect 811 2 813 4
rect 816 2 818 4
rect 821 2 823 4
rect 826 2 828 4
rect 831 2 833 4
rect 836 2 838 4
rect 841 2 843 4
rect 846 2 848 4
rect 851 2 853 4
rect 856 2 858 4
rect 861 2 863 4
rect 866 2 868 4
rect 871 2 873 4
rect 876 2 878 4
rect 881 2 883 4
rect 886 2 888 4
rect 891 2 893 4
rect 896 2 898 4
rect 901 2 903 4
rect 906 2 908 4
rect 911 2 913 4
rect 916 2 918 4
rect 921 2 923 4
rect 926 2 928 4
rect 931 2 933 4
rect 936 2 938 4
rect 941 2 943 4
rect 946 2 948 4
rect 951 2 953 4
rect 956 2 958 4
rect 961 2 963 4
rect 966 2 968 4
rect 971 2 973 4
rect 976 2 978 4
rect 981 2 983 4
rect 986 2 988 4
rect 991 2 993 4
rect 996 2 998 4
<< metal1 >>
rect 330 344 1000 670
rect 330 0 655 344
rect 674 0 1000 327
<< metal2 >>
rect 330 441 1000 670
rect 330 0 560 441
rect 576 344 1000 423
rect 576 0 655 344
rect 674 246 1000 327
rect 674 0 753 246
rect 769 0 1000 230
<< gv1 >>
rect 577 420 579 422
rect 582 420 584 422
rect 587 420 589 422
rect 592 420 594 422
rect 597 420 599 422
rect 602 420 604 422
rect 607 420 609 422
rect 612 420 614 422
rect 617 420 619 422
rect 622 420 624 422
rect 627 420 629 422
rect 632 420 634 422
rect 637 420 639 422
rect 642 420 644 422
rect 647 420 649 422
rect 652 420 654 422
rect 657 420 659 422
rect 662 420 664 422
rect 667 420 669 422
rect 672 420 674 422
rect 677 420 679 422
rect 682 420 684 422
rect 687 420 689 422
rect 692 420 694 422
rect 697 420 699 422
rect 702 420 704 422
rect 707 420 709 422
rect 712 420 714 422
rect 717 420 719 422
rect 722 420 724 422
rect 727 420 729 422
rect 732 420 734 422
rect 737 420 739 422
rect 742 420 744 422
rect 747 420 749 422
rect 752 420 754 422
rect 757 420 759 422
rect 762 420 764 422
rect 767 420 769 422
rect 772 420 774 422
rect 777 420 779 422
rect 782 420 784 422
rect 787 420 789 422
rect 792 420 794 422
rect 797 420 799 422
rect 802 420 804 422
rect 807 420 809 422
rect 812 420 814 422
rect 817 420 819 422
rect 822 420 824 422
rect 827 420 829 422
rect 832 420 834 422
rect 837 420 839 422
rect 842 420 844 422
rect 847 420 849 422
rect 852 420 854 422
rect 857 420 859 422
rect 862 420 864 422
rect 867 420 869 422
rect 872 420 874 422
rect 877 420 879 422
rect 882 420 884 422
rect 887 420 889 422
rect 892 420 894 422
rect 897 420 899 422
rect 902 420 904 422
rect 907 420 909 422
rect 912 420 914 422
rect 917 420 919 422
rect 922 420 924 422
rect 927 420 929 422
rect 932 420 934 422
rect 937 420 939 422
rect 942 420 944 422
rect 947 420 949 422
rect 952 420 954 422
rect 957 420 959 422
rect 962 420 964 422
rect 967 420 969 422
rect 972 420 974 422
rect 977 420 979 422
rect 982 420 984 422
rect 987 420 989 422
rect 992 420 994 422
rect 997 420 999 422
rect 577 415 579 417
rect 582 415 584 417
rect 587 415 589 417
rect 592 415 594 417
rect 597 415 599 417
rect 602 415 604 417
rect 607 415 609 417
rect 612 415 614 417
rect 617 415 619 417
rect 622 415 624 417
rect 627 415 629 417
rect 632 415 634 417
rect 637 415 639 417
rect 642 415 644 417
rect 647 415 649 417
rect 652 415 654 417
rect 657 415 659 417
rect 662 415 664 417
rect 667 415 669 417
rect 672 415 674 417
rect 677 415 679 417
rect 682 415 684 417
rect 687 415 689 417
rect 692 415 694 417
rect 697 415 699 417
rect 702 415 704 417
rect 707 415 709 417
rect 712 415 714 417
rect 717 415 719 417
rect 722 415 724 417
rect 727 415 729 417
rect 732 415 734 417
rect 737 415 739 417
rect 742 415 744 417
rect 747 415 749 417
rect 752 415 754 417
rect 757 415 759 417
rect 762 415 764 417
rect 767 415 769 417
rect 772 415 774 417
rect 777 415 779 417
rect 782 415 784 417
rect 787 415 789 417
rect 792 415 794 417
rect 797 415 799 417
rect 802 415 804 417
rect 807 415 809 417
rect 812 415 814 417
rect 817 415 819 417
rect 822 415 824 417
rect 827 415 829 417
rect 832 415 834 417
rect 837 415 839 417
rect 842 415 844 417
rect 847 415 849 417
rect 852 415 854 417
rect 857 415 859 417
rect 862 415 864 417
rect 867 415 869 417
rect 872 415 874 417
rect 877 415 879 417
rect 882 415 884 417
rect 887 415 889 417
rect 892 415 894 417
rect 897 415 899 417
rect 902 415 904 417
rect 907 415 909 417
rect 912 415 914 417
rect 917 415 919 417
rect 922 415 924 417
rect 927 415 929 417
rect 932 415 934 417
rect 937 415 939 417
rect 942 415 944 417
rect 947 415 949 417
rect 952 415 954 417
rect 957 415 959 417
rect 962 415 964 417
rect 967 415 969 417
rect 972 415 974 417
rect 977 415 979 417
rect 982 415 984 417
rect 987 415 989 417
rect 992 415 994 417
rect 997 415 999 417
rect 577 410 579 412
rect 582 410 584 412
rect 587 410 589 412
rect 592 410 594 412
rect 597 410 599 412
rect 602 410 604 412
rect 607 410 609 412
rect 612 410 614 412
rect 617 410 619 412
rect 622 410 624 412
rect 627 410 629 412
rect 632 410 634 412
rect 637 410 639 412
rect 642 410 644 412
rect 647 410 649 412
rect 652 410 654 412
rect 657 410 659 412
rect 662 410 664 412
rect 667 410 669 412
rect 672 410 674 412
rect 677 410 679 412
rect 682 410 684 412
rect 687 410 689 412
rect 692 410 694 412
rect 697 410 699 412
rect 702 410 704 412
rect 707 410 709 412
rect 712 410 714 412
rect 717 410 719 412
rect 722 410 724 412
rect 727 410 729 412
rect 732 410 734 412
rect 737 410 739 412
rect 742 410 744 412
rect 747 410 749 412
rect 752 410 754 412
rect 757 410 759 412
rect 762 410 764 412
rect 767 410 769 412
rect 772 410 774 412
rect 777 410 779 412
rect 782 410 784 412
rect 787 410 789 412
rect 792 410 794 412
rect 797 410 799 412
rect 802 410 804 412
rect 807 410 809 412
rect 812 410 814 412
rect 817 410 819 412
rect 822 410 824 412
rect 827 410 829 412
rect 832 410 834 412
rect 837 410 839 412
rect 842 410 844 412
rect 847 410 849 412
rect 852 410 854 412
rect 857 410 859 412
rect 862 410 864 412
rect 867 410 869 412
rect 872 410 874 412
rect 877 410 879 412
rect 882 410 884 412
rect 887 410 889 412
rect 892 410 894 412
rect 897 410 899 412
rect 902 410 904 412
rect 907 410 909 412
rect 912 410 914 412
rect 917 410 919 412
rect 922 410 924 412
rect 927 410 929 412
rect 932 410 934 412
rect 937 410 939 412
rect 942 410 944 412
rect 947 410 949 412
rect 952 410 954 412
rect 957 410 959 412
rect 962 410 964 412
rect 967 410 969 412
rect 972 410 974 412
rect 977 410 979 412
rect 982 410 984 412
rect 987 410 989 412
rect 992 410 994 412
rect 997 410 999 412
rect 577 405 579 407
rect 582 405 584 407
rect 587 405 589 407
rect 592 405 594 407
rect 597 405 599 407
rect 602 405 604 407
rect 607 405 609 407
rect 612 405 614 407
rect 617 405 619 407
rect 622 405 624 407
rect 627 405 629 407
rect 632 405 634 407
rect 637 405 639 407
rect 642 405 644 407
rect 647 405 649 407
rect 652 405 654 407
rect 657 405 659 407
rect 662 405 664 407
rect 667 405 669 407
rect 672 405 674 407
rect 677 405 679 407
rect 682 405 684 407
rect 687 405 689 407
rect 692 405 694 407
rect 697 405 699 407
rect 702 405 704 407
rect 707 405 709 407
rect 712 405 714 407
rect 717 405 719 407
rect 722 405 724 407
rect 727 405 729 407
rect 732 405 734 407
rect 737 405 739 407
rect 742 405 744 407
rect 747 405 749 407
rect 752 405 754 407
rect 757 405 759 407
rect 762 405 764 407
rect 767 405 769 407
rect 772 405 774 407
rect 777 405 779 407
rect 782 405 784 407
rect 787 405 789 407
rect 792 405 794 407
rect 797 405 799 407
rect 802 405 804 407
rect 807 405 809 407
rect 812 405 814 407
rect 817 405 819 407
rect 822 405 824 407
rect 827 405 829 407
rect 832 405 834 407
rect 837 405 839 407
rect 842 405 844 407
rect 847 405 849 407
rect 852 405 854 407
rect 857 405 859 407
rect 862 405 864 407
rect 867 405 869 407
rect 872 405 874 407
rect 877 405 879 407
rect 882 405 884 407
rect 887 405 889 407
rect 892 405 894 407
rect 897 405 899 407
rect 902 405 904 407
rect 907 405 909 407
rect 912 405 914 407
rect 917 405 919 407
rect 922 405 924 407
rect 927 405 929 407
rect 932 405 934 407
rect 937 405 939 407
rect 942 405 944 407
rect 947 405 949 407
rect 952 405 954 407
rect 957 405 959 407
rect 962 405 964 407
rect 967 405 969 407
rect 972 405 974 407
rect 977 405 979 407
rect 982 405 984 407
rect 987 405 989 407
rect 992 405 994 407
rect 997 405 999 407
rect 577 400 579 402
rect 582 400 584 402
rect 587 400 589 402
rect 592 400 594 402
rect 597 400 599 402
rect 602 400 604 402
rect 607 400 609 402
rect 612 400 614 402
rect 617 400 619 402
rect 622 400 624 402
rect 627 400 629 402
rect 632 400 634 402
rect 637 400 639 402
rect 642 400 644 402
rect 647 400 649 402
rect 652 400 654 402
rect 657 400 659 402
rect 662 400 664 402
rect 667 400 669 402
rect 672 400 674 402
rect 677 400 679 402
rect 682 400 684 402
rect 687 400 689 402
rect 692 400 694 402
rect 697 400 699 402
rect 702 400 704 402
rect 707 400 709 402
rect 712 400 714 402
rect 717 400 719 402
rect 722 400 724 402
rect 727 400 729 402
rect 732 400 734 402
rect 737 400 739 402
rect 742 400 744 402
rect 747 400 749 402
rect 752 400 754 402
rect 757 400 759 402
rect 762 400 764 402
rect 767 400 769 402
rect 772 400 774 402
rect 777 400 779 402
rect 782 400 784 402
rect 787 400 789 402
rect 792 400 794 402
rect 797 400 799 402
rect 802 400 804 402
rect 807 400 809 402
rect 812 400 814 402
rect 817 400 819 402
rect 822 400 824 402
rect 827 400 829 402
rect 832 400 834 402
rect 837 400 839 402
rect 842 400 844 402
rect 847 400 849 402
rect 852 400 854 402
rect 857 400 859 402
rect 862 400 864 402
rect 867 400 869 402
rect 872 400 874 402
rect 877 400 879 402
rect 882 400 884 402
rect 887 400 889 402
rect 892 400 894 402
rect 897 400 899 402
rect 902 400 904 402
rect 907 400 909 402
rect 912 400 914 402
rect 917 400 919 402
rect 922 400 924 402
rect 927 400 929 402
rect 932 400 934 402
rect 937 400 939 402
rect 942 400 944 402
rect 947 400 949 402
rect 952 400 954 402
rect 957 400 959 402
rect 962 400 964 402
rect 967 400 969 402
rect 972 400 974 402
rect 977 400 979 402
rect 982 400 984 402
rect 987 400 989 402
rect 992 400 994 402
rect 997 400 999 402
rect 577 395 579 397
rect 582 395 584 397
rect 587 395 589 397
rect 592 395 594 397
rect 597 395 599 397
rect 602 395 604 397
rect 607 395 609 397
rect 612 395 614 397
rect 617 395 619 397
rect 622 395 624 397
rect 627 395 629 397
rect 632 395 634 397
rect 637 395 639 397
rect 642 395 644 397
rect 647 395 649 397
rect 652 395 654 397
rect 657 395 659 397
rect 662 395 664 397
rect 667 395 669 397
rect 672 395 674 397
rect 677 395 679 397
rect 682 395 684 397
rect 687 395 689 397
rect 692 395 694 397
rect 697 395 699 397
rect 702 395 704 397
rect 707 395 709 397
rect 712 395 714 397
rect 717 395 719 397
rect 722 395 724 397
rect 727 395 729 397
rect 732 395 734 397
rect 737 395 739 397
rect 742 395 744 397
rect 747 395 749 397
rect 752 395 754 397
rect 757 395 759 397
rect 762 395 764 397
rect 767 395 769 397
rect 772 395 774 397
rect 777 395 779 397
rect 782 395 784 397
rect 787 395 789 397
rect 792 395 794 397
rect 797 395 799 397
rect 802 395 804 397
rect 807 395 809 397
rect 812 395 814 397
rect 817 395 819 397
rect 822 395 824 397
rect 827 395 829 397
rect 832 395 834 397
rect 837 395 839 397
rect 842 395 844 397
rect 847 395 849 397
rect 852 395 854 397
rect 857 395 859 397
rect 862 395 864 397
rect 867 395 869 397
rect 872 395 874 397
rect 877 395 879 397
rect 882 395 884 397
rect 887 395 889 397
rect 892 395 894 397
rect 897 395 899 397
rect 902 395 904 397
rect 907 395 909 397
rect 912 395 914 397
rect 917 395 919 397
rect 922 395 924 397
rect 927 395 929 397
rect 932 395 934 397
rect 937 395 939 397
rect 942 395 944 397
rect 947 395 949 397
rect 952 395 954 397
rect 957 395 959 397
rect 962 395 964 397
rect 967 395 969 397
rect 972 395 974 397
rect 977 395 979 397
rect 982 395 984 397
rect 987 395 989 397
rect 992 395 994 397
rect 997 395 999 397
rect 577 390 579 392
rect 582 390 584 392
rect 587 390 589 392
rect 592 390 594 392
rect 597 390 599 392
rect 602 390 604 392
rect 607 390 609 392
rect 612 390 614 392
rect 617 390 619 392
rect 622 390 624 392
rect 627 390 629 392
rect 632 390 634 392
rect 637 390 639 392
rect 642 390 644 392
rect 647 390 649 392
rect 652 390 654 392
rect 657 390 659 392
rect 662 390 664 392
rect 667 390 669 392
rect 672 390 674 392
rect 677 390 679 392
rect 682 390 684 392
rect 687 390 689 392
rect 692 390 694 392
rect 697 390 699 392
rect 702 390 704 392
rect 707 390 709 392
rect 712 390 714 392
rect 717 390 719 392
rect 722 390 724 392
rect 727 390 729 392
rect 732 390 734 392
rect 737 390 739 392
rect 742 390 744 392
rect 747 390 749 392
rect 752 390 754 392
rect 757 390 759 392
rect 762 390 764 392
rect 767 390 769 392
rect 772 390 774 392
rect 777 390 779 392
rect 782 390 784 392
rect 787 390 789 392
rect 792 390 794 392
rect 797 390 799 392
rect 802 390 804 392
rect 807 390 809 392
rect 812 390 814 392
rect 817 390 819 392
rect 822 390 824 392
rect 827 390 829 392
rect 832 390 834 392
rect 837 390 839 392
rect 842 390 844 392
rect 847 390 849 392
rect 852 390 854 392
rect 857 390 859 392
rect 862 390 864 392
rect 867 390 869 392
rect 872 390 874 392
rect 877 390 879 392
rect 882 390 884 392
rect 887 390 889 392
rect 892 390 894 392
rect 897 390 899 392
rect 902 390 904 392
rect 907 390 909 392
rect 912 390 914 392
rect 917 390 919 392
rect 922 390 924 392
rect 927 390 929 392
rect 932 390 934 392
rect 937 390 939 392
rect 942 390 944 392
rect 947 390 949 392
rect 952 390 954 392
rect 957 390 959 392
rect 962 390 964 392
rect 967 390 969 392
rect 972 390 974 392
rect 977 390 979 392
rect 982 390 984 392
rect 987 390 989 392
rect 992 390 994 392
rect 997 390 999 392
rect 577 385 579 387
rect 582 385 584 387
rect 587 385 589 387
rect 592 385 594 387
rect 597 385 599 387
rect 602 385 604 387
rect 607 385 609 387
rect 612 385 614 387
rect 617 385 619 387
rect 622 385 624 387
rect 627 385 629 387
rect 632 385 634 387
rect 637 385 639 387
rect 642 385 644 387
rect 647 385 649 387
rect 652 385 654 387
rect 657 385 659 387
rect 662 385 664 387
rect 667 385 669 387
rect 672 385 674 387
rect 677 385 679 387
rect 682 385 684 387
rect 687 385 689 387
rect 692 385 694 387
rect 697 385 699 387
rect 702 385 704 387
rect 707 385 709 387
rect 712 385 714 387
rect 717 385 719 387
rect 722 385 724 387
rect 727 385 729 387
rect 732 385 734 387
rect 737 385 739 387
rect 742 385 744 387
rect 747 385 749 387
rect 752 385 754 387
rect 757 385 759 387
rect 762 385 764 387
rect 767 385 769 387
rect 772 385 774 387
rect 777 385 779 387
rect 782 385 784 387
rect 787 385 789 387
rect 792 385 794 387
rect 797 385 799 387
rect 802 385 804 387
rect 807 385 809 387
rect 812 385 814 387
rect 817 385 819 387
rect 822 385 824 387
rect 827 385 829 387
rect 832 385 834 387
rect 837 385 839 387
rect 842 385 844 387
rect 847 385 849 387
rect 852 385 854 387
rect 857 385 859 387
rect 862 385 864 387
rect 867 385 869 387
rect 872 385 874 387
rect 877 385 879 387
rect 882 385 884 387
rect 887 385 889 387
rect 892 385 894 387
rect 897 385 899 387
rect 902 385 904 387
rect 907 385 909 387
rect 912 385 914 387
rect 917 385 919 387
rect 922 385 924 387
rect 927 385 929 387
rect 932 385 934 387
rect 937 385 939 387
rect 942 385 944 387
rect 947 385 949 387
rect 952 385 954 387
rect 957 385 959 387
rect 962 385 964 387
rect 967 385 969 387
rect 972 385 974 387
rect 977 385 979 387
rect 982 385 984 387
rect 987 385 989 387
rect 992 385 994 387
rect 997 385 999 387
rect 577 380 579 382
rect 582 380 584 382
rect 587 380 589 382
rect 592 380 594 382
rect 597 380 599 382
rect 602 380 604 382
rect 607 380 609 382
rect 612 380 614 382
rect 617 380 619 382
rect 622 380 624 382
rect 627 380 629 382
rect 632 380 634 382
rect 637 380 639 382
rect 642 380 644 382
rect 647 380 649 382
rect 652 380 654 382
rect 657 380 659 382
rect 662 380 664 382
rect 667 380 669 382
rect 672 380 674 382
rect 677 380 679 382
rect 682 380 684 382
rect 687 380 689 382
rect 692 380 694 382
rect 697 380 699 382
rect 702 380 704 382
rect 707 380 709 382
rect 712 380 714 382
rect 717 380 719 382
rect 722 380 724 382
rect 727 380 729 382
rect 732 380 734 382
rect 737 380 739 382
rect 742 380 744 382
rect 747 380 749 382
rect 752 380 754 382
rect 757 380 759 382
rect 762 380 764 382
rect 767 380 769 382
rect 772 380 774 382
rect 777 380 779 382
rect 782 380 784 382
rect 787 380 789 382
rect 792 380 794 382
rect 797 380 799 382
rect 802 380 804 382
rect 807 380 809 382
rect 812 380 814 382
rect 817 380 819 382
rect 822 380 824 382
rect 827 380 829 382
rect 832 380 834 382
rect 837 380 839 382
rect 842 380 844 382
rect 847 380 849 382
rect 852 380 854 382
rect 857 380 859 382
rect 862 380 864 382
rect 867 380 869 382
rect 872 380 874 382
rect 877 380 879 382
rect 882 380 884 382
rect 887 380 889 382
rect 892 380 894 382
rect 897 380 899 382
rect 902 380 904 382
rect 907 380 909 382
rect 912 380 914 382
rect 917 380 919 382
rect 922 380 924 382
rect 927 380 929 382
rect 932 380 934 382
rect 937 380 939 382
rect 942 380 944 382
rect 947 380 949 382
rect 952 380 954 382
rect 957 380 959 382
rect 962 380 964 382
rect 967 380 969 382
rect 972 380 974 382
rect 977 380 979 382
rect 982 380 984 382
rect 987 380 989 382
rect 992 380 994 382
rect 997 380 999 382
rect 577 375 579 377
rect 582 375 584 377
rect 587 375 589 377
rect 592 375 594 377
rect 597 375 599 377
rect 602 375 604 377
rect 607 375 609 377
rect 612 375 614 377
rect 617 375 619 377
rect 622 375 624 377
rect 627 375 629 377
rect 632 375 634 377
rect 637 375 639 377
rect 642 375 644 377
rect 647 375 649 377
rect 652 375 654 377
rect 657 375 659 377
rect 662 375 664 377
rect 667 375 669 377
rect 672 375 674 377
rect 677 375 679 377
rect 682 375 684 377
rect 687 375 689 377
rect 692 375 694 377
rect 697 375 699 377
rect 702 375 704 377
rect 707 375 709 377
rect 712 375 714 377
rect 717 375 719 377
rect 722 375 724 377
rect 727 375 729 377
rect 732 375 734 377
rect 737 375 739 377
rect 742 375 744 377
rect 747 375 749 377
rect 752 375 754 377
rect 757 375 759 377
rect 762 375 764 377
rect 767 375 769 377
rect 772 375 774 377
rect 777 375 779 377
rect 782 375 784 377
rect 787 375 789 377
rect 792 375 794 377
rect 797 375 799 377
rect 802 375 804 377
rect 807 375 809 377
rect 812 375 814 377
rect 817 375 819 377
rect 822 375 824 377
rect 827 375 829 377
rect 832 375 834 377
rect 837 375 839 377
rect 842 375 844 377
rect 847 375 849 377
rect 852 375 854 377
rect 857 375 859 377
rect 862 375 864 377
rect 867 375 869 377
rect 872 375 874 377
rect 877 375 879 377
rect 882 375 884 377
rect 887 375 889 377
rect 892 375 894 377
rect 897 375 899 377
rect 902 375 904 377
rect 907 375 909 377
rect 912 375 914 377
rect 917 375 919 377
rect 922 375 924 377
rect 927 375 929 377
rect 932 375 934 377
rect 937 375 939 377
rect 942 375 944 377
rect 947 375 949 377
rect 952 375 954 377
rect 957 375 959 377
rect 962 375 964 377
rect 967 375 969 377
rect 972 375 974 377
rect 977 375 979 377
rect 982 375 984 377
rect 987 375 989 377
rect 992 375 994 377
rect 997 375 999 377
rect 577 370 579 372
rect 582 370 584 372
rect 587 370 589 372
rect 592 370 594 372
rect 597 370 599 372
rect 602 370 604 372
rect 607 370 609 372
rect 612 370 614 372
rect 617 370 619 372
rect 622 370 624 372
rect 627 370 629 372
rect 632 370 634 372
rect 637 370 639 372
rect 642 370 644 372
rect 647 370 649 372
rect 652 370 654 372
rect 657 370 659 372
rect 662 370 664 372
rect 667 370 669 372
rect 672 370 674 372
rect 677 370 679 372
rect 682 370 684 372
rect 687 370 689 372
rect 692 370 694 372
rect 697 370 699 372
rect 702 370 704 372
rect 707 370 709 372
rect 712 370 714 372
rect 717 370 719 372
rect 722 370 724 372
rect 727 370 729 372
rect 732 370 734 372
rect 737 370 739 372
rect 742 370 744 372
rect 747 370 749 372
rect 752 370 754 372
rect 757 370 759 372
rect 762 370 764 372
rect 767 370 769 372
rect 772 370 774 372
rect 777 370 779 372
rect 782 370 784 372
rect 787 370 789 372
rect 792 370 794 372
rect 797 370 799 372
rect 802 370 804 372
rect 807 370 809 372
rect 812 370 814 372
rect 817 370 819 372
rect 822 370 824 372
rect 827 370 829 372
rect 832 370 834 372
rect 837 370 839 372
rect 842 370 844 372
rect 847 370 849 372
rect 852 370 854 372
rect 857 370 859 372
rect 862 370 864 372
rect 867 370 869 372
rect 872 370 874 372
rect 877 370 879 372
rect 882 370 884 372
rect 887 370 889 372
rect 892 370 894 372
rect 897 370 899 372
rect 902 370 904 372
rect 907 370 909 372
rect 912 370 914 372
rect 917 370 919 372
rect 922 370 924 372
rect 927 370 929 372
rect 932 370 934 372
rect 937 370 939 372
rect 942 370 944 372
rect 947 370 949 372
rect 952 370 954 372
rect 957 370 959 372
rect 962 370 964 372
rect 967 370 969 372
rect 972 370 974 372
rect 977 370 979 372
rect 982 370 984 372
rect 987 370 989 372
rect 992 370 994 372
rect 997 370 999 372
rect 577 365 579 367
rect 582 365 584 367
rect 587 365 589 367
rect 592 365 594 367
rect 597 365 599 367
rect 602 365 604 367
rect 607 365 609 367
rect 612 365 614 367
rect 617 365 619 367
rect 622 365 624 367
rect 627 365 629 367
rect 632 365 634 367
rect 637 365 639 367
rect 642 365 644 367
rect 647 365 649 367
rect 652 365 654 367
rect 657 365 659 367
rect 662 365 664 367
rect 667 365 669 367
rect 672 365 674 367
rect 677 365 679 367
rect 682 365 684 367
rect 687 365 689 367
rect 692 365 694 367
rect 697 365 699 367
rect 702 365 704 367
rect 707 365 709 367
rect 712 365 714 367
rect 717 365 719 367
rect 722 365 724 367
rect 727 365 729 367
rect 732 365 734 367
rect 737 365 739 367
rect 742 365 744 367
rect 747 365 749 367
rect 752 365 754 367
rect 757 365 759 367
rect 762 365 764 367
rect 767 365 769 367
rect 772 365 774 367
rect 777 365 779 367
rect 782 365 784 367
rect 787 365 789 367
rect 792 365 794 367
rect 797 365 799 367
rect 802 365 804 367
rect 807 365 809 367
rect 812 365 814 367
rect 817 365 819 367
rect 822 365 824 367
rect 827 365 829 367
rect 832 365 834 367
rect 837 365 839 367
rect 842 365 844 367
rect 847 365 849 367
rect 852 365 854 367
rect 857 365 859 367
rect 862 365 864 367
rect 867 365 869 367
rect 872 365 874 367
rect 877 365 879 367
rect 882 365 884 367
rect 887 365 889 367
rect 892 365 894 367
rect 897 365 899 367
rect 902 365 904 367
rect 907 365 909 367
rect 912 365 914 367
rect 917 365 919 367
rect 922 365 924 367
rect 927 365 929 367
rect 932 365 934 367
rect 937 365 939 367
rect 942 365 944 367
rect 947 365 949 367
rect 952 365 954 367
rect 957 365 959 367
rect 962 365 964 367
rect 967 365 969 367
rect 972 365 974 367
rect 977 365 979 367
rect 982 365 984 367
rect 987 365 989 367
rect 992 365 994 367
rect 997 365 999 367
rect 577 360 579 362
rect 582 360 584 362
rect 587 360 589 362
rect 592 360 594 362
rect 597 360 599 362
rect 602 360 604 362
rect 607 360 609 362
rect 612 360 614 362
rect 617 360 619 362
rect 622 360 624 362
rect 627 360 629 362
rect 632 360 634 362
rect 637 360 639 362
rect 642 360 644 362
rect 647 360 649 362
rect 652 360 654 362
rect 657 360 659 362
rect 662 360 664 362
rect 667 360 669 362
rect 672 360 674 362
rect 677 360 679 362
rect 682 360 684 362
rect 687 360 689 362
rect 692 360 694 362
rect 697 360 699 362
rect 702 360 704 362
rect 707 360 709 362
rect 712 360 714 362
rect 717 360 719 362
rect 722 360 724 362
rect 727 360 729 362
rect 732 360 734 362
rect 737 360 739 362
rect 742 360 744 362
rect 747 360 749 362
rect 752 360 754 362
rect 757 360 759 362
rect 762 360 764 362
rect 767 360 769 362
rect 772 360 774 362
rect 777 360 779 362
rect 782 360 784 362
rect 787 360 789 362
rect 792 360 794 362
rect 797 360 799 362
rect 802 360 804 362
rect 807 360 809 362
rect 812 360 814 362
rect 817 360 819 362
rect 822 360 824 362
rect 827 360 829 362
rect 832 360 834 362
rect 837 360 839 362
rect 842 360 844 362
rect 847 360 849 362
rect 852 360 854 362
rect 857 360 859 362
rect 862 360 864 362
rect 867 360 869 362
rect 872 360 874 362
rect 877 360 879 362
rect 882 360 884 362
rect 887 360 889 362
rect 892 360 894 362
rect 897 360 899 362
rect 902 360 904 362
rect 907 360 909 362
rect 912 360 914 362
rect 917 360 919 362
rect 922 360 924 362
rect 927 360 929 362
rect 932 360 934 362
rect 937 360 939 362
rect 942 360 944 362
rect 947 360 949 362
rect 952 360 954 362
rect 957 360 959 362
rect 962 360 964 362
rect 967 360 969 362
rect 972 360 974 362
rect 977 360 979 362
rect 982 360 984 362
rect 987 360 989 362
rect 992 360 994 362
rect 997 360 999 362
rect 577 355 579 357
rect 582 355 584 357
rect 587 355 589 357
rect 592 355 594 357
rect 597 355 599 357
rect 602 355 604 357
rect 607 355 609 357
rect 612 355 614 357
rect 617 355 619 357
rect 622 355 624 357
rect 627 355 629 357
rect 632 355 634 357
rect 637 355 639 357
rect 642 355 644 357
rect 647 355 649 357
rect 652 355 654 357
rect 657 355 659 357
rect 662 355 664 357
rect 667 355 669 357
rect 672 355 674 357
rect 677 355 679 357
rect 682 355 684 357
rect 687 355 689 357
rect 692 355 694 357
rect 697 355 699 357
rect 702 355 704 357
rect 707 355 709 357
rect 712 355 714 357
rect 717 355 719 357
rect 722 355 724 357
rect 727 355 729 357
rect 732 355 734 357
rect 737 355 739 357
rect 742 355 744 357
rect 747 355 749 357
rect 752 355 754 357
rect 757 355 759 357
rect 762 355 764 357
rect 767 355 769 357
rect 772 355 774 357
rect 777 355 779 357
rect 782 355 784 357
rect 787 355 789 357
rect 792 355 794 357
rect 797 355 799 357
rect 802 355 804 357
rect 807 355 809 357
rect 812 355 814 357
rect 817 355 819 357
rect 822 355 824 357
rect 827 355 829 357
rect 832 355 834 357
rect 837 355 839 357
rect 842 355 844 357
rect 847 355 849 357
rect 852 355 854 357
rect 857 355 859 357
rect 862 355 864 357
rect 867 355 869 357
rect 872 355 874 357
rect 877 355 879 357
rect 882 355 884 357
rect 887 355 889 357
rect 892 355 894 357
rect 897 355 899 357
rect 902 355 904 357
rect 907 355 909 357
rect 912 355 914 357
rect 917 355 919 357
rect 922 355 924 357
rect 927 355 929 357
rect 932 355 934 357
rect 937 355 939 357
rect 942 355 944 357
rect 947 355 949 357
rect 952 355 954 357
rect 957 355 959 357
rect 962 355 964 357
rect 967 355 969 357
rect 972 355 974 357
rect 977 355 979 357
rect 982 355 984 357
rect 987 355 989 357
rect 992 355 994 357
rect 997 355 999 357
rect 577 350 579 352
rect 582 350 584 352
rect 587 350 589 352
rect 592 350 594 352
rect 597 350 599 352
rect 602 350 604 352
rect 607 350 609 352
rect 612 350 614 352
rect 617 350 619 352
rect 622 350 624 352
rect 627 350 629 352
rect 632 350 634 352
rect 637 350 639 352
rect 642 350 644 352
rect 647 350 649 352
rect 652 350 654 352
rect 657 350 659 352
rect 662 350 664 352
rect 667 350 669 352
rect 672 350 674 352
rect 677 350 679 352
rect 682 350 684 352
rect 687 350 689 352
rect 692 350 694 352
rect 697 350 699 352
rect 702 350 704 352
rect 707 350 709 352
rect 712 350 714 352
rect 717 350 719 352
rect 722 350 724 352
rect 727 350 729 352
rect 732 350 734 352
rect 737 350 739 352
rect 742 350 744 352
rect 747 350 749 352
rect 752 350 754 352
rect 757 350 759 352
rect 762 350 764 352
rect 767 350 769 352
rect 772 350 774 352
rect 777 350 779 352
rect 782 350 784 352
rect 787 350 789 352
rect 792 350 794 352
rect 797 350 799 352
rect 802 350 804 352
rect 807 350 809 352
rect 812 350 814 352
rect 817 350 819 352
rect 822 350 824 352
rect 827 350 829 352
rect 832 350 834 352
rect 837 350 839 352
rect 842 350 844 352
rect 847 350 849 352
rect 852 350 854 352
rect 857 350 859 352
rect 862 350 864 352
rect 867 350 869 352
rect 872 350 874 352
rect 877 350 879 352
rect 882 350 884 352
rect 887 350 889 352
rect 892 350 894 352
rect 897 350 899 352
rect 902 350 904 352
rect 907 350 909 352
rect 912 350 914 352
rect 917 350 919 352
rect 922 350 924 352
rect 927 350 929 352
rect 932 350 934 352
rect 937 350 939 352
rect 942 350 944 352
rect 947 350 949 352
rect 952 350 954 352
rect 957 350 959 352
rect 962 350 964 352
rect 967 350 969 352
rect 972 350 974 352
rect 977 350 979 352
rect 982 350 984 352
rect 987 350 989 352
rect 992 350 994 352
rect 997 350 999 352
rect 577 345 579 347
rect 582 345 584 347
rect 587 345 589 347
rect 592 345 594 347
rect 597 345 599 347
rect 602 345 604 347
rect 607 345 609 347
rect 612 345 614 347
rect 617 345 619 347
rect 622 345 624 347
rect 627 345 629 347
rect 632 345 634 347
rect 637 345 639 347
rect 642 345 644 347
rect 647 345 649 347
rect 652 345 654 347
rect 657 345 659 347
rect 662 345 664 347
rect 667 345 669 347
rect 672 345 674 347
rect 677 345 679 347
rect 682 345 684 347
rect 687 345 689 347
rect 692 345 694 347
rect 697 345 699 347
rect 702 345 704 347
rect 707 345 709 347
rect 712 345 714 347
rect 717 345 719 347
rect 722 345 724 347
rect 727 345 729 347
rect 732 345 734 347
rect 737 345 739 347
rect 742 345 744 347
rect 747 345 749 347
rect 752 345 754 347
rect 757 345 759 347
rect 762 345 764 347
rect 767 345 769 347
rect 772 345 774 347
rect 777 345 779 347
rect 782 345 784 347
rect 787 345 789 347
rect 792 345 794 347
rect 797 345 799 347
rect 802 345 804 347
rect 807 345 809 347
rect 812 345 814 347
rect 817 345 819 347
rect 822 345 824 347
rect 827 345 829 347
rect 832 345 834 347
rect 837 345 839 347
rect 842 345 844 347
rect 847 345 849 347
rect 852 345 854 347
rect 857 345 859 347
rect 862 345 864 347
rect 867 345 869 347
rect 872 345 874 347
rect 877 345 879 347
rect 882 345 884 347
rect 887 345 889 347
rect 892 345 894 347
rect 897 345 899 347
rect 902 345 904 347
rect 907 345 909 347
rect 912 345 914 347
rect 917 345 919 347
rect 922 345 924 347
rect 927 345 929 347
rect 932 345 934 347
rect 937 345 939 347
rect 942 345 944 347
rect 947 345 949 347
rect 952 345 954 347
rect 957 345 959 347
rect 962 345 964 347
rect 967 345 969 347
rect 972 345 974 347
rect 977 345 979 347
rect 982 345 984 347
rect 987 345 989 347
rect 992 345 994 347
rect 997 345 999 347
rect 577 339 579 341
rect 582 339 584 341
rect 587 339 589 341
rect 592 339 594 341
rect 597 339 599 341
rect 602 339 604 341
rect 607 339 609 341
rect 612 339 614 341
rect 617 339 619 341
rect 622 339 624 341
rect 627 339 629 341
rect 632 339 634 341
rect 637 339 639 341
rect 642 339 644 341
rect 647 339 649 341
rect 652 339 654 341
rect 577 334 579 336
rect 582 334 584 336
rect 587 334 589 336
rect 592 334 594 336
rect 597 334 599 336
rect 602 334 604 336
rect 607 334 609 336
rect 612 334 614 336
rect 617 334 619 336
rect 622 334 624 336
rect 627 334 629 336
rect 632 334 634 336
rect 637 334 639 336
rect 642 334 644 336
rect 647 334 649 336
rect 652 334 654 336
rect 577 329 579 331
rect 582 329 584 331
rect 587 329 589 331
rect 592 329 594 331
rect 597 329 599 331
rect 602 329 604 331
rect 607 329 609 331
rect 612 329 614 331
rect 617 329 619 331
rect 622 329 624 331
rect 627 329 629 331
rect 632 329 634 331
rect 637 329 639 331
rect 642 329 644 331
rect 647 329 649 331
rect 652 329 654 331
rect 577 324 579 326
rect 582 324 584 326
rect 587 324 589 326
rect 592 324 594 326
rect 597 324 599 326
rect 602 324 604 326
rect 607 324 609 326
rect 612 324 614 326
rect 617 324 619 326
rect 622 324 624 326
rect 627 324 629 326
rect 632 324 634 326
rect 637 324 639 326
rect 642 324 644 326
rect 647 324 649 326
rect 652 324 654 326
rect 676 323 678 325
rect 681 323 683 325
rect 686 323 688 325
rect 691 323 693 325
rect 696 323 698 325
rect 701 323 703 325
rect 706 323 708 325
rect 711 323 713 325
rect 716 323 718 325
rect 721 323 723 325
rect 726 323 728 325
rect 731 323 733 325
rect 736 323 738 325
rect 741 323 743 325
rect 746 323 748 325
rect 751 323 753 325
rect 756 323 758 325
rect 761 323 763 325
rect 766 323 768 325
rect 771 323 773 325
rect 776 323 778 325
rect 781 323 783 325
rect 786 323 788 325
rect 791 323 793 325
rect 796 323 798 325
rect 801 323 803 325
rect 806 323 808 325
rect 811 323 813 325
rect 816 323 818 325
rect 821 323 823 325
rect 826 323 828 325
rect 831 323 833 325
rect 836 323 838 325
rect 841 323 843 325
rect 846 323 848 325
rect 851 323 853 325
rect 856 323 858 325
rect 861 323 863 325
rect 866 323 868 325
rect 871 323 873 325
rect 876 323 878 325
rect 881 323 883 325
rect 886 323 888 325
rect 891 323 893 325
rect 896 323 898 325
rect 901 323 903 325
rect 906 323 908 325
rect 911 323 913 325
rect 916 323 918 325
rect 921 323 923 325
rect 926 323 928 325
rect 931 323 933 325
rect 936 323 938 325
rect 941 323 943 325
rect 946 323 948 325
rect 951 323 953 325
rect 956 323 958 325
rect 961 323 963 325
rect 966 323 968 325
rect 971 323 973 325
rect 976 323 978 325
rect 981 323 983 325
rect 986 323 988 325
rect 991 323 993 325
rect 996 323 998 325
rect 577 319 579 321
rect 582 319 584 321
rect 587 319 589 321
rect 592 319 594 321
rect 597 319 599 321
rect 602 319 604 321
rect 607 319 609 321
rect 612 319 614 321
rect 617 319 619 321
rect 622 319 624 321
rect 627 319 629 321
rect 632 319 634 321
rect 637 319 639 321
rect 642 319 644 321
rect 647 319 649 321
rect 652 319 654 321
rect 676 318 678 320
rect 681 318 683 320
rect 686 318 688 320
rect 691 318 693 320
rect 696 318 698 320
rect 701 318 703 320
rect 706 318 708 320
rect 711 318 713 320
rect 716 318 718 320
rect 721 318 723 320
rect 726 318 728 320
rect 731 318 733 320
rect 736 318 738 320
rect 741 318 743 320
rect 746 318 748 320
rect 751 318 753 320
rect 756 318 758 320
rect 761 318 763 320
rect 766 318 768 320
rect 771 318 773 320
rect 776 318 778 320
rect 781 318 783 320
rect 786 318 788 320
rect 791 318 793 320
rect 796 318 798 320
rect 801 318 803 320
rect 806 318 808 320
rect 811 318 813 320
rect 816 318 818 320
rect 821 318 823 320
rect 826 318 828 320
rect 831 318 833 320
rect 836 318 838 320
rect 841 318 843 320
rect 846 318 848 320
rect 851 318 853 320
rect 856 318 858 320
rect 861 318 863 320
rect 866 318 868 320
rect 871 318 873 320
rect 876 318 878 320
rect 881 318 883 320
rect 886 318 888 320
rect 891 318 893 320
rect 896 318 898 320
rect 901 318 903 320
rect 906 318 908 320
rect 911 318 913 320
rect 916 318 918 320
rect 921 318 923 320
rect 926 318 928 320
rect 931 318 933 320
rect 936 318 938 320
rect 941 318 943 320
rect 946 318 948 320
rect 951 318 953 320
rect 956 318 958 320
rect 961 318 963 320
rect 966 318 968 320
rect 971 318 973 320
rect 976 318 978 320
rect 981 318 983 320
rect 986 318 988 320
rect 991 318 993 320
rect 996 318 998 320
rect 577 314 579 316
rect 582 314 584 316
rect 587 314 589 316
rect 592 314 594 316
rect 597 314 599 316
rect 602 314 604 316
rect 607 314 609 316
rect 612 314 614 316
rect 617 314 619 316
rect 622 314 624 316
rect 627 314 629 316
rect 632 314 634 316
rect 637 314 639 316
rect 642 314 644 316
rect 647 314 649 316
rect 652 314 654 316
rect 676 313 678 315
rect 681 313 683 315
rect 686 313 688 315
rect 691 313 693 315
rect 696 313 698 315
rect 701 313 703 315
rect 706 313 708 315
rect 711 313 713 315
rect 716 313 718 315
rect 721 313 723 315
rect 726 313 728 315
rect 731 313 733 315
rect 736 313 738 315
rect 741 313 743 315
rect 746 313 748 315
rect 751 313 753 315
rect 756 313 758 315
rect 761 313 763 315
rect 766 313 768 315
rect 771 313 773 315
rect 776 313 778 315
rect 781 313 783 315
rect 786 313 788 315
rect 791 313 793 315
rect 796 313 798 315
rect 801 313 803 315
rect 806 313 808 315
rect 811 313 813 315
rect 816 313 818 315
rect 821 313 823 315
rect 826 313 828 315
rect 831 313 833 315
rect 836 313 838 315
rect 841 313 843 315
rect 846 313 848 315
rect 851 313 853 315
rect 856 313 858 315
rect 861 313 863 315
rect 866 313 868 315
rect 871 313 873 315
rect 876 313 878 315
rect 881 313 883 315
rect 886 313 888 315
rect 891 313 893 315
rect 896 313 898 315
rect 901 313 903 315
rect 906 313 908 315
rect 911 313 913 315
rect 916 313 918 315
rect 921 313 923 315
rect 926 313 928 315
rect 931 313 933 315
rect 936 313 938 315
rect 941 313 943 315
rect 946 313 948 315
rect 951 313 953 315
rect 956 313 958 315
rect 961 313 963 315
rect 966 313 968 315
rect 971 313 973 315
rect 976 313 978 315
rect 981 313 983 315
rect 986 313 988 315
rect 991 313 993 315
rect 996 313 998 315
rect 577 309 579 311
rect 582 309 584 311
rect 587 309 589 311
rect 592 309 594 311
rect 597 309 599 311
rect 602 309 604 311
rect 607 309 609 311
rect 612 309 614 311
rect 617 309 619 311
rect 622 309 624 311
rect 627 309 629 311
rect 632 309 634 311
rect 637 309 639 311
rect 642 309 644 311
rect 647 309 649 311
rect 652 309 654 311
rect 676 308 678 310
rect 681 308 683 310
rect 686 308 688 310
rect 691 308 693 310
rect 696 308 698 310
rect 701 308 703 310
rect 706 308 708 310
rect 711 308 713 310
rect 716 308 718 310
rect 721 308 723 310
rect 726 308 728 310
rect 731 308 733 310
rect 736 308 738 310
rect 741 308 743 310
rect 746 308 748 310
rect 751 308 753 310
rect 756 308 758 310
rect 761 308 763 310
rect 766 308 768 310
rect 771 308 773 310
rect 776 308 778 310
rect 781 308 783 310
rect 786 308 788 310
rect 791 308 793 310
rect 796 308 798 310
rect 801 308 803 310
rect 806 308 808 310
rect 811 308 813 310
rect 816 308 818 310
rect 821 308 823 310
rect 826 308 828 310
rect 831 308 833 310
rect 836 308 838 310
rect 841 308 843 310
rect 846 308 848 310
rect 851 308 853 310
rect 856 308 858 310
rect 861 308 863 310
rect 866 308 868 310
rect 871 308 873 310
rect 876 308 878 310
rect 881 308 883 310
rect 886 308 888 310
rect 891 308 893 310
rect 896 308 898 310
rect 901 308 903 310
rect 906 308 908 310
rect 911 308 913 310
rect 916 308 918 310
rect 921 308 923 310
rect 926 308 928 310
rect 931 308 933 310
rect 936 308 938 310
rect 941 308 943 310
rect 946 308 948 310
rect 951 308 953 310
rect 956 308 958 310
rect 961 308 963 310
rect 966 308 968 310
rect 971 308 973 310
rect 976 308 978 310
rect 981 308 983 310
rect 986 308 988 310
rect 991 308 993 310
rect 996 308 998 310
rect 577 304 579 306
rect 582 304 584 306
rect 587 304 589 306
rect 592 304 594 306
rect 597 304 599 306
rect 602 304 604 306
rect 607 304 609 306
rect 612 304 614 306
rect 617 304 619 306
rect 622 304 624 306
rect 627 304 629 306
rect 632 304 634 306
rect 637 304 639 306
rect 642 304 644 306
rect 647 304 649 306
rect 652 304 654 306
rect 676 303 678 305
rect 681 303 683 305
rect 686 303 688 305
rect 691 303 693 305
rect 696 303 698 305
rect 701 303 703 305
rect 706 303 708 305
rect 711 303 713 305
rect 716 303 718 305
rect 721 303 723 305
rect 726 303 728 305
rect 731 303 733 305
rect 736 303 738 305
rect 741 303 743 305
rect 746 303 748 305
rect 751 303 753 305
rect 756 303 758 305
rect 761 303 763 305
rect 766 303 768 305
rect 771 303 773 305
rect 776 303 778 305
rect 781 303 783 305
rect 786 303 788 305
rect 791 303 793 305
rect 796 303 798 305
rect 801 303 803 305
rect 806 303 808 305
rect 811 303 813 305
rect 816 303 818 305
rect 821 303 823 305
rect 826 303 828 305
rect 831 303 833 305
rect 836 303 838 305
rect 841 303 843 305
rect 846 303 848 305
rect 851 303 853 305
rect 856 303 858 305
rect 861 303 863 305
rect 866 303 868 305
rect 871 303 873 305
rect 876 303 878 305
rect 881 303 883 305
rect 886 303 888 305
rect 891 303 893 305
rect 896 303 898 305
rect 901 303 903 305
rect 906 303 908 305
rect 911 303 913 305
rect 916 303 918 305
rect 921 303 923 305
rect 926 303 928 305
rect 931 303 933 305
rect 936 303 938 305
rect 941 303 943 305
rect 946 303 948 305
rect 951 303 953 305
rect 956 303 958 305
rect 961 303 963 305
rect 966 303 968 305
rect 971 303 973 305
rect 976 303 978 305
rect 981 303 983 305
rect 986 303 988 305
rect 991 303 993 305
rect 996 303 998 305
rect 577 299 579 301
rect 582 299 584 301
rect 587 299 589 301
rect 592 299 594 301
rect 597 299 599 301
rect 602 299 604 301
rect 607 299 609 301
rect 612 299 614 301
rect 617 299 619 301
rect 622 299 624 301
rect 627 299 629 301
rect 632 299 634 301
rect 637 299 639 301
rect 642 299 644 301
rect 647 299 649 301
rect 652 299 654 301
rect 676 298 678 300
rect 681 298 683 300
rect 686 298 688 300
rect 691 298 693 300
rect 696 298 698 300
rect 701 298 703 300
rect 706 298 708 300
rect 711 298 713 300
rect 716 298 718 300
rect 721 298 723 300
rect 726 298 728 300
rect 731 298 733 300
rect 736 298 738 300
rect 741 298 743 300
rect 746 298 748 300
rect 751 298 753 300
rect 756 298 758 300
rect 761 298 763 300
rect 766 298 768 300
rect 771 298 773 300
rect 776 298 778 300
rect 781 298 783 300
rect 786 298 788 300
rect 791 298 793 300
rect 796 298 798 300
rect 801 298 803 300
rect 806 298 808 300
rect 811 298 813 300
rect 816 298 818 300
rect 821 298 823 300
rect 826 298 828 300
rect 831 298 833 300
rect 836 298 838 300
rect 841 298 843 300
rect 846 298 848 300
rect 851 298 853 300
rect 856 298 858 300
rect 861 298 863 300
rect 866 298 868 300
rect 871 298 873 300
rect 876 298 878 300
rect 881 298 883 300
rect 886 298 888 300
rect 891 298 893 300
rect 896 298 898 300
rect 901 298 903 300
rect 906 298 908 300
rect 911 298 913 300
rect 916 298 918 300
rect 921 298 923 300
rect 926 298 928 300
rect 931 298 933 300
rect 936 298 938 300
rect 941 298 943 300
rect 946 298 948 300
rect 951 298 953 300
rect 956 298 958 300
rect 961 298 963 300
rect 966 298 968 300
rect 971 298 973 300
rect 976 298 978 300
rect 981 298 983 300
rect 986 298 988 300
rect 991 298 993 300
rect 996 298 998 300
rect 577 294 579 296
rect 582 294 584 296
rect 587 294 589 296
rect 592 294 594 296
rect 597 294 599 296
rect 602 294 604 296
rect 607 294 609 296
rect 612 294 614 296
rect 617 294 619 296
rect 622 294 624 296
rect 627 294 629 296
rect 632 294 634 296
rect 637 294 639 296
rect 642 294 644 296
rect 647 294 649 296
rect 652 294 654 296
rect 676 293 678 295
rect 681 293 683 295
rect 686 293 688 295
rect 691 293 693 295
rect 696 293 698 295
rect 701 293 703 295
rect 706 293 708 295
rect 711 293 713 295
rect 716 293 718 295
rect 721 293 723 295
rect 726 293 728 295
rect 731 293 733 295
rect 736 293 738 295
rect 741 293 743 295
rect 746 293 748 295
rect 751 293 753 295
rect 756 293 758 295
rect 761 293 763 295
rect 766 293 768 295
rect 771 293 773 295
rect 776 293 778 295
rect 781 293 783 295
rect 786 293 788 295
rect 791 293 793 295
rect 796 293 798 295
rect 801 293 803 295
rect 806 293 808 295
rect 811 293 813 295
rect 816 293 818 295
rect 821 293 823 295
rect 826 293 828 295
rect 831 293 833 295
rect 836 293 838 295
rect 841 293 843 295
rect 846 293 848 295
rect 851 293 853 295
rect 856 293 858 295
rect 861 293 863 295
rect 866 293 868 295
rect 871 293 873 295
rect 876 293 878 295
rect 881 293 883 295
rect 886 293 888 295
rect 891 293 893 295
rect 896 293 898 295
rect 901 293 903 295
rect 906 293 908 295
rect 911 293 913 295
rect 916 293 918 295
rect 921 293 923 295
rect 926 293 928 295
rect 931 293 933 295
rect 936 293 938 295
rect 941 293 943 295
rect 946 293 948 295
rect 951 293 953 295
rect 956 293 958 295
rect 961 293 963 295
rect 966 293 968 295
rect 971 293 973 295
rect 976 293 978 295
rect 981 293 983 295
rect 986 293 988 295
rect 991 293 993 295
rect 996 293 998 295
rect 577 289 579 291
rect 582 289 584 291
rect 587 289 589 291
rect 592 289 594 291
rect 597 289 599 291
rect 602 289 604 291
rect 607 289 609 291
rect 612 289 614 291
rect 617 289 619 291
rect 622 289 624 291
rect 627 289 629 291
rect 632 289 634 291
rect 637 289 639 291
rect 642 289 644 291
rect 647 289 649 291
rect 652 289 654 291
rect 676 288 678 290
rect 681 288 683 290
rect 686 288 688 290
rect 691 288 693 290
rect 696 288 698 290
rect 701 288 703 290
rect 706 288 708 290
rect 711 288 713 290
rect 716 288 718 290
rect 721 288 723 290
rect 726 288 728 290
rect 731 288 733 290
rect 736 288 738 290
rect 741 288 743 290
rect 746 288 748 290
rect 751 288 753 290
rect 756 288 758 290
rect 761 288 763 290
rect 766 288 768 290
rect 771 288 773 290
rect 776 288 778 290
rect 781 288 783 290
rect 786 288 788 290
rect 791 288 793 290
rect 796 288 798 290
rect 801 288 803 290
rect 806 288 808 290
rect 811 288 813 290
rect 816 288 818 290
rect 821 288 823 290
rect 826 288 828 290
rect 831 288 833 290
rect 836 288 838 290
rect 841 288 843 290
rect 846 288 848 290
rect 851 288 853 290
rect 856 288 858 290
rect 861 288 863 290
rect 866 288 868 290
rect 871 288 873 290
rect 876 288 878 290
rect 881 288 883 290
rect 886 288 888 290
rect 891 288 893 290
rect 896 288 898 290
rect 901 288 903 290
rect 906 288 908 290
rect 911 288 913 290
rect 916 288 918 290
rect 921 288 923 290
rect 926 288 928 290
rect 931 288 933 290
rect 936 288 938 290
rect 941 288 943 290
rect 946 288 948 290
rect 951 288 953 290
rect 956 288 958 290
rect 961 288 963 290
rect 966 288 968 290
rect 971 288 973 290
rect 976 288 978 290
rect 981 288 983 290
rect 986 288 988 290
rect 991 288 993 290
rect 996 288 998 290
rect 577 284 579 286
rect 582 284 584 286
rect 587 284 589 286
rect 592 284 594 286
rect 597 284 599 286
rect 602 284 604 286
rect 607 284 609 286
rect 612 284 614 286
rect 617 284 619 286
rect 622 284 624 286
rect 627 284 629 286
rect 632 284 634 286
rect 637 284 639 286
rect 642 284 644 286
rect 647 284 649 286
rect 652 284 654 286
rect 676 283 678 285
rect 681 283 683 285
rect 686 283 688 285
rect 691 283 693 285
rect 696 283 698 285
rect 701 283 703 285
rect 706 283 708 285
rect 711 283 713 285
rect 716 283 718 285
rect 721 283 723 285
rect 726 283 728 285
rect 731 283 733 285
rect 736 283 738 285
rect 741 283 743 285
rect 746 283 748 285
rect 751 283 753 285
rect 756 283 758 285
rect 761 283 763 285
rect 766 283 768 285
rect 771 283 773 285
rect 776 283 778 285
rect 781 283 783 285
rect 786 283 788 285
rect 791 283 793 285
rect 796 283 798 285
rect 801 283 803 285
rect 806 283 808 285
rect 811 283 813 285
rect 816 283 818 285
rect 821 283 823 285
rect 826 283 828 285
rect 831 283 833 285
rect 836 283 838 285
rect 841 283 843 285
rect 846 283 848 285
rect 851 283 853 285
rect 856 283 858 285
rect 861 283 863 285
rect 866 283 868 285
rect 871 283 873 285
rect 876 283 878 285
rect 881 283 883 285
rect 886 283 888 285
rect 891 283 893 285
rect 896 283 898 285
rect 901 283 903 285
rect 906 283 908 285
rect 911 283 913 285
rect 916 283 918 285
rect 921 283 923 285
rect 926 283 928 285
rect 931 283 933 285
rect 936 283 938 285
rect 941 283 943 285
rect 946 283 948 285
rect 951 283 953 285
rect 956 283 958 285
rect 961 283 963 285
rect 966 283 968 285
rect 971 283 973 285
rect 976 283 978 285
rect 981 283 983 285
rect 986 283 988 285
rect 991 283 993 285
rect 996 283 998 285
rect 577 279 579 281
rect 582 279 584 281
rect 587 279 589 281
rect 592 279 594 281
rect 597 279 599 281
rect 602 279 604 281
rect 607 279 609 281
rect 612 279 614 281
rect 617 279 619 281
rect 622 279 624 281
rect 627 279 629 281
rect 632 279 634 281
rect 637 279 639 281
rect 642 279 644 281
rect 647 279 649 281
rect 652 279 654 281
rect 676 278 678 280
rect 681 278 683 280
rect 686 278 688 280
rect 691 278 693 280
rect 696 278 698 280
rect 701 278 703 280
rect 706 278 708 280
rect 711 278 713 280
rect 716 278 718 280
rect 721 278 723 280
rect 726 278 728 280
rect 731 278 733 280
rect 736 278 738 280
rect 741 278 743 280
rect 746 278 748 280
rect 751 278 753 280
rect 756 278 758 280
rect 761 278 763 280
rect 766 278 768 280
rect 771 278 773 280
rect 776 278 778 280
rect 781 278 783 280
rect 786 278 788 280
rect 791 278 793 280
rect 796 278 798 280
rect 801 278 803 280
rect 806 278 808 280
rect 811 278 813 280
rect 816 278 818 280
rect 821 278 823 280
rect 826 278 828 280
rect 831 278 833 280
rect 836 278 838 280
rect 841 278 843 280
rect 846 278 848 280
rect 851 278 853 280
rect 856 278 858 280
rect 861 278 863 280
rect 866 278 868 280
rect 871 278 873 280
rect 876 278 878 280
rect 881 278 883 280
rect 886 278 888 280
rect 891 278 893 280
rect 896 278 898 280
rect 901 278 903 280
rect 906 278 908 280
rect 911 278 913 280
rect 916 278 918 280
rect 921 278 923 280
rect 926 278 928 280
rect 931 278 933 280
rect 936 278 938 280
rect 941 278 943 280
rect 946 278 948 280
rect 951 278 953 280
rect 956 278 958 280
rect 961 278 963 280
rect 966 278 968 280
rect 971 278 973 280
rect 976 278 978 280
rect 981 278 983 280
rect 986 278 988 280
rect 991 278 993 280
rect 996 278 998 280
rect 577 274 579 276
rect 582 274 584 276
rect 587 274 589 276
rect 592 274 594 276
rect 597 274 599 276
rect 602 274 604 276
rect 607 274 609 276
rect 612 274 614 276
rect 617 274 619 276
rect 622 274 624 276
rect 627 274 629 276
rect 632 274 634 276
rect 637 274 639 276
rect 642 274 644 276
rect 647 274 649 276
rect 652 274 654 276
rect 676 273 678 275
rect 681 273 683 275
rect 686 273 688 275
rect 691 273 693 275
rect 696 273 698 275
rect 701 273 703 275
rect 706 273 708 275
rect 711 273 713 275
rect 716 273 718 275
rect 721 273 723 275
rect 726 273 728 275
rect 731 273 733 275
rect 736 273 738 275
rect 741 273 743 275
rect 746 273 748 275
rect 751 273 753 275
rect 756 273 758 275
rect 761 273 763 275
rect 766 273 768 275
rect 771 273 773 275
rect 776 273 778 275
rect 781 273 783 275
rect 786 273 788 275
rect 791 273 793 275
rect 796 273 798 275
rect 801 273 803 275
rect 806 273 808 275
rect 811 273 813 275
rect 816 273 818 275
rect 821 273 823 275
rect 826 273 828 275
rect 831 273 833 275
rect 836 273 838 275
rect 841 273 843 275
rect 846 273 848 275
rect 851 273 853 275
rect 856 273 858 275
rect 861 273 863 275
rect 866 273 868 275
rect 871 273 873 275
rect 876 273 878 275
rect 881 273 883 275
rect 886 273 888 275
rect 891 273 893 275
rect 896 273 898 275
rect 901 273 903 275
rect 906 273 908 275
rect 911 273 913 275
rect 916 273 918 275
rect 921 273 923 275
rect 926 273 928 275
rect 931 273 933 275
rect 936 273 938 275
rect 941 273 943 275
rect 946 273 948 275
rect 951 273 953 275
rect 956 273 958 275
rect 961 273 963 275
rect 966 273 968 275
rect 971 273 973 275
rect 976 273 978 275
rect 981 273 983 275
rect 986 273 988 275
rect 991 273 993 275
rect 996 273 998 275
rect 577 269 579 271
rect 582 269 584 271
rect 587 269 589 271
rect 592 269 594 271
rect 597 269 599 271
rect 602 269 604 271
rect 607 269 609 271
rect 612 269 614 271
rect 617 269 619 271
rect 622 269 624 271
rect 627 269 629 271
rect 632 269 634 271
rect 637 269 639 271
rect 642 269 644 271
rect 647 269 649 271
rect 652 269 654 271
rect 676 268 678 270
rect 681 268 683 270
rect 686 268 688 270
rect 691 268 693 270
rect 696 268 698 270
rect 701 268 703 270
rect 706 268 708 270
rect 711 268 713 270
rect 716 268 718 270
rect 721 268 723 270
rect 726 268 728 270
rect 731 268 733 270
rect 736 268 738 270
rect 741 268 743 270
rect 746 268 748 270
rect 751 268 753 270
rect 756 268 758 270
rect 761 268 763 270
rect 766 268 768 270
rect 771 268 773 270
rect 776 268 778 270
rect 781 268 783 270
rect 786 268 788 270
rect 791 268 793 270
rect 796 268 798 270
rect 801 268 803 270
rect 806 268 808 270
rect 811 268 813 270
rect 816 268 818 270
rect 821 268 823 270
rect 826 268 828 270
rect 831 268 833 270
rect 836 268 838 270
rect 841 268 843 270
rect 846 268 848 270
rect 851 268 853 270
rect 856 268 858 270
rect 861 268 863 270
rect 866 268 868 270
rect 871 268 873 270
rect 876 268 878 270
rect 881 268 883 270
rect 886 268 888 270
rect 891 268 893 270
rect 896 268 898 270
rect 901 268 903 270
rect 906 268 908 270
rect 911 268 913 270
rect 916 268 918 270
rect 921 268 923 270
rect 926 268 928 270
rect 931 268 933 270
rect 936 268 938 270
rect 941 268 943 270
rect 946 268 948 270
rect 951 268 953 270
rect 956 268 958 270
rect 961 268 963 270
rect 966 268 968 270
rect 971 268 973 270
rect 976 268 978 270
rect 981 268 983 270
rect 986 268 988 270
rect 991 268 993 270
rect 996 268 998 270
rect 577 264 579 266
rect 582 264 584 266
rect 587 264 589 266
rect 592 264 594 266
rect 597 264 599 266
rect 602 264 604 266
rect 607 264 609 266
rect 612 264 614 266
rect 617 264 619 266
rect 622 264 624 266
rect 627 264 629 266
rect 632 264 634 266
rect 637 264 639 266
rect 642 264 644 266
rect 647 264 649 266
rect 652 264 654 266
rect 676 263 678 265
rect 681 263 683 265
rect 686 263 688 265
rect 691 263 693 265
rect 696 263 698 265
rect 701 263 703 265
rect 706 263 708 265
rect 711 263 713 265
rect 716 263 718 265
rect 721 263 723 265
rect 726 263 728 265
rect 731 263 733 265
rect 736 263 738 265
rect 741 263 743 265
rect 746 263 748 265
rect 751 263 753 265
rect 756 263 758 265
rect 761 263 763 265
rect 766 263 768 265
rect 771 263 773 265
rect 776 263 778 265
rect 781 263 783 265
rect 786 263 788 265
rect 791 263 793 265
rect 796 263 798 265
rect 801 263 803 265
rect 806 263 808 265
rect 811 263 813 265
rect 816 263 818 265
rect 821 263 823 265
rect 826 263 828 265
rect 831 263 833 265
rect 836 263 838 265
rect 841 263 843 265
rect 846 263 848 265
rect 851 263 853 265
rect 856 263 858 265
rect 861 263 863 265
rect 866 263 868 265
rect 871 263 873 265
rect 876 263 878 265
rect 881 263 883 265
rect 886 263 888 265
rect 891 263 893 265
rect 896 263 898 265
rect 901 263 903 265
rect 906 263 908 265
rect 911 263 913 265
rect 916 263 918 265
rect 921 263 923 265
rect 926 263 928 265
rect 931 263 933 265
rect 936 263 938 265
rect 941 263 943 265
rect 946 263 948 265
rect 951 263 953 265
rect 956 263 958 265
rect 961 263 963 265
rect 966 263 968 265
rect 971 263 973 265
rect 976 263 978 265
rect 981 263 983 265
rect 986 263 988 265
rect 991 263 993 265
rect 996 263 998 265
rect 577 259 579 261
rect 582 259 584 261
rect 587 259 589 261
rect 592 259 594 261
rect 597 259 599 261
rect 602 259 604 261
rect 607 259 609 261
rect 612 259 614 261
rect 617 259 619 261
rect 622 259 624 261
rect 627 259 629 261
rect 632 259 634 261
rect 637 259 639 261
rect 642 259 644 261
rect 647 259 649 261
rect 652 259 654 261
rect 676 258 678 260
rect 681 258 683 260
rect 686 258 688 260
rect 691 258 693 260
rect 696 258 698 260
rect 701 258 703 260
rect 706 258 708 260
rect 711 258 713 260
rect 716 258 718 260
rect 721 258 723 260
rect 726 258 728 260
rect 731 258 733 260
rect 736 258 738 260
rect 741 258 743 260
rect 746 258 748 260
rect 751 258 753 260
rect 756 258 758 260
rect 761 258 763 260
rect 766 258 768 260
rect 771 258 773 260
rect 776 258 778 260
rect 781 258 783 260
rect 786 258 788 260
rect 791 258 793 260
rect 796 258 798 260
rect 801 258 803 260
rect 806 258 808 260
rect 811 258 813 260
rect 816 258 818 260
rect 821 258 823 260
rect 826 258 828 260
rect 831 258 833 260
rect 836 258 838 260
rect 841 258 843 260
rect 846 258 848 260
rect 851 258 853 260
rect 856 258 858 260
rect 861 258 863 260
rect 866 258 868 260
rect 871 258 873 260
rect 876 258 878 260
rect 881 258 883 260
rect 886 258 888 260
rect 891 258 893 260
rect 896 258 898 260
rect 901 258 903 260
rect 906 258 908 260
rect 911 258 913 260
rect 916 258 918 260
rect 921 258 923 260
rect 926 258 928 260
rect 931 258 933 260
rect 936 258 938 260
rect 941 258 943 260
rect 946 258 948 260
rect 951 258 953 260
rect 956 258 958 260
rect 961 258 963 260
rect 966 258 968 260
rect 971 258 973 260
rect 976 258 978 260
rect 981 258 983 260
rect 986 258 988 260
rect 991 258 993 260
rect 996 258 998 260
rect 577 254 579 256
rect 582 254 584 256
rect 587 254 589 256
rect 592 254 594 256
rect 597 254 599 256
rect 602 254 604 256
rect 607 254 609 256
rect 612 254 614 256
rect 617 254 619 256
rect 622 254 624 256
rect 627 254 629 256
rect 632 254 634 256
rect 637 254 639 256
rect 642 254 644 256
rect 647 254 649 256
rect 652 254 654 256
rect 676 253 678 255
rect 681 253 683 255
rect 686 253 688 255
rect 691 253 693 255
rect 696 253 698 255
rect 701 253 703 255
rect 706 253 708 255
rect 711 253 713 255
rect 716 253 718 255
rect 721 253 723 255
rect 726 253 728 255
rect 731 253 733 255
rect 736 253 738 255
rect 741 253 743 255
rect 746 253 748 255
rect 751 253 753 255
rect 756 253 758 255
rect 761 253 763 255
rect 766 253 768 255
rect 771 253 773 255
rect 776 253 778 255
rect 781 253 783 255
rect 786 253 788 255
rect 791 253 793 255
rect 796 253 798 255
rect 801 253 803 255
rect 806 253 808 255
rect 811 253 813 255
rect 816 253 818 255
rect 821 253 823 255
rect 826 253 828 255
rect 831 253 833 255
rect 836 253 838 255
rect 841 253 843 255
rect 846 253 848 255
rect 851 253 853 255
rect 856 253 858 255
rect 861 253 863 255
rect 866 253 868 255
rect 871 253 873 255
rect 876 253 878 255
rect 881 253 883 255
rect 886 253 888 255
rect 891 253 893 255
rect 896 253 898 255
rect 901 253 903 255
rect 906 253 908 255
rect 911 253 913 255
rect 916 253 918 255
rect 921 253 923 255
rect 926 253 928 255
rect 931 253 933 255
rect 936 253 938 255
rect 941 253 943 255
rect 946 253 948 255
rect 951 253 953 255
rect 956 253 958 255
rect 961 253 963 255
rect 966 253 968 255
rect 971 253 973 255
rect 976 253 978 255
rect 981 253 983 255
rect 986 253 988 255
rect 991 253 993 255
rect 996 253 998 255
rect 577 249 579 251
rect 582 249 584 251
rect 587 249 589 251
rect 592 249 594 251
rect 597 249 599 251
rect 602 249 604 251
rect 607 249 609 251
rect 612 249 614 251
rect 617 249 619 251
rect 622 249 624 251
rect 627 249 629 251
rect 632 249 634 251
rect 637 249 639 251
rect 642 249 644 251
rect 647 249 649 251
rect 652 249 654 251
rect 676 248 678 250
rect 681 248 683 250
rect 686 248 688 250
rect 691 248 693 250
rect 696 248 698 250
rect 701 248 703 250
rect 706 248 708 250
rect 711 248 713 250
rect 716 248 718 250
rect 721 248 723 250
rect 726 248 728 250
rect 731 248 733 250
rect 736 248 738 250
rect 741 248 743 250
rect 746 248 748 250
rect 751 248 753 250
rect 756 248 758 250
rect 761 248 763 250
rect 766 248 768 250
rect 771 248 773 250
rect 776 248 778 250
rect 781 248 783 250
rect 786 248 788 250
rect 791 248 793 250
rect 796 248 798 250
rect 801 248 803 250
rect 806 248 808 250
rect 811 248 813 250
rect 816 248 818 250
rect 821 248 823 250
rect 826 248 828 250
rect 831 248 833 250
rect 836 248 838 250
rect 841 248 843 250
rect 846 248 848 250
rect 851 248 853 250
rect 856 248 858 250
rect 861 248 863 250
rect 866 248 868 250
rect 871 248 873 250
rect 876 248 878 250
rect 881 248 883 250
rect 886 248 888 250
rect 891 248 893 250
rect 896 248 898 250
rect 901 248 903 250
rect 906 248 908 250
rect 911 248 913 250
rect 916 248 918 250
rect 921 248 923 250
rect 926 248 928 250
rect 931 248 933 250
rect 936 248 938 250
rect 941 248 943 250
rect 946 248 948 250
rect 951 248 953 250
rect 956 248 958 250
rect 961 248 963 250
rect 966 248 968 250
rect 971 248 973 250
rect 976 248 978 250
rect 981 248 983 250
rect 986 248 988 250
rect 991 248 993 250
rect 996 248 998 250
rect 577 244 579 246
rect 582 244 584 246
rect 587 244 589 246
rect 592 244 594 246
rect 597 244 599 246
rect 602 244 604 246
rect 607 244 609 246
rect 612 244 614 246
rect 617 244 619 246
rect 622 244 624 246
rect 627 244 629 246
rect 632 244 634 246
rect 637 244 639 246
rect 642 244 644 246
rect 647 244 649 246
rect 652 244 654 246
rect 675 241 677 243
rect 680 241 682 243
rect 685 241 687 243
rect 690 241 692 243
rect 695 241 697 243
rect 700 241 702 243
rect 705 241 707 243
rect 710 241 712 243
rect 715 241 717 243
rect 720 241 722 243
rect 725 241 727 243
rect 730 241 732 243
rect 735 241 737 243
rect 740 241 742 243
rect 745 241 747 243
rect 750 241 752 243
rect 577 239 579 241
rect 582 239 584 241
rect 587 239 589 241
rect 592 239 594 241
rect 597 239 599 241
rect 602 239 604 241
rect 607 239 609 241
rect 612 239 614 241
rect 617 239 619 241
rect 622 239 624 241
rect 627 239 629 241
rect 632 239 634 241
rect 637 239 639 241
rect 642 239 644 241
rect 647 239 649 241
rect 652 239 654 241
rect 675 236 677 238
rect 680 236 682 238
rect 685 236 687 238
rect 690 236 692 238
rect 695 236 697 238
rect 700 236 702 238
rect 705 236 707 238
rect 710 236 712 238
rect 715 236 717 238
rect 720 236 722 238
rect 725 236 727 238
rect 730 236 732 238
rect 735 236 737 238
rect 740 236 742 238
rect 745 236 747 238
rect 750 236 752 238
rect 577 234 579 236
rect 582 234 584 236
rect 587 234 589 236
rect 592 234 594 236
rect 597 234 599 236
rect 602 234 604 236
rect 607 234 609 236
rect 612 234 614 236
rect 617 234 619 236
rect 622 234 624 236
rect 627 234 629 236
rect 632 234 634 236
rect 637 234 639 236
rect 642 234 644 236
rect 647 234 649 236
rect 652 234 654 236
rect 675 231 677 233
rect 680 231 682 233
rect 685 231 687 233
rect 690 231 692 233
rect 695 231 697 233
rect 700 231 702 233
rect 705 231 707 233
rect 710 231 712 233
rect 715 231 717 233
rect 720 231 722 233
rect 725 231 727 233
rect 730 231 732 233
rect 735 231 737 233
rect 740 231 742 233
rect 745 231 747 233
rect 750 231 752 233
rect 577 229 579 231
rect 582 229 584 231
rect 587 229 589 231
rect 592 229 594 231
rect 597 229 599 231
rect 602 229 604 231
rect 607 229 609 231
rect 612 229 614 231
rect 617 229 619 231
rect 622 229 624 231
rect 627 229 629 231
rect 632 229 634 231
rect 637 229 639 231
rect 642 229 644 231
rect 647 229 649 231
rect 652 229 654 231
rect 675 226 677 228
rect 680 226 682 228
rect 685 226 687 228
rect 690 226 692 228
rect 695 226 697 228
rect 700 226 702 228
rect 705 226 707 228
rect 710 226 712 228
rect 715 226 717 228
rect 720 226 722 228
rect 725 226 727 228
rect 730 226 732 228
rect 735 226 737 228
rect 740 226 742 228
rect 745 226 747 228
rect 750 226 752 228
rect 577 224 579 226
rect 582 224 584 226
rect 587 224 589 226
rect 592 224 594 226
rect 597 224 599 226
rect 602 224 604 226
rect 607 224 609 226
rect 612 224 614 226
rect 617 224 619 226
rect 622 224 624 226
rect 627 224 629 226
rect 632 224 634 226
rect 637 224 639 226
rect 642 224 644 226
rect 647 224 649 226
rect 652 224 654 226
rect 675 221 677 223
rect 680 221 682 223
rect 685 221 687 223
rect 690 221 692 223
rect 695 221 697 223
rect 700 221 702 223
rect 705 221 707 223
rect 710 221 712 223
rect 715 221 717 223
rect 720 221 722 223
rect 725 221 727 223
rect 730 221 732 223
rect 735 221 737 223
rect 740 221 742 223
rect 745 221 747 223
rect 750 221 752 223
rect 577 219 579 221
rect 582 219 584 221
rect 587 219 589 221
rect 592 219 594 221
rect 597 219 599 221
rect 602 219 604 221
rect 607 219 609 221
rect 612 219 614 221
rect 617 219 619 221
rect 622 219 624 221
rect 627 219 629 221
rect 632 219 634 221
rect 637 219 639 221
rect 642 219 644 221
rect 647 219 649 221
rect 652 219 654 221
rect 675 216 677 218
rect 680 216 682 218
rect 685 216 687 218
rect 690 216 692 218
rect 695 216 697 218
rect 700 216 702 218
rect 705 216 707 218
rect 710 216 712 218
rect 715 216 717 218
rect 720 216 722 218
rect 725 216 727 218
rect 730 216 732 218
rect 735 216 737 218
rect 740 216 742 218
rect 745 216 747 218
rect 750 216 752 218
rect 577 214 579 216
rect 582 214 584 216
rect 587 214 589 216
rect 592 214 594 216
rect 597 214 599 216
rect 602 214 604 216
rect 607 214 609 216
rect 612 214 614 216
rect 617 214 619 216
rect 622 214 624 216
rect 627 214 629 216
rect 632 214 634 216
rect 637 214 639 216
rect 642 214 644 216
rect 647 214 649 216
rect 652 214 654 216
rect 675 211 677 213
rect 680 211 682 213
rect 685 211 687 213
rect 690 211 692 213
rect 695 211 697 213
rect 700 211 702 213
rect 705 211 707 213
rect 710 211 712 213
rect 715 211 717 213
rect 720 211 722 213
rect 725 211 727 213
rect 730 211 732 213
rect 735 211 737 213
rect 740 211 742 213
rect 745 211 747 213
rect 750 211 752 213
rect 577 209 579 211
rect 582 209 584 211
rect 587 209 589 211
rect 592 209 594 211
rect 597 209 599 211
rect 602 209 604 211
rect 607 209 609 211
rect 612 209 614 211
rect 617 209 619 211
rect 622 209 624 211
rect 627 209 629 211
rect 632 209 634 211
rect 637 209 639 211
rect 642 209 644 211
rect 647 209 649 211
rect 652 209 654 211
rect 675 206 677 208
rect 680 206 682 208
rect 685 206 687 208
rect 690 206 692 208
rect 695 206 697 208
rect 700 206 702 208
rect 705 206 707 208
rect 710 206 712 208
rect 715 206 717 208
rect 720 206 722 208
rect 725 206 727 208
rect 730 206 732 208
rect 735 206 737 208
rect 740 206 742 208
rect 745 206 747 208
rect 750 206 752 208
rect 577 204 579 206
rect 582 204 584 206
rect 587 204 589 206
rect 592 204 594 206
rect 597 204 599 206
rect 602 204 604 206
rect 607 204 609 206
rect 612 204 614 206
rect 617 204 619 206
rect 622 204 624 206
rect 627 204 629 206
rect 632 204 634 206
rect 637 204 639 206
rect 642 204 644 206
rect 647 204 649 206
rect 652 204 654 206
rect 675 201 677 203
rect 680 201 682 203
rect 685 201 687 203
rect 690 201 692 203
rect 695 201 697 203
rect 700 201 702 203
rect 705 201 707 203
rect 710 201 712 203
rect 715 201 717 203
rect 720 201 722 203
rect 725 201 727 203
rect 730 201 732 203
rect 735 201 737 203
rect 740 201 742 203
rect 745 201 747 203
rect 750 201 752 203
rect 577 199 579 201
rect 582 199 584 201
rect 587 199 589 201
rect 592 199 594 201
rect 597 199 599 201
rect 602 199 604 201
rect 607 199 609 201
rect 612 199 614 201
rect 617 199 619 201
rect 622 199 624 201
rect 627 199 629 201
rect 632 199 634 201
rect 637 199 639 201
rect 642 199 644 201
rect 647 199 649 201
rect 652 199 654 201
rect 675 196 677 198
rect 680 196 682 198
rect 685 196 687 198
rect 690 196 692 198
rect 695 196 697 198
rect 700 196 702 198
rect 705 196 707 198
rect 710 196 712 198
rect 715 196 717 198
rect 720 196 722 198
rect 725 196 727 198
rect 730 196 732 198
rect 735 196 737 198
rect 740 196 742 198
rect 745 196 747 198
rect 750 196 752 198
rect 577 194 579 196
rect 582 194 584 196
rect 587 194 589 196
rect 592 194 594 196
rect 597 194 599 196
rect 602 194 604 196
rect 607 194 609 196
rect 612 194 614 196
rect 617 194 619 196
rect 622 194 624 196
rect 627 194 629 196
rect 632 194 634 196
rect 637 194 639 196
rect 642 194 644 196
rect 647 194 649 196
rect 652 194 654 196
rect 675 191 677 193
rect 680 191 682 193
rect 685 191 687 193
rect 690 191 692 193
rect 695 191 697 193
rect 700 191 702 193
rect 705 191 707 193
rect 710 191 712 193
rect 715 191 717 193
rect 720 191 722 193
rect 725 191 727 193
rect 730 191 732 193
rect 735 191 737 193
rect 740 191 742 193
rect 745 191 747 193
rect 750 191 752 193
rect 577 189 579 191
rect 582 189 584 191
rect 587 189 589 191
rect 592 189 594 191
rect 597 189 599 191
rect 602 189 604 191
rect 607 189 609 191
rect 612 189 614 191
rect 617 189 619 191
rect 622 189 624 191
rect 627 189 629 191
rect 632 189 634 191
rect 637 189 639 191
rect 642 189 644 191
rect 647 189 649 191
rect 652 189 654 191
rect 675 186 677 188
rect 680 186 682 188
rect 685 186 687 188
rect 690 186 692 188
rect 695 186 697 188
rect 700 186 702 188
rect 705 186 707 188
rect 710 186 712 188
rect 715 186 717 188
rect 720 186 722 188
rect 725 186 727 188
rect 730 186 732 188
rect 735 186 737 188
rect 740 186 742 188
rect 745 186 747 188
rect 750 186 752 188
rect 577 184 579 186
rect 582 184 584 186
rect 587 184 589 186
rect 592 184 594 186
rect 597 184 599 186
rect 602 184 604 186
rect 607 184 609 186
rect 612 184 614 186
rect 617 184 619 186
rect 622 184 624 186
rect 627 184 629 186
rect 632 184 634 186
rect 637 184 639 186
rect 642 184 644 186
rect 647 184 649 186
rect 652 184 654 186
rect 675 181 677 183
rect 680 181 682 183
rect 685 181 687 183
rect 690 181 692 183
rect 695 181 697 183
rect 700 181 702 183
rect 705 181 707 183
rect 710 181 712 183
rect 715 181 717 183
rect 720 181 722 183
rect 725 181 727 183
rect 730 181 732 183
rect 735 181 737 183
rect 740 181 742 183
rect 745 181 747 183
rect 750 181 752 183
rect 577 179 579 181
rect 582 179 584 181
rect 587 179 589 181
rect 592 179 594 181
rect 597 179 599 181
rect 602 179 604 181
rect 607 179 609 181
rect 612 179 614 181
rect 617 179 619 181
rect 622 179 624 181
rect 627 179 629 181
rect 632 179 634 181
rect 637 179 639 181
rect 642 179 644 181
rect 647 179 649 181
rect 652 179 654 181
rect 675 176 677 178
rect 680 176 682 178
rect 685 176 687 178
rect 690 176 692 178
rect 695 176 697 178
rect 700 176 702 178
rect 705 176 707 178
rect 710 176 712 178
rect 715 176 717 178
rect 720 176 722 178
rect 725 176 727 178
rect 730 176 732 178
rect 735 176 737 178
rect 740 176 742 178
rect 745 176 747 178
rect 750 176 752 178
rect 577 174 579 176
rect 582 174 584 176
rect 587 174 589 176
rect 592 174 594 176
rect 597 174 599 176
rect 602 174 604 176
rect 607 174 609 176
rect 612 174 614 176
rect 617 174 619 176
rect 622 174 624 176
rect 627 174 629 176
rect 632 174 634 176
rect 637 174 639 176
rect 642 174 644 176
rect 647 174 649 176
rect 652 174 654 176
rect 675 171 677 173
rect 680 171 682 173
rect 685 171 687 173
rect 690 171 692 173
rect 695 171 697 173
rect 700 171 702 173
rect 705 171 707 173
rect 710 171 712 173
rect 715 171 717 173
rect 720 171 722 173
rect 725 171 727 173
rect 730 171 732 173
rect 735 171 737 173
rect 740 171 742 173
rect 745 171 747 173
rect 750 171 752 173
rect 577 169 579 171
rect 582 169 584 171
rect 587 169 589 171
rect 592 169 594 171
rect 597 169 599 171
rect 602 169 604 171
rect 607 169 609 171
rect 612 169 614 171
rect 617 169 619 171
rect 622 169 624 171
rect 627 169 629 171
rect 632 169 634 171
rect 637 169 639 171
rect 642 169 644 171
rect 647 169 649 171
rect 652 169 654 171
rect 675 166 677 168
rect 680 166 682 168
rect 685 166 687 168
rect 690 166 692 168
rect 695 166 697 168
rect 700 166 702 168
rect 705 166 707 168
rect 710 166 712 168
rect 715 166 717 168
rect 720 166 722 168
rect 725 166 727 168
rect 730 166 732 168
rect 735 166 737 168
rect 740 166 742 168
rect 745 166 747 168
rect 750 166 752 168
rect 577 164 579 166
rect 582 164 584 166
rect 587 164 589 166
rect 592 164 594 166
rect 597 164 599 166
rect 602 164 604 166
rect 607 164 609 166
rect 612 164 614 166
rect 617 164 619 166
rect 622 164 624 166
rect 627 164 629 166
rect 632 164 634 166
rect 637 164 639 166
rect 642 164 644 166
rect 647 164 649 166
rect 652 164 654 166
rect 675 161 677 163
rect 680 161 682 163
rect 685 161 687 163
rect 690 161 692 163
rect 695 161 697 163
rect 700 161 702 163
rect 705 161 707 163
rect 710 161 712 163
rect 715 161 717 163
rect 720 161 722 163
rect 725 161 727 163
rect 730 161 732 163
rect 735 161 737 163
rect 740 161 742 163
rect 745 161 747 163
rect 750 161 752 163
rect 577 159 579 161
rect 582 159 584 161
rect 587 159 589 161
rect 592 159 594 161
rect 597 159 599 161
rect 602 159 604 161
rect 607 159 609 161
rect 612 159 614 161
rect 617 159 619 161
rect 622 159 624 161
rect 627 159 629 161
rect 632 159 634 161
rect 637 159 639 161
rect 642 159 644 161
rect 647 159 649 161
rect 652 159 654 161
rect 675 156 677 158
rect 680 156 682 158
rect 685 156 687 158
rect 690 156 692 158
rect 695 156 697 158
rect 700 156 702 158
rect 705 156 707 158
rect 710 156 712 158
rect 715 156 717 158
rect 720 156 722 158
rect 725 156 727 158
rect 730 156 732 158
rect 735 156 737 158
rect 740 156 742 158
rect 745 156 747 158
rect 750 156 752 158
rect 577 154 579 156
rect 582 154 584 156
rect 587 154 589 156
rect 592 154 594 156
rect 597 154 599 156
rect 602 154 604 156
rect 607 154 609 156
rect 612 154 614 156
rect 617 154 619 156
rect 622 154 624 156
rect 627 154 629 156
rect 632 154 634 156
rect 637 154 639 156
rect 642 154 644 156
rect 647 154 649 156
rect 652 154 654 156
rect 675 151 677 153
rect 680 151 682 153
rect 685 151 687 153
rect 690 151 692 153
rect 695 151 697 153
rect 700 151 702 153
rect 705 151 707 153
rect 710 151 712 153
rect 715 151 717 153
rect 720 151 722 153
rect 725 151 727 153
rect 730 151 732 153
rect 735 151 737 153
rect 740 151 742 153
rect 745 151 747 153
rect 750 151 752 153
rect 577 149 579 151
rect 582 149 584 151
rect 587 149 589 151
rect 592 149 594 151
rect 597 149 599 151
rect 602 149 604 151
rect 607 149 609 151
rect 612 149 614 151
rect 617 149 619 151
rect 622 149 624 151
rect 627 149 629 151
rect 632 149 634 151
rect 637 149 639 151
rect 642 149 644 151
rect 647 149 649 151
rect 652 149 654 151
rect 675 146 677 148
rect 680 146 682 148
rect 685 146 687 148
rect 690 146 692 148
rect 695 146 697 148
rect 700 146 702 148
rect 705 146 707 148
rect 710 146 712 148
rect 715 146 717 148
rect 720 146 722 148
rect 725 146 727 148
rect 730 146 732 148
rect 735 146 737 148
rect 740 146 742 148
rect 745 146 747 148
rect 750 146 752 148
rect 577 144 579 146
rect 582 144 584 146
rect 587 144 589 146
rect 592 144 594 146
rect 597 144 599 146
rect 602 144 604 146
rect 607 144 609 146
rect 612 144 614 146
rect 617 144 619 146
rect 622 144 624 146
rect 627 144 629 146
rect 632 144 634 146
rect 637 144 639 146
rect 642 144 644 146
rect 647 144 649 146
rect 652 144 654 146
rect 675 141 677 143
rect 680 141 682 143
rect 685 141 687 143
rect 690 141 692 143
rect 695 141 697 143
rect 700 141 702 143
rect 705 141 707 143
rect 710 141 712 143
rect 715 141 717 143
rect 720 141 722 143
rect 725 141 727 143
rect 730 141 732 143
rect 735 141 737 143
rect 740 141 742 143
rect 745 141 747 143
rect 750 141 752 143
rect 577 139 579 141
rect 582 139 584 141
rect 587 139 589 141
rect 592 139 594 141
rect 597 139 599 141
rect 602 139 604 141
rect 607 139 609 141
rect 612 139 614 141
rect 617 139 619 141
rect 622 139 624 141
rect 627 139 629 141
rect 632 139 634 141
rect 637 139 639 141
rect 642 139 644 141
rect 647 139 649 141
rect 652 139 654 141
rect 675 136 677 138
rect 680 136 682 138
rect 685 136 687 138
rect 690 136 692 138
rect 695 136 697 138
rect 700 136 702 138
rect 705 136 707 138
rect 710 136 712 138
rect 715 136 717 138
rect 720 136 722 138
rect 725 136 727 138
rect 730 136 732 138
rect 735 136 737 138
rect 740 136 742 138
rect 745 136 747 138
rect 750 136 752 138
rect 577 134 579 136
rect 582 134 584 136
rect 587 134 589 136
rect 592 134 594 136
rect 597 134 599 136
rect 602 134 604 136
rect 607 134 609 136
rect 612 134 614 136
rect 617 134 619 136
rect 622 134 624 136
rect 627 134 629 136
rect 632 134 634 136
rect 637 134 639 136
rect 642 134 644 136
rect 647 134 649 136
rect 652 134 654 136
rect 675 131 677 133
rect 680 131 682 133
rect 685 131 687 133
rect 690 131 692 133
rect 695 131 697 133
rect 700 131 702 133
rect 705 131 707 133
rect 710 131 712 133
rect 715 131 717 133
rect 720 131 722 133
rect 725 131 727 133
rect 730 131 732 133
rect 735 131 737 133
rect 740 131 742 133
rect 745 131 747 133
rect 750 131 752 133
rect 577 129 579 131
rect 582 129 584 131
rect 587 129 589 131
rect 592 129 594 131
rect 597 129 599 131
rect 602 129 604 131
rect 607 129 609 131
rect 612 129 614 131
rect 617 129 619 131
rect 622 129 624 131
rect 627 129 629 131
rect 632 129 634 131
rect 637 129 639 131
rect 642 129 644 131
rect 647 129 649 131
rect 652 129 654 131
rect 675 126 677 128
rect 680 126 682 128
rect 685 126 687 128
rect 690 126 692 128
rect 695 126 697 128
rect 700 126 702 128
rect 705 126 707 128
rect 710 126 712 128
rect 715 126 717 128
rect 720 126 722 128
rect 725 126 727 128
rect 730 126 732 128
rect 735 126 737 128
rect 740 126 742 128
rect 745 126 747 128
rect 750 126 752 128
rect 577 124 579 126
rect 582 124 584 126
rect 587 124 589 126
rect 592 124 594 126
rect 597 124 599 126
rect 602 124 604 126
rect 607 124 609 126
rect 612 124 614 126
rect 617 124 619 126
rect 622 124 624 126
rect 627 124 629 126
rect 632 124 634 126
rect 637 124 639 126
rect 642 124 644 126
rect 647 124 649 126
rect 652 124 654 126
rect 675 121 677 123
rect 680 121 682 123
rect 685 121 687 123
rect 690 121 692 123
rect 695 121 697 123
rect 700 121 702 123
rect 705 121 707 123
rect 710 121 712 123
rect 715 121 717 123
rect 720 121 722 123
rect 725 121 727 123
rect 730 121 732 123
rect 735 121 737 123
rect 740 121 742 123
rect 745 121 747 123
rect 750 121 752 123
rect 577 119 579 121
rect 582 119 584 121
rect 587 119 589 121
rect 592 119 594 121
rect 597 119 599 121
rect 602 119 604 121
rect 607 119 609 121
rect 612 119 614 121
rect 617 119 619 121
rect 622 119 624 121
rect 627 119 629 121
rect 632 119 634 121
rect 637 119 639 121
rect 642 119 644 121
rect 647 119 649 121
rect 652 119 654 121
rect 675 116 677 118
rect 680 116 682 118
rect 685 116 687 118
rect 690 116 692 118
rect 695 116 697 118
rect 700 116 702 118
rect 705 116 707 118
rect 710 116 712 118
rect 715 116 717 118
rect 720 116 722 118
rect 725 116 727 118
rect 730 116 732 118
rect 735 116 737 118
rect 740 116 742 118
rect 745 116 747 118
rect 750 116 752 118
rect 577 114 579 116
rect 582 114 584 116
rect 587 114 589 116
rect 592 114 594 116
rect 597 114 599 116
rect 602 114 604 116
rect 607 114 609 116
rect 612 114 614 116
rect 617 114 619 116
rect 622 114 624 116
rect 627 114 629 116
rect 632 114 634 116
rect 637 114 639 116
rect 642 114 644 116
rect 647 114 649 116
rect 652 114 654 116
rect 675 111 677 113
rect 680 111 682 113
rect 685 111 687 113
rect 690 111 692 113
rect 695 111 697 113
rect 700 111 702 113
rect 705 111 707 113
rect 710 111 712 113
rect 715 111 717 113
rect 720 111 722 113
rect 725 111 727 113
rect 730 111 732 113
rect 735 111 737 113
rect 740 111 742 113
rect 745 111 747 113
rect 750 111 752 113
rect 577 109 579 111
rect 582 109 584 111
rect 587 109 589 111
rect 592 109 594 111
rect 597 109 599 111
rect 602 109 604 111
rect 607 109 609 111
rect 612 109 614 111
rect 617 109 619 111
rect 622 109 624 111
rect 627 109 629 111
rect 632 109 634 111
rect 637 109 639 111
rect 642 109 644 111
rect 647 109 649 111
rect 652 109 654 111
rect 675 106 677 108
rect 680 106 682 108
rect 685 106 687 108
rect 690 106 692 108
rect 695 106 697 108
rect 700 106 702 108
rect 705 106 707 108
rect 710 106 712 108
rect 715 106 717 108
rect 720 106 722 108
rect 725 106 727 108
rect 730 106 732 108
rect 735 106 737 108
rect 740 106 742 108
rect 745 106 747 108
rect 750 106 752 108
rect 577 104 579 106
rect 582 104 584 106
rect 587 104 589 106
rect 592 104 594 106
rect 597 104 599 106
rect 602 104 604 106
rect 607 104 609 106
rect 612 104 614 106
rect 617 104 619 106
rect 622 104 624 106
rect 627 104 629 106
rect 632 104 634 106
rect 637 104 639 106
rect 642 104 644 106
rect 647 104 649 106
rect 652 104 654 106
rect 675 101 677 103
rect 680 101 682 103
rect 685 101 687 103
rect 690 101 692 103
rect 695 101 697 103
rect 700 101 702 103
rect 705 101 707 103
rect 710 101 712 103
rect 715 101 717 103
rect 720 101 722 103
rect 725 101 727 103
rect 730 101 732 103
rect 735 101 737 103
rect 740 101 742 103
rect 745 101 747 103
rect 750 101 752 103
rect 577 99 579 101
rect 582 99 584 101
rect 587 99 589 101
rect 592 99 594 101
rect 597 99 599 101
rect 602 99 604 101
rect 607 99 609 101
rect 612 99 614 101
rect 617 99 619 101
rect 622 99 624 101
rect 627 99 629 101
rect 632 99 634 101
rect 637 99 639 101
rect 642 99 644 101
rect 647 99 649 101
rect 652 99 654 101
rect 675 96 677 98
rect 680 96 682 98
rect 685 96 687 98
rect 690 96 692 98
rect 695 96 697 98
rect 700 96 702 98
rect 705 96 707 98
rect 710 96 712 98
rect 715 96 717 98
rect 720 96 722 98
rect 725 96 727 98
rect 730 96 732 98
rect 735 96 737 98
rect 740 96 742 98
rect 745 96 747 98
rect 750 96 752 98
rect 577 94 579 96
rect 582 94 584 96
rect 587 94 589 96
rect 592 94 594 96
rect 597 94 599 96
rect 602 94 604 96
rect 607 94 609 96
rect 612 94 614 96
rect 617 94 619 96
rect 622 94 624 96
rect 627 94 629 96
rect 632 94 634 96
rect 637 94 639 96
rect 642 94 644 96
rect 647 94 649 96
rect 652 94 654 96
rect 675 91 677 93
rect 680 91 682 93
rect 685 91 687 93
rect 690 91 692 93
rect 695 91 697 93
rect 700 91 702 93
rect 705 91 707 93
rect 710 91 712 93
rect 715 91 717 93
rect 720 91 722 93
rect 725 91 727 93
rect 730 91 732 93
rect 735 91 737 93
rect 740 91 742 93
rect 745 91 747 93
rect 750 91 752 93
rect 577 89 579 91
rect 582 89 584 91
rect 587 89 589 91
rect 592 89 594 91
rect 597 89 599 91
rect 602 89 604 91
rect 607 89 609 91
rect 612 89 614 91
rect 617 89 619 91
rect 622 89 624 91
rect 627 89 629 91
rect 632 89 634 91
rect 637 89 639 91
rect 642 89 644 91
rect 647 89 649 91
rect 652 89 654 91
rect 675 86 677 88
rect 680 86 682 88
rect 685 86 687 88
rect 690 86 692 88
rect 695 86 697 88
rect 700 86 702 88
rect 705 86 707 88
rect 710 86 712 88
rect 715 86 717 88
rect 720 86 722 88
rect 725 86 727 88
rect 730 86 732 88
rect 735 86 737 88
rect 740 86 742 88
rect 745 86 747 88
rect 750 86 752 88
rect 577 84 579 86
rect 582 84 584 86
rect 587 84 589 86
rect 592 84 594 86
rect 597 84 599 86
rect 602 84 604 86
rect 607 84 609 86
rect 612 84 614 86
rect 617 84 619 86
rect 622 84 624 86
rect 627 84 629 86
rect 632 84 634 86
rect 637 84 639 86
rect 642 84 644 86
rect 647 84 649 86
rect 652 84 654 86
rect 675 81 677 83
rect 680 81 682 83
rect 685 81 687 83
rect 690 81 692 83
rect 695 81 697 83
rect 700 81 702 83
rect 705 81 707 83
rect 710 81 712 83
rect 715 81 717 83
rect 720 81 722 83
rect 725 81 727 83
rect 730 81 732 83
rect 735 81 737 83
rect 740 81 742 83
rect 745 81 747 83
rect 750 81 752 83
rect 577 79 579 81
rect 582 79 584 81
rect 587 79 589 81
rect 592 79 594 81
rect 597 79 599 81
rect 602 79 604 81
rect 607 79 609 81
rect 612 79 614 81
rect 617 79 619 81
rect 622 79 624 81
rect 627 79 629 81
rect 632 79 634 81
rect 637 79 639 81
rect 642 79 644 81
rect 647 79 649 81
rect 652 79 654 81
rect 675 76 677 78
rect 680 76 682 78
rect 685 76 687 78
rect 690 76 692 78
rect 695 76 697 78
rect 700 76 702 78
rect 705 76 707 78
rect 710 76 712 78
rect 715 76 717 78
rect 720 76 722 78
rect 725 76 727 78
rect 730 76 732 78
rect 735 76 737 78
rect 740 76 742 78
rect 745 76 747 78
rect 750 76 752 78
rect 577 74 579 76
rect 582 74 584 76
rect 587 74 589 76
rect 592 74 594 76
rect 597 74 599 76
rect 602 74 604 76
rect 607 74 609 76
rect 612 74 614 76
rect 617 74 619 76
rect 622 74 624 76
rect 627 74 629 76
rect 632 74 634 76
rect 637 74 639 76
rect 642 74 644 76
rect 647 74 649 76
rect 652 74 654 76
rect 675 71 677 73
rect 680 71 682 73
rect 685 71 687 73
rect 690 71 692 73
rect 695 71 697 73
rect 700 71 702 73
rect 705 71 707 73
rect 710 71 712 73
rect 715 71 717 73
rect 720 71 722 73
rect 725 71 727 73
rect 730 71 732 73
rect 735 71 737 73
rect 740 71 742 73
rect 745 71 747 73
rect 750 71 752 73
rect 577 69 579 71
rect 582 69 584 71
rect 587 69 589 71
rect 592 69 594 71
rect 597 69 599 71
rect 602 69 604 71
rect 607 69 609 71
rect 612 69 614 71
rect 617 69 619 71
rect 622 69 624 71
rect 627 69 629 71
rect 632 69 634 71
rect 637 69 639 71
rect 642 69 644 71
rect 647 69 649 71
rect 652 69 654 71
rect 675 66 677 68
rect 680 66 682 68
rect 685 66 687 68
rect 690 66 692 68
rect 695 66 697 68
rect 700 66 702 68
rect 705 66 707 68
rect 710 66 712 68
rect 715 66 717 68
rect 720 66 722 68
rect 725 66 727 68
rect 730 66 732 68
rect 735 66 737 68
rect 740 66 742 68
rect 745 66 747 68
rect 750 66 752 68
rect 577 64 579 66
rect 582 64 584 66
rect 587 64 589 66
rect 592 64 594 66
rect 597 64 599 66
rect 602 64 604 66
rect 607 64 609 66
rect 612 64 614 66
rect 617 64 619 66
rect 622 64 624 66
rect 627 64 629 66
rect 632 64 634 66
rect 637 64 639 66
rect 642 64 644 66
rect 647 64 649 66
rect 652 64 654 66
rect 675 61 677 63
rect 680 61 682 63
rect 685 61 687 63
rect 690 61 692 63
rect 695 61 697 63
rect 700 61 702 63
rect 705 61 707 63
rect 710 61 712 63
rect 715 61 717 63
rect 720 61 722 63
rect 725 61 727 63
rect 730 61 732 63
rect 735 61 737 63
rect 740 61 742 63
rect 745 61 747 63
rect 750 61 752 63
rect 577 59 579 61
rect 582 59 584 61
rect 587 59 589 61
rect 592 59 594 61
rect 597 59 599 61
rect 602 59 604 61
rect 607 59 609 61
rect 612 59 614 61
rect 617 59 619 61
rect 622 59 624 61
rect 627 59 629 61
rect 632 59 634 61
rect 637 59 639 61
rect 642 59 644 61
rect 647 59 649 61
rect 652 59 654 61
rect 675 56 677 58
rect 680 56 682 58
rect 685 56 687 58
rect 690 56 692 58
rect 695 56 697 58
rect 700 56 702 58
rect 705 56 707 58
rect 710 56 712 58
rect 715 56 717 58
rect 720 56 722 58
rect 725 56 727 58
rect 730 56 732 58
rect 735 56 737 58
rect 740 56 742 58
rect 745 56 747 58
rect 750 56 752 58
rect 577 54 579 56
rect 582 54 584 56
rect 587 54 589 56
rect 592 54 594 56
rect 597 54 599 56
rect 602 54 604 56
rect 607 54 609 56
rect 612 54 614 56
rect 617 54 619 56
rect 622 54 624 56
rect 627 54 629 56
rect 632 54 634 56
rect 637 54 639 56
rect 642 54 644 56
rect 647 54 649 56
rect 652 54 654 56
rect 675 51 677 53
rect 680 51 682 53
rect 685 51 687 53
rect 690 51 692 53
rect 695 51 697 53
rect 700 51 702 53
rect 705 51 707 53
rect 710 51 712 53
rect 715 51 717 53
rect 720 51 722 53
rect 725 51 727 53
rect 730 51 732 53
rect 735 51 737 53
rect 740 51 742 53
rect 745 51 747 53
rect 750 51 752 53
rect 577 49 579 51
rect 582 49 584 51
rect 587 49 589 51
rect 592 49 594 51
rect 597 49 599 51
rect 602 49 604 51
rect 607 49 609 51
rect 612 49 614 51
rect 617 49 619 51
rect 622 49 624 51
rect 627 49 629 51
rect 632 49 634 51
rect 637 49 639 51
rect 642 49 644 51
rect 647 49 649 51
rect 652 49 654 51
rect 675 46 677 48
rect 680 46 682 48
rect 685 46 687 48
rect 690 46 692 48
rect 695 46 697 48
rect 700 46 702 48
rect 705 46 707 48
rect 710 46 712 48
rect 715 46 717 48
rect 720 46 722 48
rect 725 46 727 48
rect 730 46 732 48
rect 735 46 737 48
rect 740 46 742 48
rect 745 46 747 48
rect 750 46 752 48
rect 577 44 579 46
rect 582 44 584 46
rect 587 44 589 46
rect 592 44 594 46
rect 597 44 599 46
rect 602 44 604 46
rect 607 44 609 46
rect 612 44 614 46
rect 617 44 619 46
rect 622 44 624 46
rect 627 44 629 46
rect 632 44 634 46
rect 637 44 639 46
rect 642 44 644 46
rect 647 44 649 46
rect 652 44 654 46
rect 675 41 677 43
rect 680 41 682 43
rect 685 41 687 43
rect 690 41 692 43
rect 695 41 697 43
rect 700 41 702 43
rect 705 41 707 43
rect 710 41 712 43
rect 715 41 717 43
rect 720 41 722 43
rect 725 41 727 43
rect 730 41 732 43
rect 735 41 737 43
rect 740 41 742 43
rect 745 41 747 43
rect 750 41 752 43
rect 577 39 579 41
rect 582 39 584 41
rect 587 39 589 41
rect 592 39 594 41
rect 597 39 599 41
rect 602 39 604 41
rect 607 39 609 41
rect 612 39 614 41
rect 617 39 619 41
rect 622 39 624 41
rect 627 39 629 41
rect 632 39 634 41
rect 637 39 639 41
rect 642 39 644 41
rect 647 39 649 41
rect 652 39 654 41
rect 675 36 677 38
rect 680 36 682 38
rect 685 36 687 38
rect 690 36 692 38
rect 695 36 697 38
rect 700 36 702 38
rect 705 36 707 38
rect 710 36 712 38
rect 715 36 717 38
rect 720 36 722 38
rect 725 36 727 38
rect 730 36 732 38
rect 735 36 737 38
rect 740 36 742 38
rect 745 36 747 38
rect 750 36 752 38
rect 577 34 579 36
rect 582 34 584 36
rect 587 34 589 36
rect 592 34 594 36
rect 597 34 599 36
rect 602 34 604 36
rect 607 34 609 36
rect 612 34 614 36
rect 617 34 619 36
rect 622 34 624 36
rect 627 34 629 36
rect 632 34 634 36
rect 637 34 639 36
rect 642 34 644 36
rect 647 34 649 36
rect 652 34 654 36
rect 675 31 677 33
rect 680 31 682 33
rect 685 31 687 33
rect 690 31 692 33
rect 695 31 697 33
rect 700 31 702 33
rect 705 31 707 33
rect 710 31 712 33
rect 715 31 717 33
rect 720 31 722 33
rect 725 31 727 33
rect 730 31 732 33
rect 735 31 737 33
rect 740 31 742 33
rect 745 31 747 33
rect 750 31 752 33
rect 577 29 579 31
rect 582 29 584 31
rect 587 29 589 31
rect 592 29 594 31
rect 597 29 599 31
rect 602 29 604 31
rect 607 29 609 31
rect 612 29 614 31
rect 617 29 619 31
rect 622 29 624 31
rect 627 29 629 31
rect 632 29 634 31
rect 637 29 639 31
rect 642 29 644 31
rect 647 29 649 31
rect 652 29 654 31
rect 675 26 677 28
rect 680 26 682 28
rect 685 26 687 28
rect 690 26 692 28
rect 695 26 697 28
rect 700 26 702 28
rect 705 26 707 28
rect 710 26 712 28
rect 715 26 717 28
rect 720 26 722 28
rect 725 26 727 28
rect 730 26 732 28
rect 735 26 737 28
rect 740 26 742 28
rect 745 26 747 28
rect 750 26 752 28
rect 577 24 579 26
rect 582 24 584 26
rect 587 24 589 26
rect 592 24 594 26
rect 597 24 599 26
rect 602 24 604 26
rect 607 24 609 26
rect 612 24 614 26
rect 617 24 619 26
rect 622 24 624 26
rect 627 24 629 26
rect 632 24 634 26
rect 637 24 639 26
rect 642 24 644 26
rect 647 24 649 26
rect 652 24 654 26
rect 675 21 677 23
rect 680 21 682 23
rect 685 21 687 23
rect 690 21 692 23
rect 695 21 697 23
rect 700 21 702 23
rect 705 21 707 23
rect 710 21 712 23
rect 715 21 717 23
rect 720 21 722 23
rect 725 21 727 23
rect 730 21 732 23
rect 735 21 737 23
rect 740 21 742 23
rect 745 21 747 23
rect 750 21 752 23
rect 577 19 579 21
rect 582 19 584 21
rect 587 19 589 21
rect 592 19 594 21
rect 597 19 599 21
rect 602 19 604 21
rect 607 19 609 21
rect 612 19 614 21
rect 617 19 619 21
rect 622 19 624 21
rect 627 19 629 21
rect 632 19 634 21
rect 637 19 639 21
rect 642 19 644 21
rect 647 19 649 21
rect 652 19 654 21
rect 675 16 677 18
rect 680 16 682 18
rect 685 16 687 18
rect 690 16 692 18
rect 695 16 697 18
rect 700 16 702 18
rect 705 16 707 18
rect 710 16 712 18
rect 715 16 717 18
rect 720 16 722 18
rect 725 16 727 18
rect 730 16 732 18
rect 735 16 737 18
rect 740 16 742 18
rect 745 16 747 18
rect 750 16 752 18
rect 577 14 579 16
rect 582 14 584 16
rect 587 14 589 16
rect 592 14 594 16
rect 597 14 599 16
rect 602 14 604 16
rect 607 14 609 16
rect 612 14 614 16
rect 617 14 619 16
rect 622 14 624 16
rect 627 14 629 16
rect 632 14 634 16
rect 637 14 639 16
rect 642 14 644 16
rect 647 14 649 16
rect 652 14 654 16
rect 675 11 677 13
rect 680 11 682 13
rect 685 11 687 13
rect 690 11 692 13
rect 695 11 697 13
rect 700 11 702 13
rect 705 11 707 13
rect 710 11 712 13
rect 715 11 717 13
rect 720 11 722 13
rect 725 11 727 13
rect 730 11 732 13
rect 735 11 737 13
rect 740 11 742 13
rect 745 11 747 13
rect 750 11 752 13
rect 577 9 579 11
rect 582 9 584 11
rect 587 9 589 11
rect 592 9 594 11
rect 597 9 599 11
rect 602 9 604 11
rect 607 9 609 11
rect 612 9 614 11
rect 617 9 619 11
rect 622 9 624 11
rect 627 9 629 11
rect 632 9 634 11
rect 637 9 639 11
rect 642 9 644 11
rect 647 9 649 11
rect 652 9 654 11
rect 675 6 677 8
rect 680 6 682 8
rect 685 6 687 8
rect 690 6 692 8
rect 695 6 697 8
rect 700 6 702 8
rect 705 6 707 8
rect 710 6 712 8
rect 715 6 717 8
rect 720 6 722 8
rect 725 6 727 8
rect 730 6 732 8
rect 735 6 737 8
rect 740 6 742 8
rect 745 6 747 8
rect 750 6 752 8
rect 577 4 579 6
rect 582 4 584 6
rect 587 4 589 6
rect 592 4 594 6
rect 597 4 599 6
rect 602 4 604 6
rect 607 4 609 6
rect 612 4 614 6
rect 617 4 619 6
rect 622 4 624 6
rect 627 4 629 6
rect 632 4 634 6
rect 637 4 639 6
rect 642 4 644 6
rect 647 4 649 6
rect 652 4 654 6
rect 675 1 677 3
rect 680 1 682 3
rect 685 1 687 3
rect 690 1 692 3
rect 695 1 697 3
rect 700 1 702 3
rect 705 1 707 3
rect 710 1 712 3
rect 715 1 717 3
rect 720 1 722 3
rect 725 1 727 3
rect 730 1 732 3
rect 735 1 737 3
rect 740 1 742 3
rect 745 1 747 3
rect 750 1 752 3
<< end >>
